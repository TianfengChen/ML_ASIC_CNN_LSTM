VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LDO_Top_int
  CLASS BLOCK ;
  ORIGIN 0.34 96.81 ;
  FOREIGN LDO_Top_int -0.34 -96.81 ;
  SIZE 125.45 BY 47.85 ;
  SYMMETRY X Y R90 ;
  PIN SW[2]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 22.94 -49.16 23.14 -48.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.68 -62.45 23.4 -61.73 ;
      LAYER M2 ;
        RECT 22.74 -62.39 23.34 -61.79 ;
      LAYER M3 ;
        RECT 22.74 -62.39 23.34 -61.79 ;
      LAYER V2 ;
        RECT 22.74 -61.99 22.94 -61.79 ;
        RECT 22.74 -62.39 22.94 -62.19 ;
        RECT 23.14 -61.99 23.34 -61.79 ;
        RECT 23.14 -62.39 23.34 -62.19 ;
      LAYER V1 ;
        RECT 22.74 -61.99 22.94 -61.79 ;
        RECT 22.74 -62.39 22.94 -62.19 ;
        RECT 23.14 -61.99 23.34 -61.79 ;
        RECT 23.14 -62.39 23.34 -62.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -62 24.6 -61.84 ;
    END
  END SW[2]
  PIN SW[1]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 22.19 -49.16 22.39 -48.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.93 -58.78 22.65 -58.06 ;
      LAYER M2 ;
        RECT 21.99 -58.72 22.59 -58.12 ;
      LAYER M3 ;
        RECT 21.99 -58.72 22.59 -58.12 ;
      LAYER V2 ;
        RECT 21.99 -58.32 22.19 -58.12 ;
        RECT 21.99 -58.72 22.19 -58.52 ;
        RECT 22.39 -58.32 22.59 -58.12 ;
        RECT 22.39 -58.72 22.59 -58.52 ;
      LAYER V1 ;
        RECT 21.99 -58.32 22.19 -58.12 ;
        RECT 21.99 -58.72 22.19 -58.52 ;
        RECT 22.39 -58.32 22.59 -58.12 ;
        RECT 22.39 -58.72 22.59 -58.52 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -58.64 24.6 -58.48 ;
    END
  END SW[1]
  PIN SW[0]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 21.42 -49.16 21.62 -48.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.16 -55.07 21.88 -54.35 ;
      LAYER M2 ;
        RECT 21.22 -55.01 21.82 -54.41 ;
      LAYER M3 ;
        RECT 21.22 -55.01 21.82 -54.41 ;
      LAYER V2 ;
        RECT 21.22 -54.61 21.42 -54.41 ;
        RECT 21.22 -55.01 21.42 -54.81 ;
        RECT 21.62 -54.61 21.82 -54.41 ;
        RECT 21.62 -55.01 21.82 -54.81 ;
      LAYER V1 ;
        RECT 21.22 -54.61 21.42 -54.41 ;
        RECT 21.22 -55.01 21.42 -54.81 ;
        RECT 21.62 -54.61 21.82 -54.41 ;
        RECT 21.62 -55.01 21.82 -54.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -54.8 24.6 -54.64 ;
    END
  END SW[0]
  PIN VB
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 47.82 -96.81 48.22 -96.41 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1 -71.26 50.37 -71.16 ;
        RECT 50.1 -71.26 50.3 -71.06 ;
      LAYER V1 ;
        RECT 50.1 -71.26 50.3 -71.06 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.93 -71.75 33.25 -71.43 ;
        RECT 32.93 -71.35 33.25 -71.03 ;
      LAYER M2 ;
        RECT 32.92 -71.56 33.32 -71.16 ;
        RECT 32.99 -71.69 33.19 -71.09 ;
      LAYER V1 ;
        RECT 32.99 -71.29 33.19 -71.09 ;
        RECT 32.99 -71.69 33.19 -71.49 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.8 -70.23 46.96 -70.07 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.8 -68.77 47.04 -68.53 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.08 -68.77 50.32 -68.53 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.04 -71.72 50.36 -71.4 ;
      LAYER M2 ;
        RECT 50.1 -71.56 50.37 -71.46 ;
        RECT 50.1 -71.66 50.3 -71.46 ;
      LAYER V1 ;
        RECT 50.1 -71.66 50.3 -71.46 ;
    END
  END VB
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 94.63 -96.34 95.61 -95.34 ;
      LAYER V2 ;
        RECT 94.57 -95.54 94.77 -95.34 ;
        RECT 94.57 -95.94 94.77 -95.74 ;
        RECT 94.57 -96.34 94.77 -96.14 ;
        RECT 94.97 -95.54 95.17 -95.34 ;
        RECT 94.97 -95.94 95.17 -95.74 ;
        RECT 94.97 -96.34 95.17 -96.14 ;
        RECT 95.37 -95.54 95.57 -95.34 ;
        RECT 95.37 -95.94 95.57 -95.74 ;
        RECT 95.37 -96.34 95.57 -96.14 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.05 -53.02 35.05 -52.02 ;
      LAYER M3 ;
        RECT 34.05 -53.02 35.03 -52.02 ;
      LAYER V2 ;
        RECT 34.05 -52.22 34.25 -52.02 ;
        RECT 34.05 -52.62 34.25 -52.42 ;
        RECT 34.05 -53.02 34.25 -52.82 ;
        RECT 34.45 -52.22 34.65 -52.02 ;
        RECT 34.45 -52.62 34.65 -52.42 ;
        RECT 34.45 -53.02 34.65 -52.82 ;
        RECT 34.85 -52.22 35.05 -52.02 ;
        RECT 34.85 -52.62 35.05 -52.42 ;
        RECT 34.85 -53.02 35.05 -52.82 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.48 -54.26 28.76 -54 ;
        RECT 28.48 -54.29 28.75 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.48 -55.78 28.76 -55.61 ;
        RECT 28.48 -55.78 28.75 -55.49 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.44 -54.26 29.72 -54 ;
        RECT 29.44 -54.29 29.71 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.45 -55.78 29.73 -55.61 ;
        RECT 29.45 -55.78 29.72 -55.49 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.4 -54.26 30.68 -54 ;
        RECT 30.4 -54.29 30.67 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.42 -55.78 30.7 -55.49 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.36 -54.26 31.64 -54 ;
        RECT 31.36 -54.29 31.63 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.53 -55.29 31.67 -55.13 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.39 -55.78 31.67 -55.49 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4 -54.06 34.74 -53.78 ;
      LAYER M2 ;
        RECT 34.42 -54.02 34.72 -53.74 ;
      LAYER V1 ;
        RECT 34.47 -54.02 34.67 -53.82 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.12 -71.01 65.38 -70.77 ;
      LAYER M2 ;
        RECT 65.12 -71.01 65.38 -70.77 ;
      LAYER V1 ;
        RECT 65.15 -71.03 65.35 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.12 -90.61 65.38 -90.37 ;
      LAYER V1 ;
        RECT 65.15 -90.55 65.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.08 -71.01 66.34 -70.77 ;
      LAYER M2 ;
        RECT 66.08 -71.01 66.34 -70.77 ;
      LAYER V1 ;
        RECT 66.11 -71.03 66.31 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.08 -90.61 66.34 -90.37 ;
      LAYER V1 ;
        RECT 66.11 -90.55 66.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.04 -71.01 67.3 -70.77 ;
      LAYER M2 ;
        RECT 67.04 -71.01 67.3 -70.77 ;
      LAYER V1 ;
        RECT 67.07 -71.03 67.27 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.04 -90.61 67.3 -90.37 ;
      LAYER V1 ;
        RECT 67.07 -90.55 67.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68 -71.01 68.26 -70.77 ;
      LAYER M2 ;
        RECT 68 -71.01 68.26 -70.77 ;
      LAYER V1 ;
        RECT 68.03 -71.03 68.23 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 68 -90.61 68.26 -90.37 ;
      LAYER V1 ;
        RECT 68.03 -90.55 68.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.96 -71.01 69.22 -70.77 ;
      LAYER M2 ;
        RECT 68.96 -71.01 69.22 -70.77 ;
      LAYER V1 ;
        RECT 68.99 -71.03 69.19 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.96 -90.61 69.22 -90.37 ;
      LAYER V1 ;
        RECT 68.99 -90.55 69.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.92 -71.01 70.18 -70.77 ;
      LAYER M2 ;
        RECT 69.92 -71.01 70.18 -70.77 ;
      LAYER V1 ;
        RECT 69.95 -71.03 70.15 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.92 -90.61 70.18 -90.37 ;
      LAYER V1 ;
        RECT 69.95 -90.55 70.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.88 -71.01 71.14 -70.77 ;
      LAYER M2 ;
        RECT 70.88 -71.01 71.14 -70.77 ;
      LAYER V1 ;
        RECT 70.91 -71.03 71.11 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.88 -90.61 71.14 -90.37 ;
      LAYER V1 ;
        RECT 70.91 -90.55 71.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.84 -71.01 72.1 -70.77 ;
      LAYER M2 ;
        RECT 71.84 -71.01 72.1 -70.77 ;
      LAYER V1 ;
        RECT 71.87 -71.03 72.07 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.84 -90.61 72.1 -90.37 ;
      LAYER V1 ;
        RECT 71.87 -90.55 72.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.8 -71.01 73.06 -70.77 ;
      LAYER M2 ;
        RECT 72.8 -71.01 73.06 -70.77 ;
      LAYER V1 ;
        RECT 72.83 -71.03 73.03 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.8 -90.61 73.06 -90.37 ;
      LAYER V1 ;
        RECT 72.83 -90.55 73.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.76 -71.01 74.02 -70.77 ;
      LAYER M2 ;
        RECT 73.76 -71.01 74.02 -70.77 ;
      LAYER V1 ;
        RECT 73.79 -71.03 73.99 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.76 -90.61 74.02 -90.37 ;
      LAYER V1 ;
        RECT 73.79 -90.55 73.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.72 -71.01 74.98 -70.77 ;
      LAYER M2 ;
        RECT 74.72 -71.01 74.98 -70.77 ;
      LAYER V1 ;
        RECT 74.75 -71.03 74.95 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.72 -90.61 74.98 -90.37 ;
      LAYER V1 ;
        RECT 74.75 -90.55 74.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.68 -71.01 75.94 -70.77 ;
      LAYER M2 ;
        RECT 75.68 -71.01 75.94 -70.77 ;
      LAYER V1 ;
        RECT 75.71 -71.03 75.91 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.68 -90.61 75.94 -90.37 ;
      LAYER V1 ;
        RECT 75.71 -90.55 75.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.64 -71.01 76.9 -70.77 ;
      LAYER M2 ;
        RECT 76.64 -71.01 76.9 -70.77 ;
      LAYER V1 ;
        RECT 76.67 -71.03 76.87 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.64 -90.61 76.9 -90.37 ;
      LAYER V1 ;
        RECT 76.67 -90.55 76.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.6 -71.01 77.86 -70.77 ;
      LAYER M2 ;
        RECT 77.6 -71.01 77.86 -70.77 ;
      LAYER V1 ;
        RECT 77.63 -71.03 77.83 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.6 -90.61 77.86 -90.37 ;
      LAYER V1 ;
        RECT 77.63 -90.55 77.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.56 -71.01 78.82 -70.77 ;
      LAYER M2 ;
        RECT 78.56 -71.01 78.82 -70.77 ;
      LAYER V1 ;
        RECT 78.59 -71.03 78.79 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.56 -90.61 78.82 -90.37 ;
      LAYER V1 ;
        RECT 78.59 -90.55 78.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.52 -71.01 79.78 -70.77 ;
      LAYER M2 ;
        RECT 79.52 -71.01 79.78 -70.77 ;
      LAYER V1 ;
        RECT 79.55 -71.03 79.75 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.52 -90.61 79.78 -90.37 ;
      LAYER V1 ;
        RECT 79.55 -90.55 79.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.48 -71.01 80.74 -70.77 ;
      LAYER M2 ;
        RECT 80.48 -71.01 80.74 -70.77 ;
      LAYER V1 ;
        RECT 80.51 -71.03 80.71 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.48 -90.61 80.74 -90.37 ;
      LAYER V1 ;
        RECT 80.51 -90.55 80.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.44 -71.01 81.7 -70.77 ;
      LAYER M2 ;
        RECT 81.44 -71.01 81.7 -70.77 ;
      LAYER V1 ;
        RECT 81.47 -71.03 81.67 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.44 -90.61 81.7 -90.37 ;
      LAYER V1 ;
        RECT 81.47 -90.55 81.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.4 -71.01 82.66 -70.77 ;
      LAYER M2 ;
        RECT 82.4 -71.01 82.66 -70.77 ;
      LAYER V1 ;
        RECT 82.43 -71.03 82.63 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.4 -90.61 82.66 -90.37 ;
      LAYER V1 ;
        RECT 82.43 -90.55 82.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.36 -71.01 83.62 -70.77 ;
      LAYER M2 ;
        RECT 83.36 -71.01 83.62 -70.77 ;
      LAYER V1 ;
        RECT 83.39 -71.03 83.59 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.36 -90.61 83.62 -90.37 ;
      LAYER V1 ;
        RECT 83.39 -90.55 83.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.32 -71.01 84.58 -70.77 ;
      LAYER M2 ;
        RECT 84.32 -71.01 84.58 -70.77 ;
      LAYER V1 ;
        RECT 84.35 -71.03 84.55 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.32 -90.61 84.58 -90.37 ;
      LAYER V1 ;
        RECT 84.35 -90.55 84.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.28 -71.01 85.54 -70.77 ;
      LAYER M2 ;
        RECT 85.28 -71.01 85.54 -70.77 ;
      LAYER V1 ;
        RECT 85.31 -71.03 85.51 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.28 -90.61 85.54 -90.37 ;
      LAYER V1 ;
        RECT 85.31 -90.55 85.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.24 -71.01 86.5 -70.77 ;
      LAYER M2 ;
        RECT 86.24 -71.01 86.5 -70.77 ;
      LAYER V1 ;
        RECT 86.27 -71.03 86.47 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.24 -90.61 86.5 -90.37 ;
      LAYER V1 ;
        RECT 86.27 -90.55 86.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.2 -71.01 87.46 -70.77 ;
      LAYER M2 ;
        RECT 87.2 -71.01 87.46 -70.77 ;
      LAYER V1 ;
        RECT 87.23 -71.03 87.43 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.2 -90.61 87.46 -90.37 ;
      LAYER V1 ;
        RECT 87.23 -90.55 87.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.16 -71.01 88.42 -70.77 ;
      LAYER M2 ;
        RECT 88.16 -71.01 88.42 -70.77 ;
      LAYER V1 ;
        RECT 88.19 -71.03 88.39 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.16 -90.61 88.42 -90.37 ;
      LAYER V1 ;
        RECT 88.19 -90.55 88.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.12 -71.01 89.38 -70.77 ;
      LAYER M2 ;
        RECT 89.12 -71.01 89.38 -70.77 ;
      LAYER V1 ;
        RECT 89.15 -71.03 89.35 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.12 -90.61 89.38 -90.37 ;
      LAYER V1 ;
        RECT 89.15 -90.55 89.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.08 -71.01 90.34 -70.77 ;
      LAYER M2 ;
        RECT 90.08 -71.01 90.34 -70.77 ;
      LAYER V1 ;
        RECT 90.11 -71.03 90.31 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.08 -90.61 90.34 -90.37 ;
      LAYER V1 ;
        RECT 90.11 -90.55 90.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.04 -71.01 91.3 -70.77 ;
      LAYER M2 ;
        RECT 91.04 -71.01 91.3 -70.77 ;
      LAYER V1 ;
        RECT 91.07 -71.03 91.27 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.04 -90.61 91.3 -90.37 ;
      LAYER V1 ;
        RECT 91.07 -90.55 91.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92 -71.01 92.26 -70.77 ;
      LAYER M2 ;
        RECT 92 -71.01 92.26 -70.77 ;
      LAYER V1 ;
        RECT 92.03 -71.03 92.23 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 92 -90.61 92.26 -90.37 ;
      LAYER V1 ;
        RECT 92.03 -90.55 92.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.96 -71.01 93.22 -70.77 ;
      LAYER M2 ;
        RECT 92.96 -71.01 93.22 -70.77 ;
      LAYER V1 ;
        RECT 92.99 -71.03 93.19 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.96 -90.61 93.22 -90.37 ;
      LAYER V1 ;
        RECT 92.99 -90.55 93.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.92 -71.01 94.18 -70.77 ;
      LAYER M2 ;
        RECT 93.92 -71.01 94.18 -70.77 ;
      LAYER V1 ;
        RECT 93.95 -71.03 94.15 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.92 -90.61 94.18 -90.37 ;
      LAYER V1 ;
        RECT 93.95 -90.55 94.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.88 -71.01 95.14 -70.77 ;
      LAYER M2 ;
        RECT 94.88 -71.01 95.14 -70.77 ;
      LAYER V1 ;
        RECT 94.91 -71.03 95.11 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.88 -90.61 95.14 -90.37 ;
      LAYER V1 ;
        RECT 94.91 -90.55 95.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.84 -71.01 96.1 -70.77 ;
      LAYER M2 ;
        RECT 95.84 -71.01 96.1 -70.77 ;
      LAYER V1 ;
        RECT 95.87 -71.03 96.07 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.84 -90.61 96.1 -90.37 ;
      LAYER V1 ;
        RECT 95.87 -90.55 96.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.8 -71.01 97.06 -70.77 ;
      LAYER M2 ;
        RECT 96.8 -71.01 97.06 -70.77 ;
      LAYER V1 ;
        RECT 96.83 -71.03 97.03 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.8 -90.61 97.06 -90.37 ;
      LAYER V1 ;
        RECT 96.83 -90.55 97.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.76 -71.01 98.02 -70.77 ;
      LAYER M2 ;
        RECT 97.76 -71.01 98.02 -70.77 ;
      LAYER V1 ;
        RECT 97.79 -71.03 97.99 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.76 -90.61 98.02 -90.37 ;
      LAYER V1 ;
        RECT 97.79 -90.55 97.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.72 -71.01 98.98 -70.77 ;
      LAYER M2 ;
        RECT 98.72 -71.01 98.98 -70.77 ;
      LAYER V1 ;
        RECT 98.75 -71.03 98.95 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.72 -90.61 98.98 -90.37 ;
      LAYER V1 ;
        RECT 98.75 -90.55 98.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.68 -71.01 99.94 -70.77 ;
      LAYER M2 ;
        RECT 99.68 -71.01 99.94 -70.77 ;
      LAYER V1 ;
        RECT 99.71 -71.03 99.91 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.68 -90.61 99.94 -90.37 ;
      LAYER V1 ;
        RECT 99.71 -90.55 99.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.64 -71.01 100.9 -70.77 ;
      LAYER M2 ;
        RECT 100.64 -71.01 100.9 -70.77 ;
      LAYER V1 ;
        RECT 100.67 -71.03 100.87 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.64 -90.61 100.9 -90.37 ;
      LAYER V1 ;
        RECT 100.67 -90.55 100.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.6 -71.01 101.86 -70.77 ;
      LAYER M2 ;
        RECT 101.6 -71.01 101.86 -70.77 ;
      LAYER V1 ;
        RECT 101.63 -71.03 101.83 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.6 -90.61 101.86 -90.37 ;
      LAYER V1 ;
        RECT 101.63 -90.55 101.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.56 -71.01 102.82 -70.77 ;
      LAYER M2 ;
        RECT 102.56 -71.01 102.82 -70.77 ;
      LAYER V1 ;
        RECT 102.59 -71.03 102.79 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.56 -90.61 102.82 -90.37 ;
      LAYER V1 ;
        RECT 102.59 -90.55 102.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.52 -71.01 103.78 -70.77 ;
      LAYER M2 ;
        RECT 103.52 -71.01 103.78 -70.77 ;
      LAYER V1 ;
        RECT 103.55 -71.03 103.75 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.52 -90.61 103.78 -90.37 ;
      LAYER V1 ;
        RECT 103.55 -90.55 103.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.48 -71.01 104.74 -70.77 ;
      LAYER M2 ;
        RECT 104.48 -71.01 104.74 -70.77 ;
      LAYER V1 ;
        RECT 104.51 -71.03 104.71 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.48 -90.61 104.74 -90.37 ;
      LAYER V1 ;
        RECT 104.51 -90.55 104.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.44 -71.01 105.7 -70.77 ;
      LAYER M2 ;
        RECT 105.44 -71.01 105.7 -70.77 ;
      LAYER V1 ;
        RECT 105.47 -71.03 105.67 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.44 -90.61 105.7 -90.37 ;
      LAYER V1 ;
        RECT 105.47 -90.55 105.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.4 -71.01 106.66 -70.77 ;
      LAYER M2 ;
        RECT 106.4 -71.01 106.66 -70.77 ;
      LAYER V1 ;
        RECT 106.43 -71.03 106.63 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.4 -90.61 106.66 -90.37 ;
      LAYER V1 ;
        RECT 106.43 -90.55 106.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.36 -71.01 107.62 -70.77 ;
      LAYER M2 ;
        RECT 107.36 -71.01 107.62 -70.77 ;
      LAYER V1 ;
        RECT 107.39 -71.03 107.59 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.36 -90.61 107.62 -90.37 ;
      LAYER V1 ;
        RECT 107.39 -90.55 107.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.32 -71.01 108.58 -70.77 ;
      LAYER M2 ;
        RECT 108.32 -71.01 108.58 -70.77 ;
      LAYER V1 ;
        RECT 108.35 -71.03 108.55 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.32 -90.61 108.58 -90.37 ;
      LAYER V1 ;
        RECT 108.35 -90.55 108.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.28 -71.01 109.54 -70.77 ;
      LAYER M2 ;
        RECT 109.28 -71.01 109.54 -70.77 ;
      LAYER V1 ;
        RECT 109.31 -71.03 109.51 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.28 -90.61 109.54 -90.37 ;
      LAYER V1 ;
        RECT 109.31 -90.55 109.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.24 -71.01 110.5 -70.77 ;
      LAYER M2 ;
        RECT 110.24 -71.01 110.5 -70.77 ;
      LAYER V1 ;
        RECT 110.27 -71.03 110.47 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.24 -90.61 110.5 -90.37 ;
      LAYER V1 ;
        RECT 110.27 -90.55 110.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.2 -71.01 111.46 -70.77 ;
      LAYER M2 ;
        RECT 111.2 -71.01 111.46 -70.77 ;
      LAYER V1 ;
        RECT 111.23 -71.03 111.43 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.2 -90.61 111.46 -90.37 ;
      LAYER V1 ;
        RECT 111.23 -90.55 111.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.16 -71.01 112.42 -70.77 ;
      LAYER M2 ;
        RECT 112.16 -71.01 112.42 -70.77 ;
      LAYER V1 ;
        RECT 112.19 -71.03 112.39 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.16 -90.61 112.42 -90.37 ;
      LAYER V1 ;
        RECT 112.19 -90.55 112.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.12 -71.01 113.38 -70.77 ;
      LAYER M2 ;
        RECT 113.12 -71.01 113.38 -70.77 ;
      LAYER V1 ;
        RECT 113.15 -71.03 113.35 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.12 -90.61 113.38 -90.37 ;
      LAYER V1 ;
        RECT 113.15 -90.55 113.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.08 -71.01 114.34 -70.77 ;
      LAYER M2 ;
        RECT 114.08 -71.01 114.34 -70.77 ;
      LAYER V1 ;
        RECT 114.11 -71.03 114.31 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.08 -90.61 114.34 -90.37 ;
      LAYER V1 ;
        RECT 114.11 -90.55 114.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.04 -71.01 115.3 -70.77 ;
      LAYER M2 ;
        RECT 115.04 -71.01 115.3 -70.77 ;
      LAYER V1 ;
        RECT 115.07 -71.03 115.27 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.04 -90.61 115.3 -90.37 ;
      LAYER V1 ;
        RECT 115.07 -90.55 115.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116 -71.01 116.26 -70.77 ;
      LAYER M2 ;
        RECT 116 -71.01 116.26 -70.77 ;
      LAYER V1 ;
        RECT 116.03 -71.03 116.23 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 116 -90.61 116.26 -90.37 ;
      LAYER V1 ;
        RECT 116.03 -90.55 116.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.96 -71.01 117.22 -70.77 ;
      LAYER M2 ;
        RECT 116.96 -71.01 117.22 -70.77 ;
      LAYER V1 ;
        RECT 116.99 -71.03 117.19 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.96 -90.61 117.22 -90.37 ;
      LAYER V1 ;
        RECT 116.99 -90.55 117.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.92 -71.01 118.18 -70.77 ;
      LAYER M2 ;
        RECT 117.92 -71.01 118.18 -70.77 ;
      LAYER V1 ;
        RECT 117.95 -71.03 118.15 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.92 -90.61 118.18 -90.37 ;
      LAYER V1 ;
        RECT 117.95 -90.55 118.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.88 -71.01 119.14 -70.77 ;
      LAYER M2 ;
        RECT 118.88 -71.01 119.14 -70.77 ;
      LAYER V1 ;
        RECT 118.91 -71.03 119.11 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.88 -90.61 119.14 -90.37 ;
      LAYER V1 ;
        RECT 118.91 -90.55 119.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.84 -71.01 120.1 -70.77 ;
      LAYER M2 ;
        RECT 119.84 -71.01 120.1 -70.77 ;
      LAYER V1 ;
        RECT 119.87 -71.03 120.07 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.84 -90.61 120.1 -90.37 ;
      LAYER V1 ;
        RECT 119.87 -90.55 120.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.8 -71.01 121.06 -70.77 ;
      LAYER M2 ;
        RECT 120.8 -71.01 121.06 -70.77 ;
      LAYER V1 ;
        RECT 120.83 -71.03 121.03 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.8 -90.61 121.06 -90.37 ;
      LAYER V1 ;
        RECT 120.83 -90.55 121.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.76 -71.01 122.02 -70.77 ;
      LAYER M2 ;
        RECT 121.76 -71.01 122.02 -70.77 ;
      LAYER V1 ;
        RECT 121.79 -71.03 121.99 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.76 -90.61 122.02 -90.37 ;
      LAYER V1 ;
        RECT 121.79 -90.55 121.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.72 -71.01 122.98 -70.77 ;
      LAYER M2 ;
        RECT 122.72 -71.01 122.98 -70.77 ;
      LAYER V1 ;
        RECT 122.75 -71.03 122.95 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.72 -90.61 122.98 -90.37 ;
      LAYER V1 ;
        RECT 122.75 -90.55 122.95 -90.35 ;
    END
  END DVDD
  PIN AVDD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 7.38 -61.17 9.38 -59.17 ;
      LAYER V1 ;
        RECT 7.38 -59.45 7.58 -59.25 ;
        RECT 7.38 -59.85 7.58 -59.65 ;
        RECT 7.38 -60.25 7.58 -60.05 ;
        RECT 7.38 -60.65 7.58 -60.45 ;
        RECT 7.38 -61.05 7.58 -60.85 ;
        RECT 7.78 -59.45 7.98 -59.25 ;
        RECT 7.78 -59.85 7.98 -59.65 ;
        RECT 7.78 -60.25 7.98 -60.05 ;
        RECT 7.78 -60.65 7.98 -60.45 ;
        RECT 7.78 -61.05 7.98 -60.85 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.1 -67.25 22.1 -65.25 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.55 -65.95 101.55 -50.95 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.9 -69.65 124.78 -68.77 ;
      LAYER V1 ;
        RECT 123.94 -69.09 124.14 -68.89 ;
        RECT 123.94 -69.53 124.14 -69.33 ;
        RECT 124.34 -69.09 124.54 -68.89 ;
        RECT 124.34 -69.53 124.54 -69.33 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.01 -60.63 4.17 -60.47 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.32 -61.91 8.04 -61.19 ;
      LAYER M2 ;
        RECT 7.38 -61.85 7.98 -61.25 ;
      LAYER V1 ;
        RECT 7.38 -61.45 7.58 -61.25 ;
        RECT 7.38 -61.85 7.58 -61.65 ;
        RECT 7.78 -61.45 7.98 -61.25 ;
        RECT 7.78 -61.85 7.98 -61.65 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -55.47 24.44 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -58.09 24.44 -57.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -62.67 24.44 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.98 -56.88 24.46 -56.4 ;
      LAYER M2 ;
        RECT 24.08 -57.14 24.68 -56.54 ;
      LAYER V1 ;
        RECT 24.08 -56.74 24.28 -56.54 ;
        RECT 24.48 -56.74 24.68 -56.54 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.98 -64.08 24.46 -63.6 ;
      LAYER M2 ;
        RECT 24.08 -63.94 24.68 -63.34 ;
      LAYER V1 ;
        RECT 24.08 -63.94 24.28 -63.74 ;
        RECT 24.48 -63.94 24.68 -63.74 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -55.47 25.4 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -58.09 25.4 -57.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -62.67 25.4 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.67 -69.21 25.93 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.86 -72.92 26.02 -72.76 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.79 -69.8 26.09 -69.5 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -55.47 26.36 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -55.89 26.36 -55.61 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -58.09 26.36 -57.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -62.67 26.36 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -63.09 26.36 -62.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -55.59 26.84 -55.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -57.98 26.84 -57.7 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -62.79 26.84 -62.5 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -55.59 27.8 -55.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -57.98 27.8 -57.7 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -62.79 27.8 -62.5 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.52 -72.92 28.68 -72.76 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.33 -69.42 28.8 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.12 -72.92 31.28 -72.76 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.05 -68.33 31.35 -68.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.05 -69.89 31.35 -69.59 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.05 -69.21 32.31 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.14 -68.35 36.46 -68.03 ;
      LAYER M2 ;
        RECT 36.13 -68.33 36.43 -68.03 ;
      LAYER V1 ;
        RECT 36.2 -68.29 36.4 -68.09 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.55 -68.35 36.87 -68.03 ;
      LAYER V1 ;
        RECT 36.6 -68.29 36.8 -68.09 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.57 -70.21 36.87 -69.91 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.64 -69.59 47.8 -69.43 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.57 -72.2 47.87 -71.9 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.57 -72.64 47.87 -72.34 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.38 -73.01 51.54 -72.85 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.31 -69.99 51.61 -69.69 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.31 -69.16 51.63 -68.84 ;
        RECT 51.19 -69.3 51.45 -69.04 ;
      LAYER M2 ;
        RECT 51.31 -69.55 51.61 -69.25 ;
      LAYER V1 ;
        RECT 51.37 -69.1 51.57 -68.9 ;
        RECT 51.37 -69.5 51.57 -69.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.8 -69.38 54.14 -69.04 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.99 -73.01 54.15 -72.85 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.92 -70.1 54.22 -69.8 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.44 -69.3 56.7 -69.04 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.63 -73.01 56.79 -72.85 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.57 -70.08 56.87 -69.78 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.56 -69.3 57.82 -69.04 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.32 -69.65 64.2 -68.77 ;
      LAYER M2 ;
        RECT 63.32 -69.65 64.2 -68.77 ;
      LAYER V1 ;
        RECT 63.54 -69.09 63.74 -68.89 ;
        RECT 63.54 -69.53 63.74 -69.33 ;
        RECT 63.94 -69.09 64.14 -68.89 ;
        RECT 63.94 -69.53 64.14 -69.33 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.32 -92.61 64.2 -91.73 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6 -71.03 65.86 -70.77 ;
      LAYER V1 ;
        RECT 65.63 -71.03 65.83 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6 -90.61 65.86 -90.35 ;
      LAYER M2 ;
        RECT 65.6 -90.61 65.86 -90.35 ;
      LAYER V1 ;
        RECT 65.63 -90.55 65.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.56 -71.03 66.82 -70.77 ;
      LAYER V1 ;
        RECT 66.59 -71.03 66.79 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.56 -90.61 66.82 -90.35 ;
      LAYER M2 ;
        RECT 66.56 -90.61 66.82 -90.35 ;
      LAYER V1 ;
        RECT 66.59 -90.55 66.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.52 -71.03 67.78 -70.77 ;
      LAYER V1 ;
        RECT 67.55 -71.03 67.75 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.52 -90.61 67.78 -90.35 ;
      LAYER M2 ;
        RECT 67.52 -90.61 67.78 -90.35 ;
      LAYER V1 ;
        RECT 67.55 -90.55 67.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.48 -71.03 68.74 -70.77 ;
      LAYER V1 ;
        RECT 68.51 -71.03 68.71 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.48 -90.61 68.74 -90.35 ;
      LAYER M2 ;
        RECT 68.48 -90.61 68.74 -90.35 ;
      LAYER V1 ;
        RECT 68.51 -90.55 68.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.44 -71.03 69.7 -70.77 ;
      LAYER V1 ;
        RECT 69.47 -71.03 69.67 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.44 -90.61 69.7 -90.35 ;
      LAYER M2 ;
        RECT 69.44 -90.61 69.7 -90.35 ;
      LAYER V1 ;
        RECT 69.47 -90.55 69.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4 -71.03 70.66 -70.77 ;
      LAYER V1 ;
        RECT 70.43 -71.03 70.63 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4 -90.61 70.66 -90.35 ;
      LAYER M2 ;
        RECT 70.4 -90.61 70.66 -90.35 ;
      LAYER V1 ;
        RECT 70.43 -90.55 70.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.36 -71.03 71.62 -70.77 ;
      LAYER V1 ;
        RECT 71.39 -71.03 71.59 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.36 -90.61 71.62 -90.35 ;
      LAYER M2 ;
        RECT 71.36 -90.61 71.62 -90.35 ;
      LAYER V1 ;
        RECT 71.39 -90.55 71.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.32 -71.03 72.58 -70.77 ;
      LAYER V1 ;
        RECT 72.35 -71.03 72.55 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.32 -90.61 72.58 -90.35 ;
      LAYER M2 ;
        RECT 72.32 -90.61 72.58 -90.35 ;
      LAYER V1 ;
        RECT 72.35 -90.55 72.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.28 -71.03 73.54 -70.77 ;
      LAYER V1 ;
        RECT 73.31 -71.03 73.51 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.28 -90.61 73.54 -90.35 ;
      LAYER M2 ;
        RECT 73.28 -90.61 73.54 -90.35 ;
      LAYER V1 ;
        RECT 73.31 -90.55 73.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.24 -71.03 74.5 -70.77 ;
      LAYER V1 ;
        RECT 74.27 -71.03 74.47 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.24 -90.61 74.5 -90.35 ;
      LAYER M2 ;
        RECT 74.24 -90.61 74.5 -90.35 ;
      LAYER V1 ;
        RECT 74.27 -90.55 74.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2 -71.03 75.46 -70.77 ;
      LAYER V1 ;
        RECT 75.23 -71.03 75.43 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2 -90.61 75.46 -90.35 ;
      LAYER M2 ;
        RECT 75.2 -90.61 75.46 -90.35 ;
      LAYER V1 ;
        RECT 75.23 -90.55 75.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.16 -71.03 76.42 -70.77 ;
      LAYER V1 ;
        RECT 76.19 -71.03 76.39 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.16 -90.61 76.42 -90.35 ;
      LAYER M2 ;
        RECT 76.16 -90.61 76.42 -90.35 ;
      LAYER V1 ;
        RECT 76.19 -90.55 76.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.12 -71.03 77.38 -70.77 ;
      LAYER V1 ;
        RECT 77.15 -71.03 77.35 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.12 -90.61 77.38 -90.35 ;
      LAYER M2 ;
        RECT 77.12 -90.61 77.38 -90.35 ;
      LAYER V1 ;
        RECT 77.15 -90.55 77.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.08 -71.03 78.34 -70.77 ;
      LAYER V1 ;
        RECT 78.11 -71.03 78.31 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.08 -90.61 78.34 -90.35 ;
      LAYER M2 ;
        RECT 78.08 -90.61 78.34 -90.35 ;
      LAYER V1 ;
        RECT 78.11 -90.55 78.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.04 -71.03 79.3 -70.77 ;
      LAYER V1 ;
        RECT 79.07 -71.03 79.27 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.04 -90.61 79.3 -90.35 ;
      LAYER M2 ;
        RECT 79.04 -90.61 79.3 -90.35 ;
      LAYER V1 ;
        RECT 79.07 -90.55 79.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80 -71.03 80.26 -70.77 ;
      LAYER V1 ;
        RECT 80.03 -71.03 80.23 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 80 -90.61 80.26 -90.35 ;
      LAYER M2 ;
        RECT 80 -90.61 80.26 -90.35 ;
      LAYER V1 ;
        RECT 80.03 -90.55 80.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.96 -71.03 81.22 -70.77 ;
      LAYER V1 ;
        RECT 80.99 -71.03 81.19 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.96 -90.61 81.22 -90.35 ;
      LAYER M2 ;
        RECT 80.96 -90.61 81.22 -90.35 ;
      LAYER V1 ;
        RECT 80.99 -90.55 81.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.92 -71.03 82.18 -70.77 ;
      LAYER V1 ;
        RECT 81.95 -71.03 82.15 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.92 -90.61 82.18 -90.35 ;
      LAYER M2 ;
        RECT 81.92 -90.61 82.18 -90.35 ;
      LAYER V1 ;
        RECT 81.95 -90.55 82.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.88 -71.03 83.14 -70.77 ;
      LAYER V1 ;
        RECT 82.91 -71.03 83.11 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.88 -90.61 83.14 -90.35 ;
      LAYER M2 ;
        RECT 82.88 -90.61 83.14 -90.35 ;
      LAYER V1 ;
        RECT 82.91 -90.55 83.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.84 -71.03 84.1 -70.77 ;
      LAYER V1 ;
        RECT 83.87 -71.03 84.07 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.84 -90.61 84.1 -90.35 ;
      LAYER M2 ;
        RECT 83.84 -90.61 84.1 -90.35 ;
      LAYER V1 ;
        RECT 83.87 -90.55 84.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8 -71.03 85.06 -70.77 ;
      LAYER V1 ;
        RECT 84.83 -71.03 85.03 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8 -90.61 85.06 -90.35 ;
      LAYER M2 ;
        RECT 84.8 -90.61 85.06 -90.35 ;
      LAYER V1 ;
        RECT 84.83 -90.55 85.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.76 -71.03 86.02 -70.77 ;
      LAYER V1 ;
        RECT 85.79 -71.03 85.99 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.76 -90.61 86.02 -90.35 ;
      LAYER M2 ;
        RECT 85.76 -90.61 86.02 -90.35 ;
      LAYER V1 ;
        RECT 85.79 -90.55 85.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.72 -71.03 86.98 -70.77 ;
      LAYER V1 ;
        RECT 86.75 -71.03 86.95 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.72 -90.61 86.98 -90.35 ;
      LAYER M2 ;
        RECT 86.72 -90.61 86.98 -90.35 ;
      LAYER V1 ;
        RECT 86.75 -90.55 86.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.68 -71.03 87.94 -70.77 ;
      LAYER V1 ;
        RECT 87.71 -71.03 87.91 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.68 -90.61 87.94 -90.35 ;
      LAYER M2 ;
        RECT 87.68 -90.61 87.94 -90.35 ;
      LAYER V1 ;
        RECT 87.71 -90.55 87.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.64 -71.03 88.9 -70.77 ;
      LAYER V1 ;
        RECT 88.67 -71.03 88.87 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.64 -90.61 88.9 -90.35 ;
      LAYER M2 ;
        RECT 88.64 -90.61 88.9 -90.35 ;
      LAYER V1 ;
        RECT 88.67 -90.55 88.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.6 -71.03 89.86 -70.77 ;
      LAYER V1 ;
        RECT 89.63 -71.03 89.83 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.6 -90.61 89.86 -90.35 ;
      LAYER M2 ;
        RECT 89.6 -90.61 89.86 -90.35 ;
      LAYER V1 ;
        RECT 89.63 -90.55 89.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.56 -71.03 90.82 -70.77 ;
      LAYER V1 ;
        RECT 90.59 -71.03 90.79 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.56 -90.61 90.82 -90.35 ;
      LAYER M2 ;
        RECT 90.56 -90.61 90.82 -90.35 ;
      LAYER V1 ;
        RECT 90.59 -90.55 90.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.52 -71.03 91.78 -70.77 ;
      LAYER V1 ;
        RECT 91.55 -71.03 91.75 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.52 -90.61 91.78 -90.35 ;
      LAYER M2 ;
        RECT 91.52 -90.61 91.78 -90.35 ;
      LAYER V1 ;
        RECT 91.55 -90.55 91.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.48 -71.03 92.74 -70.77 ;
      LAYER V1 ;
        RECT 92.51 -71.03 92.71 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.48 -90.61 92.74 -90.35 ;
      LAYER M2 ;
        RECT 92.48 -90.61 92.74 -90.35 ;
      LAYER V1 ;
        RECT 92.51 -90.55 92.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.44 -71.03 93.7 -70.77 ;
      LAYER V1 ;
        RECT 93.47 -71.03 93.67 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.44 -90.61 93.7 -90.35 ;
      LAYER M2 ;
        RECT 93.44 -90.61 93.7 -90.35 ;
      LAYER V1 ;
        RECT 93.47 -90.55 93.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4 -71.03 94.66 -70.77 ;
      LAYER V1 ;
        RECT 94.43 -71.03 94.63 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4 -90.61 94.66 -90.35 ;
      LAYER M2 ;
        RECT 94.4 -90.61 94.66 -90.35 ;
      LAYER V1 ;
        RECT 94.43 -90.55 94.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.36 -71.03 95.62 -70.77 ;
      LAYER V1 ;
        RECT 95.39 -71.03 95.59 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.36 -90.61 95.62 -90.35 ;
      LAYER M2 ;
        RECT 95.36 -90.61 95.62 -90.35 ;
      LAYER V1 ;
        RECT 95.39 -90.55 95.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.32 -71.03 96.58 -70.77 ;
      LAYER V1 ;
        RECT 96.35 -71.03 96.55 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.32 -90.61 96.58 -90.35 ;
      LAYER M2 ;
        RECT 96.32 -90.61 96.58 -90.35 ;
      LAYER V1 ;
        RECT 96.35 -90.55 96.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.28 -71.03 97.54 -70.77 ;
      LAYER V1 ;
        RECT 97.31 -71.03 97.51 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.28 -90.61 97.54 -90.35 ;
      LAYER M2 ;
        RECT 97.28 -90.61 97.54 -90.35 ;
      LAYER V1 ;
        RECT 97.31 -90.55 97.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.24 -71.03 98.5 -70.77 ;
      LAYER V1 ;
        RECT 98.27 -71.03 98.47 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.24 -90.61 98.5 -90.35 ;
      LAYER M2 ;
        RECT 98.24 -90.61 98.5 -90.35 ;
      LAYER V1 ;
        RECT 98.27 -90.55 98.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.2 -71.03 99.46 -70.77 ;
      LAYER V1 ;
        RECT 99.23 -71.03 99.43 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.2 -90.61 99.46 -90.35 ;
      LAYER M2 ;
        RECT 99.2 -90.61 99.46 -90.35 ;
      LAYER V1 ;
        RECT 99.23 -90.55 99.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.16 -71.03 100.42 -70.77 ;
      LAYER V1 ;
        RECT 100.19 -71.03 100.39 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.16 -90.61 100.42 -90.35 ;
      LAYER M2 ;
        RECT 100.16 -90.61 100.42 -90.35 ;
      LAYER V1 ;
        RECT 100.19 -90.55 100.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.12 -71.03 101.38 -70.77 ;
      LAYER V1 ;
        RECT 101.15 -71.03 101.35 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.12 -90.61 101.38 -90.35 ;
      LAYER M2 ;
        RECT 101.12 -90.61 101.38 -90.35 ;
      LAYER V1 ;
        RECT 101.15 -90.55 101.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.08 -71.03 102.34 -70.77 ;
      LAYER V1 ;
        RECT 102.11 -71.03 102.31 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.08 -90.61 102.34 -90.35 ;
      LAYER M2 ;
        RECT 102.08 -90.61 102.34 -90.35 ;
      LAYER V1 ;
        RECT 102.11 -90.55 102.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.04 -71.03 103.3 -70.77 ;
      LAYER V1 ;
        RECT 103.07 -71.03 103.27 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.04 -90.61 103.3 -90.35 ;
      LAYER M2 ;
        RECT 103.04 -90.61 103.3 -90.35 ;
      LAYER V1 ;
        RECT 103.07 -90.55 103.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104 -71.03 104.26 -70.77 ;
      LAYER V1 ;
        RECT 104.03 -71.03 104.23 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 104 -90.61 104.26 -90.35 ;
      LAYER M2 ;
        RECT 104 -90.61 104.26 -90.35 ;
      LAYER V1 ;
        RECT 104.03 -90.55 104.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.96 -71.03 105.22 -70.77 ;
      LAYER V1 ;
        RECT 104.99 -71.03 105.19 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.96 -90.61 105.22 -90.35 ;
      LAYER M2 ;
        RECT 104.96 -90.61 105.22 -90.35 ;
      LAYER V1 ;
        RECT 104.99 -90.55 105.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.92 -71.03 106.18 -70.77 ;
      LAYER V1 ;
        RECT 105.95 -71.03 106.15 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.92 -90.61 106.18 -90.35 ;
      LAYER M2 ;
        RECT 105.92 -90.61 106.18 -90.35 ;
      LAYER V1 ;
        RECT 105.95 -90.55 106.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.88 -71.03 107.14 -70.77 ;
      LAYER V1 ;
        RECT 106.91 -71.03 107.11 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.88 -90.61 107.14 -90.35 ;
      LAYER M2 ;
        RECT 106.88 -90.61 107.14 -90.35 ;
      LAYER V1 ;
        RECT 106.91 -90.55 107.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.84 -71.03 108.1 -70.77 ;
      LAYER V1 ;
        RECT 107.87 -71.03 108.07 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.84 -90.61 108.1 -90.35 ;
      LAYER M2 ;
        RECT 107.84 -90.61 108.1 -90.35 ;
      LAYER V1 ;
        RECT 107.87 -90.55 108.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.8 -71.03 109.06 -70.77 ;
      LAYER V1 ;
        RECT 108.83 -71.03 109.03 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.8 -90.61 109.06 -90.35 ;
      LAYER M2 ;
        RECT 108.8 -90.61 109.06 -90.35 ;
      LAYER V1 ;
        RECT 108.83 -90.55 109.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.76 -71.03 110.02 -70.77 ;
      LAYER V1 ;
        RECT 109.79 -71.03 109.99 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.76 -90.61 110.02 -90.35 ;
      LAYER M2 ;
        RECT 109.76 -90.61 110.02 -90.35 ;
      LAYER V1 ;
        RECT 109.79 -90.55 109.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.72 -71.03 110.98 -70.77 ;
      LAYER V1 ;
        RECT 110.75 -71.03 110.95 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.72 -90.61 110.98 -90.35 ;
      LAYER M2 ;
        RECT 110.72 -90.61 110.98 -90.35 ;
      LAYER V1 ;
        RECT 110.75 -90.55 110.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.68 -71.03 111.94 -70.77 ;
      LAYER V1 ;
        RECT 111.71 -71.03 111.91 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.68 -90.61 111.94 -90.35 ;
      LAYER M2 ;
        RECT 111.68 -90.61 111.94 -90.35 ;
      LAYER V1 ;
        RECT 111.71 -90.55 111.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.64 -71.03 112.9 -70.77 ;
      LAYER V1 ;
        RECT 112.67 -71.03 112.87 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.64 -90.61 112.9 -90.35 ;
      LAYER M2 ;
        RECT 112.64 -90.61 112.9 -90.35 ;
      LAYER V1 ;
        RECT 112.67 -90.55 112.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.6 -71.03 113.86 -70.77 ;
      LAYER V1 ;
        RECT 113.63 -71.03 113.83 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.6 -90.61 113.86 -90.35 ;
      LAYER M2 ;
        RECT 113.6 -90.61 113.86 -90.35 ;
      LAYER V1 ;
        RECT 113.63 -90.55 113.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.56 -71.03 114.82 -70.77 ;
      LAYER V1 ;
        RECT 114.59 -71.03 114.79 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.56 -90.61 114.82 -90.35 ;
      LAYER M2 ;
        RECT 114.56 -90.61 114.82 -90.35 ;
      LAYER V1 ;
        RECT 114.59 -90.55 114.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.52 -71.03 115.78 -70.77 ;
      LAYER V1 ;
        RECT 115.55 -71.03 115.75 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.52 -90.61 115.78 -90.35 ;
      LAYER M2 ;
        RECT 115.52 -90.61 115.78 -90.35 ;
      LAYER V1 ;
        RECT 115.55 -90.55 115.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.48 -71.03 116.74 -70.77 ;
      LAYER V1 ;
        RECT 116.51 -71.03 116.71 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.48 -90.61 116.74 -90.35 ;
      LAYER M2 ;
        RECT 116.48 -90.61 116.74 -90.35 ;
      LAYER V1 ;
        RECT 116.51 -90.55 116.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.44 -71.03 117.7 -70.77 ;
      LAYER V1 ;
        RECT 117.47 -71.03 117.67 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.44 -90.61 117.7 -90.35 ;
      LAYER M2 ;
        RECT 117.44 -90.61 117.7 -90.35 ;
      LAYER V1 ;
        RECT 117.47 -90.55 117.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.4 -71.03 118.66 -70.77 ;
      LAYER V1 ;
        RECT 118.43 -71.03 118.63 -70.83 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.4 -90.61 118.66 -90.35 ;
      LAYER M2 ;
        RECT 118.4 -90.61 118.66 -90.35 ;
      LAYER V1 ;
        RECT 118.43 -90.55 118.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.36 -90.61 119.62 -90.35 ;
      LAYER M2 ;
        RECT 119.36 -90.61 119.62 -90.35 ;
      LAYER V1 ;
        RECT 119.39 -90.55 119.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.32 -90.61 120.58 -90.35 ;
      LAYER M2 ;
        RECT 120.32 -90.61 120.58 -90.35 ;
      LAYER V1 ;
        RECT 120.35 -90.55 120.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.28 -90.61 121.54 -90.35 ;
      LAYER M2 ;
        RECT 121.28 -90.61 121.54 -90.35 ;
      LAYER V1 ;
        RECT 121.31 -90.55 121.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.24 -90.61 122.5 -90.35 ;
      LAYER M2 ;
        RECT 122.24 -90.61 122.5 -90.35 ;
      LAYER V1 ;
        RECT 122.27 -90.55 122.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.34 -92.61 124.78 -92.17 ;
    END
  END AVDD
  PIN AVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 38.8 -69 38.98 -68.8 ;
      LAYER V2 ;
        RECT 38.78 -69 38.98 -68.8 ;
      LAYER V1 ;
        RECT 38.78 -69 38.98 -68.8 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER M3 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER M4 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER V3 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
      LAYER V2 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
      LAYER V1 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER M3 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER M4 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER V3 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
      LAYER V2 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
      LAYER V1 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.28 -53.12 27.88 -52.54 ;
      LAYER V1 ;
        RECT 27.28 -52.74 27.48 -52.54 ;
        RECT 27.28 -53.14 27.48 -52.94 ;
        RECT 27.68 -52.74 27.88 -52.54 ;
        RECT 27.68 -53.14 27.88 -52.94 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.28 -60.34 27.88 -59.76 ;
      LAYER V1 ;
        RECT 27.28 -60.34 27.48 -60.14 ;
        RECT 27.68 -60.34 27.88 -60.14 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.22 -90.74 38.82 -90.14 ;
      LAYER M3 ;
        RECT 38.22 -90.74 38.82 -90.14 ;
        RECT 38.52 -90.8 38.82 -90.14 ;
      LAYER V2 ;
        RECT 38.22 -90.34 38.42 -90.14 ;
        RECT 38.22 -90.74 38.42 -90.54 ;
        RECT 38.62 -90.34 38.82 -90.14 ;
        RECT 38.62 -90.74 38.82 -90.54 ;
      LAYER V1 ;
        RECT 38.22 -90.34 38.42 -90.14 ;
        RECT 38.22 -90.74 38.42 -90.54 ;
        RECT 38.62 -90.34 38.82 -90.14 ;
        RECT 38.62 -90.74 38.82 -90.54 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.16 -92.22 3.4 -91.98 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.01 -68.27 4.15 -68.11 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.72 -63.63 9.98 -63.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.72 -69.75 9.98 -69.51 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.87 -69.23 22.99 -68.11 ;
      LAYER M2 ;
        RECT 21.93 -69.17 22.93 -68.17 ;
      LAYER M3 ;
        RECT 21.93 -69.17 22.93 -68.17 ;
      LAYER M4 ;
        RECT 21.93 -69.17 22.91 -68.17 ;
      LAYER V3 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
      LAYER V2 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
      LAYER V1 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -54.25 24.44 -53.99 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -59.29 24.44 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.98 -60.48 24.44 -60 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -61.45 24.44 -61.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -54.25 25.4 -53.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -59.32 25.4 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -61.45 25.4 -61.16 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -54.25 26.36 -53.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -59.32 26.36 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -61.45 26.36 -61.16 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -54.25 26.84 -53.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -59.32 26.84 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -61.45 26.84 -61.16 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -54.25 27.8 -53.96 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -59.32 27.8 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -61.45 27.8 -61.16 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.92 -60.48 32.38 -60 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.16 -87.14 36.32 -87 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.32 -69.06 38.62 -68.74 ;
      LAYER M2 ;
        RECT 38.38 -69 38.56 -68.8 ;
      LAYER M3 ;
        RECT 38.38 -69 38.56 -68.8 ;
      LAYER V2 ;
        RECT 38.38 -69 38.58 -68.8 ;
      LAYER V1 ;
        RECT 38.38 -69 38.58 -68.8 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.61 -87.14 38.77 -87 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.75 -66.65 39.93 -66.45 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.15 -87.13 43.31 -86.99 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.49 -66.65 43.67 -66.45 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.75 -69.06 44.05 -68.74 ;
      LAYER M2 ;
        RECT 43.81 -69 43.99 -68.8 ;
      LAYER V1 ;
        RECT 43.79 -69 43.99 -68.8 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.6 -87.45 45.76 -86.99 ;
        RECT 45.54 -87.45 45.76 -87.05 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.54 -88.87 45.76 -88.47 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.84 -92.77 46.82 -90.77 ;
        RECT 44.84 -92.77 45.21 -90.58 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.03 -62.45 50.41 -62.05 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.18 -52.94 51.16 -50.94 ;
        RECT 49.18 -52.99 50.43 -50.94 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.82 -77.96 59.94 -76.84 ;
      LAYER M2 ;
        RECT 58.88 -77.9 59.88 -76.9 ;
      LAYER M3 ;
        RECT 58.88 -77.9 59.88 -76.9 ;
      LAYER M4 ;
        RECT 58.88 -77.9 59.88 -76.92 ;
      LAYER V3 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
      LAYER V2 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
      LAYER V1 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
    END
  END AVSS
  OBS
    LAYER M1 ;
      RECT 66.12 -69.65 124.78 -68.77 ;
      RECT 124.34 -90.25 124.78 -68.77 ;
      RECT 64.32 -70.61 124 -70.03 ;
      RECT 123.38 -91.33 124 -70.03 ;
      RECT 64.32 -91.33 64.72 -70.03 ;
      RECT 64.32 -91.33 124 -90.77 ;
      RECT -0.34 -52.04 47.26 -50.94 ;
      RECT 29.72 -52.99 47.26 -50.94 ;
      RECT -0.34 -52.07 23.2 -50.94 ;
      RECT -0.34 -52.94 22.24 -50.94 ;
      RECT -0.34 -96.32 1.66 -50.94 ;
      RECT 29.72 -53.28 32.38 -50.94 ;
      RECT 11.9 -93.67 19.95 -68.11 ;
      RECT 11.9 -93.67 21.57 -71.15 ;
      RECT 11.21 -93.67 21.57 -71.67 ;
      RECT 38.61 -92.77 38.77 -89.06 ;
      RECT 36.16 -92.77 36.32 -89.06 ;
      RECT 38.16 -92.77 38.88 -90.08 ;
      RECT 36.09 -92.77 36.39 -90.21 ;
      RECT 36.09 -92.77 42.92 -90.52 ;
      RECT 33.94 -92.77 42.92 -90.77 ;
      RECT 33.94 -96.32 35.94 -90.77 ;
      RECT 14.61 -96.32 14.85 -68.11 ;
      RECT 11.22 -96.32 11.46 -71.67 ;
      RECT 5.32 -96.32 14.85 -94.13 ;
      RECT 3.16 -96.32 14.85 -94.14 ;
      RECT -0.34 -96.32 35.94 -94.32 ;
      RECT 9.72 -66.39 9.98 -65.55 ;
      RECT 9.82 -67.59 9.98 -65.55 ;
      RECT 66.12 -92.61 122.42 -91.73 ;
      RECT 50.75 -60.13 51.15 -54.91 ;
      RECT 5.32 -93.03 9.21 -92.87 ;
      RECT 6.07 -68.27 7.8 -68.11 ;
    LAYER M1 SPACING 0.16 ;
      RECT -0.34 -50.62 125.11 -48.96 ;
      RECT 123.3 -91.85 125.11 -48.96 ;
      RECT 51.48 -68.45 125.11 -48.96 ;
      RECT 64.52 -70.61 125.11 -48.96 ;
      RECT -0.34 -53.46 48.86 -48.96 ;
      RECT 50.75 -68.52 63 -53.26 ;
      RECT 50.73 -96.81 50.87 -53.31 ;
      RECT 35.06 -61.73 125.11 -53.31 ;
      RECT -0.34 -53.64 34.08 -48.96 ;
      RECT 28.12 -53.72 34.08 -48.96 ;
      RECT 32.7 -70.71 34.08 -48.96 ;
      RECT -0.34 -53.67 24.8 -48.96 ;
      RECT -0.34 -54.03 23.84 -48.96 ;
      RECT 22.2 -56.08 23.84 -48.96 ;
      RECT 31.96 -54.81 34.08 -48.96 ;
      RECT 31.99 -59.68 34.08 -48.96 ;
      RECT 31 -54.29 31.16 -48.96 ;
      RECT 30.04 -54.29 30.2 -48.96 ;
      RECT 29.08 -54.29 29.24 -48.96 ;
      RECT 28.12 -54.29 28.28 -48.96 ;
      RECT 27.04 -54.25 27.33 -53.96 ;
      RECT 27.16 -55.48 27.33 -53.96 ;
      RECT 25.6 -54.25 25.89 -53.96 ;
      RECT 25.72 -55.89 25.89 -53.96 ;
      RECT 24.64 -54.25 24.92 -53.96 ;
      RECT 31.84 -54.29 34.08 -54 ;
      RECT 30.88 -54.29 31.16 -54 ;
      RECT 29.92 -54.29 30.2 -54 ;
      RECT 28.96 -54.29 29.24 -54 ;
      RECT 28 -54.29 28.28 -54 ;
      RECT -0.34 -60.15 20.84 -48.96 ;
      RECT 24.76 -56.08 24.92 -53.96 ;
      RECT 33.57 -96.81 35.82 -54.38 ;
      RECT 24.76 -54.87 28.16 -54.57 ;
      RECT 22.2 -54.87 24.12 -54.57 ;
      RECT 31.95 -54.81 125.11 -54.58 ;
      RECT 24.76 -54.81 125.11 -54.61 ;
      RECT 28.12 -55.17 31.21 -54.61 ;
      RECT 26.68 -54.98 31.21 -54.61 ;
      RECT 27.16 -55.12 28.16 -54.57 ;
      RECT 28.12 -55.29 28.42 -54.61 ;
      RECT 25.6 -58.09 25.76 -55.19 ;
      RECT 24.64 -56.08 24.92 -55.19 ;
      RECT 27.04 -55.59 27.32 -55.3 ;
      RECT -0.34 -57.74 23.66 -55.39 ;
      RECT 31.88 -55.78 125.11 -55.49 ;
      RECT 30.9 -55.78 31.18 -55.49 ;
      RECT 31.02 -67.71 31.18 -55.49 ;
      RECT 29.94 -55.78 30.22 -55.49 ;
      RECT 30.05 -96.81 30.22 -55.49 ;
      RECT 28.96 -55.78 29.24 -55.49 ;
      RECT 28 -57.79 28.28 -55.49 ;
      RECT 29.08 -68.63 29.24 -55.49 ;
      RECT 24.78 -57.49 25.76 -55.79 ;
      RECT -0.34 -56.08 25.76 -55.79 ;
      RECT 26.57 -57.38 28.28 -55.91 ;
      RECT 28.12 -59.72 32.12 -56 ;
      RECT 24.78 -57.38 125.11 -56.21 ;
      RECT 24.76 -59.32 24.92 -57.2 ;
      RECT -0.34 -57.49 26.36 -57.2 ;
      RECT 25.72 -59.32 25.89 -56.21 ;
      RECT 24.64 -58.09 24.92 -57.2 ;
      RECT 22.97 -59.68 23.84 -57.2 ;
      RECT 27.04 -57.98 27.32 -57.69 ;
      RECT -0.34 -60.15 21.61 -55.39 ;
      RECT 27.16 -59.32 27.33 -57.8 ;
      RECT 27.16 -58.71 125.11 -58.16 ;
      RECT 26.68 -58.71 125.11 -58.3 ;
      RECT 24.76 -58.71 125.11 -58.41 ;
      RECT 22.97 -58.71 24.12 -58.41 ;
      RECT 28 -59.28 125.11 -58.99 ;
      RECT 27.04 -59.32 27.33 -59.03 ;
      RECT 25.6 -59.32 25.89 -59.03 ;
      RECT 24.64 -59.32 24.92 -59.03 ;
      RECT 24.76 -60.84 31.6 -59.64 ;
      RECT 4.49 -60.87 23.66 -59.1 ;
      RECT -0.34 -91.66 3.69 -48.96 ;
      RECT 24.76 -60.84 32.12 -60.76 ;
      RECT 8.36 -61.41 23.84 -60.8 ;
      RECT 31.67 -68.63 35.82 -60.8 ;
      RECT 4.49 -96.81 7 -48.96 ;
      RECT -0.34 -67.79 7 -60.95 ;
      RECT 27.04 -61.45 27.33 -61.16 ;
      RECT 27.16 -62.68 27.33 -61.16 ;
      RECT 25.6 -61.45 25.89 -61.16 ;
      RECT 25.72 -63.09 25.89 -61.16 ;
      RECT 24.64 -61.45 24.92 -61.16 ;
      RECT 28 -61.49 125.11 -61.2 ;
      RECT 8.36 -63.07 22.36 -59.1 ;
      RECT 24.76 -63.28 24.92 -61.16 ;
      RECT -0.34 -61.67 7.01 -61.51 ;
      RECT 28.12 -66.13 49.71 -60.8 ;
      RECT 24.76 -62.07 49.71 -61.77 ;
      RECT 27.16 -62.32 49.71 -61.77 ;
      RECT 26.68 -62.18 49.71 -61.77 ;
      RECT 4.47 -96.81 9.4 -62.23 ;
      RECT 25.6 -63.09 25.89 -62.39 ;
      RECT 24.64 -63.28 24.92 -62.39 ;
      RECT 27.04 -62.79 27.32 -62.5 ;
      RECT 28 -66.13 49.71 -62.69 ;
      RECT -0.34 -63.07 23.84 -62.77 ;
      RECT 24.78 -68.63 25.76 -62.99 ;
      RECT 10.3 -63.28 25.76 -62.99 ;
      RECT 26.57 -66.13 125.11 -63.11 ;
      RECT 10.3 -67.79 23.66 -62.77 ;
      RECT 24.78 -66.13 125.11 -63.41 ;
      RECT 26.41 -96.81 28.01 -63.41 ;
      RECT 4.47 -69.19 21.55 -63.95 ;
      RECT 23.31 -96.81 25.35 -64.4 ;
      RECT 43.99 -68.21 125.11 -62.77 ;
      RECT 50.64 -71.08 50.87 -62.77 ;
      RECT 40.25 -86.67 43.17 -48.96 ;
      RECT -0.34 -67.71 39.43 -64.4 ;
      RECT 37.19 -68.42 46.48 -66.97 ;
      RECT 26.25 -69.18 28.01 -63.41 ;
      RECT 23.31 -68.63 30.73 -64.4 ;
      RECT 47.36 -69.11 49.76 -62.77 ;
      RECT 44.37 -86.67 46.48 -48.96 ;
      RECT 38.94 -86.67 43.43 -66.97 ;
      RECT 37.19 -96.81 38 -48.96 ;
      RECT 32.63 -69.59 36.38 -68.52 ;
      RECT 51.95 -68.72 63 -48.96 ;
      RECT 50.64 -68.72 50.99 -62.77 ;
      RECT 29.12 -96.81 30.73 -56 ;
      RECT 29.12 -69.27 31.73 -68.65 ;
      RECT 32.63 -69.59 38 -68.67 ;
      RECT 58.14 -76.52 63 -48.96 ;
      RECT 57.02 -69.46 57.24 -48.96 ;
      RECT 54.46 -69.48 56.12 -48.96 ;
      RECT 54.54 -96.81 56.12 -48.96 ;
      RECT 51.95 -96.81 53.48 -48.96 ;
      RECT 48.12 -71.08 50.87 -69.09 ;
      RECT 44.37 -69.75 47.32 -69.09 ;
      RECT 10.3 -96.81 21.55 -55.39 ;
      RECT -0.34 -91.66 9.4 -68.59 ;
      RECT 51.93 -96.81 53.48 -69.48 ;
      RECT 31.67 -70.71 36.25 -69.53 ;
      RECT 23.31 -96.81 25.47 -69.53 ;
      RECT 10.3 -96.81 25.47 -69.55 ;
      RECT 37.19 -86.67 46.48 -69.38 ;
      RECT 57.19 -76.52 63 -69.62 ;
      RECT 54.54 -96.81 56.25 -69.62 ;
      RECT 48.12 -71.08 50.99 -69.62 ;
      RECT 51.93 -96.81 53.6 -69.7 ;
      RECT 26.41 -72.44 30.73 -69.74 ;
      RECT 47.28 -71.08 50.99 -69.91 ;
      RECT 60.26 -91.41 64.8 -69.97 ;
      RECT -0.34 -91.66 25.47 -70.07 ;
      RECT -0.34 -72.44 30.73 -70.12 ;
      RECT 26.34 -96.81 28.2 -70.12 ;
      RECT 47.28 -71.08 53.6 -70.31 ;
      RECT 54.54 -70.61 125.11 -70.4 ;
      RECT 57.11 -96.81 58.5 -70.4 ;
      RECT 54.47 -96.81 56.31 -70.42 ;
      RECT -0.34 -70.71 46.48 -70.53 ;
      RECT 36.64 -96.81 38.29 -70.53 ;
      RECT 33.57 -71.58 49.72 -70.55 ;
      RECT 50.68 -72.53 64.8 -70.42 ;
      RECT -0.34 -72.44 32.61 -70.21 ;
      RECT 122.24 -90.03 122.5 -70.77 ;
      RECT 121.28 -90.03 121.54 -70.77 ;
      RECT 120.32 -90.03 120.58 -70.77 ;
      RECT 119.36 -90.03 119.62 -70.77 ;
      RECT 118.88 -90.03 125.11 -71.33 ;
      RECT 122.72 -90.05 125.11 -71.33 ;
      RECT 117.92 -90.05 118.18 -71.33 ;
      RECT 116.96 -90.05 117.22 -71.33 ;
      RECT 116 -90.05 116.26 -71.33 ;
      RECT 115.04 -90.05 115.3 -71.33 ;
      RECT 114.08 -90.05 114.34 -71.33 ;
      RECT 113.12 -90.05 113.38 -71.33 ;
      RECT 112.16 -90.05 112.42 -71.33 ;
      RECT 111.2 -90.05 111.46 -71.33 ;
      RECT 110.24 -90.05 110.5 -71.33 ;
      RECT 109.28 -90.05 109.54 -71.33 ;
      RECT 108.32 -90.05 108.58 -71.33 ;
      RECT 107.36 -90.05 107.62 -71.33 ;
      RECT 106.4 -90.05 106.66 -71.33 ;
      RECT 105.44 -90.05 105.7 -71.33 ;
      RECT 104.48 -90.05 104.74 -71.33 ;
      RECT 103.52 -90.05 103.78 -71.33 ;
      RECT 102.56 -90.05 102.82 -71.33 ;
      RECT 101.6 -90.05 101.86 -71.33 ;
      RECT 100.64 -90.05 100.9 -71.33 ;
      RECT 99.68 -90.05 99.94 -71.33 ;
      RECT 98.72 -90.05 98.98 -71.33 ;
      RECT 97.76 -90.05 98.02 -71.33 ;
      RECT 96.8 -90.05 97.06 -71.33 ;
      RECT 95.84 -90.05 96.1 -71.33 ;
      RECT 94.88 -90.05 95.14 -71.33 ;
      RECT 93.92 -90.05 94.18 -71.33 ;
      RECT 92.96 -90.05 93.22 -71.33 ;
      RECT 92 -90.05 92.26 -71.33 ;
      RECT 91.04 -90.05 91.3 -71.33 ;
      RECT 90.08 -90.05 90.34 -71.33 ;
      RECT 89.12 -90.05 89.38 -71.33 ;
      RECT 88.16 -90.05 88.42 -71.33 ;
      RECT 87.2 -90.05 87.46 -71.33 ;
      RECT 86.24 -90.05 86.5 -71.33 ;
      RECT 85.28 -90.05 85.54 -71.33 ;
      RECT 84.32 -90.05 84.58 -71.33 ;
      RECT 83.36 -90.05 83.62 -71.33 ;
      RECT 82.4 -90.05 82.66 -71.33 ;
      RECT 81.44 -90.05 81.7 -71.33 ;
      RECT 80.48 -90.05 80.74 -71.33 ;
      RECT 79.52 -90.05 79.78 -71.33 ;
      RECT 78.56 -90.05 78.82 -71.33 ;
      RECT 77.6 -90.05 77.86 -71.33 ;
      RECT 76.64 -90.05 76.9 -71.33 ;
      RECT 75.68 -90.05 75.94 -71.33 ;
      RECT 74.72 -90.05 74.98 -71.33 ;
      RECT 73.76 -90.05 74.02 -71.33 ;
      RECT 72.8 -90.05 73.06 -71.33 ;
      RECT 71.84 -90.05 72.1 -71.33 ;
      RECT 70.88 -90.05 71.14 -71.33 ;
      RECT 69.92 -90.05 70.18 -71.33 ;
      RECT 68.96 -90.05 69.22 -71.33 ;
      RECT 68 -90.05 68.26 -71.33 ;
      RECT 67.04 -90.05 67.3 -71.33 ;
      RECT 66.08 -90.05 66.34 -71.33 ;
      RECT 60.26 -90.05 65.38 -71.33 ;
      RECT 60.26 -90.03 125.11 -71.35 ;
      RECT 48.19 -96.81 49.72 -62.77 ;
      RECT 33.57 -86.67 47.25 -70.55 ;
      RECT 48.19 -96.81 51.06 -72.04 ;
      RECT 31.6 -96.81 35.84 -72.07 ;
      RECT 29 -96.81 30.8 -70.21 ;
      RECT -0.34 -91.66 25.54 -70.12 ;
      RECT 51.86 -96.81 53.67 -70.42 ;
      RECT 31.6 -86.67 51.06 -72.96 ;
      RECT 26.08 -76.52 125.11 -73.18 ;
      RECT 47.14 -96.81 58.5 -73.18 ;
      RECT 3.72 -96.81 35.84 -73.24 ;
      RECT 47.14 -96.81 63 -78.28 ;
      RECT 46.08 -90.03 125.11 -78.28 ;
      RECT 43.63 -86.73 45.28 -69.38 ;
      RECT -0.34 -86.68 42.83 -73.24 ;
      RECT 39.09 -96.81 42.83 -66.97 ;
      RECT 43.63 -90.26 45.22 -69.38 ;
      RECT 39.09 -90.26 45.22 -87.45 ;
      RECT 3.72 -96.81 44.52 -87.46 ;
      RECT -0.34 -88.15 125.11 -87.77 ;
      RECT 45.53 -90.45 64.8 -89.19 ;
      RECT 121.76 -90.05 122.02 -71.33 ;
      RECT 120.8 -90.05 121.06 -71.33 ;
      RECT 119.84 -90.05 120.1 -71.33 ;
      RECT 118.88 -90.05 119.14 -71.33 ;
      RECT -0.34 -90.26 64.8 -89.19 ;
      RECT 64.52 -96.81 124.02 -90.77 ;
      RECT -0.34 -96.81 2.84 -48.96 ;
      RECT -0.34 -96.81 44.52 -92.54 ;
      RECT 47.14 -96.81 125.11 -92.93 ;
      RECT -0.34 -96.81 125.11 -93.09 ;
      RECT 23.72 -62.07 24.12 -61.77 ;
    LAYER M2 ;
      RECT 122.72 -92.5 122.98 -72.93 ;
      RECT 121.76 -92.5 122.02 -72.93 ;
      RECT 120.8 -92.5 121.06 -72.93 ;
      RECT 119.84 -92.5 120.1 -72.93 ;
      RECT 118.88 -92.5 119.14 -72.93 ;
      RECT 117.92 -92.5 118.18 -72.93 ;
      RECT 116.96 -92.5 117.22 -72.93 ;
      RECT 116 -92.5 116.26 -72.93 ;
      RECT 115.04 -92.5 115.3 -72.93 ;
      RECT 114.08 -92.5 114.34 -72.93 ;
      RECT 113.12 -92.5 113.38 -72.93 ;
      RECT 112.16 -92.5 112.42 -72.93 ;
      RECT 111.2 -92.5 111.46 -72.93 ;
      RECT 110.24 -92.5 110.5 -72.93 ;
      RECT 109.28 -92.5 109.54 -72.93 ;
      RECT 108.32 -92.5 108.58 -72.93 ;
      RECT 107.36 -92.5 107.62 -72.93 ;
      RECT 106.4 -92.5 106.66 -72.93 ;
      RECT 105.44 -92.5 105.7 -72.93 ;
      RECT 104.48 -92.5 104.74 -72.93 ;
      RECT 103.52 -92.5 103.78 -72.93 ;
      RECT 102.56 -92.5 102.82 -72.93 ;
      RECT 101.6 -92.5 101.86 -72.93 ;
      RECT 100.64 -96.35 100.9 -72.93 ;
      RECT 99.68 -96.35 99.94 -72.93 ;
      RECT 98.72 -96.35 98.98 -72.93 ;
      RECT 97.76 -96.35 98.02 -72.93 ;
      RECT 96.8 -96.35 97.06 -72.93 ;
      RECT 95.84 -96.35 96.1 -72.93 ;
      RECT 94.88 -96.35 95.14 -72.93 ;
      RECT 93.92 -96.35 94.18 -72.93 ;
      RECT 92.96 -96.35 93.22 -72.93 ;
      RECT 92 -96.35 92.26 -72.93 ;
      RECT 91.04 -96.35 91.3 -72.93 ;
      RECT 90.08 -96.35 90.34 -72.93 ;
      RECT 89.12 -96.35 89.38 -72.93 ;
      RECT 88.16 -96.35 88.42 -72.93 ;
      RECT 87.2 -96.35 87.46 -72.93 ;
      RECT 86.24 -92.5 86.5 -72.93 ;
      RECT 85.28 -92.5 85.54 -72.93 ;
      RECT 84.32 -92.5 84.58 -72.93 ;
      RECT 83.36 -92.5 83.62 -72.93 ;
      RECT 82.4 -92.5 82.66 -72.93 ;
      RECT 81.44 -92.5 81.7 -72.93 ;
      RECT 80.48 -92.5 80.74 -72.93 ;
      RECT 79.52 -92.5 79.78 -72.93 ;
      RECT 78.56 -92.5 78.82 -72.93 ;
      RECT 77.6 -92.5 77.86 -72.93 ;
      RECT 76.64 -92.5 76.9 -72.93 ;
      RECT 75.68 -92.5 75.94 -72.93 ;
      RECT 74.72 -92.5 74.98 -72.93 ;
      RECT 73.76 -92.5 74.02 -72.93 ;
      RECT 72.8 -92.5 73.06 -72.93 ;
      RECT 71.84 -92.5 72.1 -72.93 ;
      RECT 70.88 -92.5 71.14 -72.93 ;
      RECT 69.92 -92.5 70.18 -72.93 ;
      RECT 68.96 -92.5 69.22 -72.93 ;
      RECT 68 -92.5 68.26 -72.93 ;
      RECT 67.04 -92.5 67.3 -72.93 ;
      RECT 66.08 -92.5 66.34 -72.93 ;
      RECT 65.12 -92.5 65.38 -72.93 ;
      RECT 65.12 -92.5 122.98 -92.22 ;
      RECT 86.55 -96.35 101.55 -92.22 ;
      RECT 86.55 -69.65 101.55 -67.87 ;
      RECT 66.12 -69.65 121.98 -68.77 ;
      RECT 121.28 -88.43 121.54 -68.77 ;
      RECT 120.32 -88.43 120.58 -68.77 ;
      RECT 119.36 -88.43 119.62 -68.77 ;
      RECT 118.4 -88.43 118.66 -68.77 ;
      RECT 117.44 -88.43 117.7 -68.77 ;
      RECT 116.48 -88.43 116.74 -68.77 ;
      RECT 115.52 -88.43 115.78 -68.77 ;
      RECT 114.56 -88.43 114.82 -68.77 ;
      RECT 113.6 -88.43 113.86 -68.77 ;
      RECT 112.64 -88.43 112.9 -68.77 ;
      RECT 111.68 -88.43 111.94 -68.77 ;
      RECT 110.72 -88.43 110.98 -68.77 ;
      RECT 109.76 -88.43 110.02 -68.77 ;
      RECT 108.8 -88.43 109.06 -68.77 ;
      RECT 107.84 -88.43 108.1 -68.77 ;
      RECT 106.88 -88.43 107.14 -68.77 ;
      RECT 105.92 -88.43 106.18 -68.77 ;
      RECT 104.96 -88.43 105.22 -68.77 ;
      RECT 104 -88.43 104.26 -68.77 ;
      RECT 103.04 -88.43 103.3 -68.77 ;
      RECT 102.08 -88.43 102.34 -68.77 ;
      RECT 101.12 -88.43 101.38 -67.87 ;
      RECT 100.16 -88.43 100.42 -67.87 ;
      RECT 99.2 -88.43 99.46 -67.87 ;
      RECT 98.24 -88.43 98.5 -67.87 ;
      RECT 97.28 -88.43 97.54 -67.87 ;
      RECT 96.32 -88.43 96.58 -67.87 ;
      RECT 95.36 -88.43 95.62 -67.87 ;
      RECT 94.4 -88.43 94.66 -67.87 ;
      RECT 93.44 -88.43 93.7 -67.87 ;
      RECT 92.48 -88.43 92.74 -67.87 ;
      RECT 91.52 -88.43 91.78 -67.87 ;
      RECT 90.56 -88.43 90.82 -67.87 ;
      RECT 89.6 -88.43 89.86 -67.87 ;
      RECT 88.64 -88.43 88.9 -67.87 ;
      RECT 87.68 -88.43 87.94 -67.87 ;
      RECT 86.72 -88.43 86.98 -67.87 ;
      RECT 85.76 -88.43 86.02 -68.77 ;
      RECT 84.8 -88.43 85.06 -68.77 ;
      RECT 83.84 -88.43 84.1 -68.77 ;
      RECT 82.88 -88.43 83.14 -68.77 ;
      RECT 81.92 -88.43 82.18 -68.77 ;
      RECT 80.96 -88.43 81.22 -68.77 ;
      RECT 80 -88.43 80.26 -68.77 ;
      RECT 79.04 -88.43 79.3 -68.77 ;
      RECT 78.08 -88.43 78.34 -68.77 ;
      RECT 77.12 -88.43 77.38 -68.77 ;
      RECT 76.16 -88.43 76.42 -68.77 ;
      RECT 75.2 -88.43 75.46 -68.77 ;
      RECT 74.24 -88.43 74.5 -68.77 ;
      RECT 73.28 -88.43 73.54 -68.77 ;
      RECT 72.32 -88.43 72.58 -68.77 ;
      RECT 71.36 -88.43 71.62 -68.77 ;
      RECT 70.4 -88.43 70.66 -68.77 ;
      RECT 69.44 -88.43 69.7 -68.77 ;
      RECT 68.48 -88.43 68.74 -68.77 ;
      RECT 67.52 -88.43 67.78 -68.77 ;
      RECT 66.56 -88.43 66.82 -68.77 ;
      RECT 24.02 -66.11 84.63 -65.25 ;
      RECT 38.35 -67.25 84.63 -65.25 ;
      RECT 24.02 -67.25 34.21 -65.25 ;
      RECT 38.35 -68.33 39.11 -65.25 ;
      RECT 38.35 -68.33 49.39 -68.03 ;
      RECT 35.24 -71.56 48.18 -71.16 ;
      RECT 47.82 -94.49 48.18 -71.16 ;
      RECT 47.82 -94.49 48.22 -73.58 ;
      RECT 24.08 -61.42 24.68 -59.06 ;
      RECT 11.3 -61.17 24.68 -59.17 ;
      RECT 20.1 -63.33 22.1 -59.17 ;
      RECT 122.24 -88.43 122.5 -71.57 ;
      RECT 65.6 -88.43 65.86 -71.57 ;
    LAYER M2 SPACING 0.2 ;
      RECT -0.34 -50.64 125.11 -48.96 ;
      RECT 101.85 -68.47 125.11 -48.96 ;
      RECT 51.46 -50.65 125.11 -48.96 ;
      RECT -0.34 -51.72 48.88 -48.96 ;
      RECT 51.46 -68.47 86.25 -48.96 ;
      RECT 35.35 -67.73 48.88 -48.96 ;
      RECT -0.34 -52.24 33.75 -48.96 ;
      RECT 28.18 -53.7 33.75 -48.96 ;
      RECT 33.55 -70.86 33.75 -48.96 ;
      RECT -0.34 -53.66 26.98 -48.96 ;
      RECT 50.73 -68.47 86.25 -53.24 ;
      RECT 51.31 -68.95 51.61 -53.24 ;
      RECT 35.35 -61.75 86.25 -53.29 ;
      RECT 50.71 -96.81 50.89 -53.29 ;
      RECT 35.04 -61.75 86.25 -53.32 ;
      RECT -0.34 -53.66 34.1 -53.42 ;
      RECT 28.1 -59.46 28.18 -53.42 ;
      RECT 27.14 -58.73 28.18 -53.42 ;
      RECT -0.34 -53.69 24.82 -48.96 ;
      RECT -0.34 -54.05 23.86 -48.96 ;
      RECT 22.18 -56.1 23.86 -48.96 ;
      RECT 31.94 -54.83 34.1 -53.32 ;
      RECT 32.68 -70.73 33.75 -48.96 ;
      RECT -0.34 -58.87 20.86 -48.96 ;
      RECT 33.62 -96.81 35.83 -54.36 ;
      RECT 24.9 -54.89 28.18 -54.55 ;
      RECT 26.66 -55 28.18 -54.55 ;
      RECT 22.18 -54.89 24.14 -54.55 ;
      RECT 31.93 -54.83 86.25 -54.56 ;
      RECT 24.9 -54.83 86.25 -54.59 ;
      RECT 31.97 -59.7 86.25 -54.36 ;
      RECT 27.14 -55.19 31.23 -54.59 ;
      RECT -0.34 -57.76 23.68 -55.37 ;
      RECT -0.34 -56.1 25.78 -55.77 ;
      RECT 26.66 -57.4 28.18 -55.89 ;
      RECT 28.18 -59.7 86.25 -56.08 ;
      RECT 24.76 -56.24 25.78 -55.77 ;
      RECT 24.98 -57.4 86.25 -56.19 ;
      RECT -0.34 -57.76 23.78 -57.18 ;
      RECT 24.98 -57.51 26.26 -56.19 ;
      RECT 22.95 -58.18 24.82 -57.44 ;
      RECT 22.95 -61.43 24.68 -57.44 ;
      RECT 23.7 -63.04 24.68 -57.44 ;
      RECT 26.66 -58.73 86.25 -58.28 ;
      RECT 24.9 -58.73 86.25 -58.39 ;
      RECT 27.14 -59.46 27.88 -53.42 ;
      RECT 9.68 -63.09 21.63 -55.37 ;
      RECT -0.34 -60.17 7.08 -48.96 ;
      RECT 4.47 -60.89 7.08 -48.96 ;
      RECT 23.7 -61.54 24.82 -58.94 ;
      RECT 9.68 -61.43 24.82 -59.08 ;
      RECT 9.68 -60.86 26.98 -59.62 ;
      RECT 28.18 -67.73 31.62 -56.08 ;
      RECT -0.34 -91.68 3.71 -48.96 ;
      RECT 9.68 -60.86 31.62 -60.64 ;
      RECT 31.65 -68.65 35.83 -60.78 ;
      RECT 4.47 -96.81 7.02 -48.96 ;
      RECT -0.34 -67.81 7.02 -60.93 ;
      RECT 9.68 -63.09 22.38 -59.08 ;
      RECT 8.34 -63.09 22.38 -61.47 ;
      RECT 26.66 -62.2 49.73 -61.75 ;
      RECT 24.9 -62.09 49.73 -61.75 ;
      RECT 28.1 -67.73 49.73 -60.78 ;
      RECT 4.45 -96.81 9.42 -62.21 ;
      RECT 23.7 -63.04 24.82 -62.3 ;
      RECT 28.1 -67.73 86.25 -62.75 ;
      RECT 10.28 -63.3 23.78 -62.75 ;
      RECT 24.98 -68.65 25.78 -62.97 ;
      RECT 26.66 -67.73 86.25 -63.09 ;
      RECT 10.28 -64.95 23.68 -62.75 ;
      RECT 24.98 -67.73 86.25 -63.39 ;
      RECT 26.39 -96.81 28.03 -63.39 ;
      RECT 4.45 -69.21 10.91 -63.93 ;
      RECT 24.76 -67.73 86.25 -64.24 ;
      RECT 23.29 -96.81 25.37 -64.38 ;
      RECT 22.4 -67.73 86.25 -64.38 ;
      RECT -0.34 -67.81 19.8 -63.93 ;
      RECT 64.5 -70.47 123.6 -66.25 ;
      RECT -0.34 -67.81 30.75 -67.55 ;
      RECT 37.11 -68.33 125.11 -66.25 ;
      RECT 50.62 -70.86 50.89 -62.75 ;
      RECT 23.29 -68.65 30.75 -64.38 ;
      RECT 26.23 -69.2 28.03 -63.39 ;
      RECT 4.45 -67.97 21.57 -67.55 ;
      RECT 36.73 -68.33 125.11 -68.03 ;
      RECT 47.34 -69.13 49.78 -62.75 ;
      RECT 37.17 -68.44 46.5 -48.96 ;
      RECT 44.35 -86.69 46.5 -48.96 ;
      RECT 38.92 -86.69 43.45 -48.96 ;
      RECT 37.17 -89.84 38.02 -48.96 ;
      RECT 50.62 -68.54 63.02 -62.75 ;
      RECT 51.93 -68.74 63.02 -48.96 ;
      RECT 58.12 -76.54 63.02 -48.96 ;
      RECT 50.62 -68.74 51.01 -62.75 ;
      RECT 3.7 -96.81 9.42 -68.57 ;
      RECT 23.29 -68.65 35.84 -68.63 ;
      RECT 32.61 -69.61 38.02 -68.65 ;
      RECT 29.1 -69.29 31.75 -68.63 ;
      RECT 57 -69.48 57.26 -48.96 ;
      RECT 54.44 -69.5 56.14 -48.96 ;
      RECT 54.52 -96.81 56.14 -48.96 ;
      RECT 51.93 -96.81 53.5 -48.96 ;
      RECT 38.86 -69 43.51 -68.8 ;
      RECT 50.6 -70.86 50.89 -69.07 ;
      RECT 48.1 -70.76 50.89 -69.07 ;
      RECT 44.35 -69.77 47.34 -69.07 ;
      RECT 10.28 -96.81 10.91 -48.96 ;
      RECT 29.1 -96.81 30.75 -56.08 ;
      RECT 51.91 -96.81 53.5 -69.46 ;
      RECT 23.29 -96.81 25.49 -69.51 ;
      RECT 21.87 -96.81 25.49 -69.53 ;
      RECT 57.17 -76.54 63.02 -69.6 ;
      RECT 54.52 -96.81 56.27 -69.6 ;
      RECT 48.1 -70.76 51.01 -69.6 ;
      RECT 37.17 -86.69 46.5 -69.36 ;
      RECT 31.65 -70.73 36.27 -69.51 ;
      RECT 51.91 -96.81 53.62 -69.68 ;
      RECT 26.39 -72.46 30.75 -69.72 ;
      RECT 47.82 -96.11 49.74 -69.89 ;
      RECT 123.28 -91.87 125.11 -69.95 ;
      RECT 3.7 -96.81 10.91 -70.05 ;
      RECT 21.87 -72.46 30.75 -70.1 ;
      RECT 26.32 -96.81 28.22 -70.1 ;
      RECT 47.26 -70.76 53.62 -70.29 ;
      RECT 54.52 -70.47 125.11 -70.38 ;
      RECT 57.09 -96.81 58.52 -70.38 ;
      RECT 54.45 -96.81 56.33 -70.4 ;
      RECT 122.24 -90.05 122.5 -48.96 ;
      RECT 121.28 -90.05 121.54 -48.96 ;
      RECT 120.32 -90.05 120.58 -48.96 ;
      RECT 119.36 -90.05 119.62 -48.96 ;
      RECT 118.4 -90.05 118.66 -48.96 ;
      RECT 117.44 -90.05 117.7 -48.96 ;
      RECT 116.48 -90.05 116.74 -48.96 ;
      RECT 115.52 -90.05 115.78 -48.96 ;
      RECT 114.56 -90.05 114.82 -48.96 ;
      RECT 113.6 -90.05 113.86 -48.96 ;
      RECT 112.64 -90.05 112.9 -48.96 ;
      RECT 111.68 -90.05 111.94 -48.96 ;
      RECT 110.72 -90.05 110.98 -48.96 ;
      RECT 109.76 -90.05 110.02 -48.96 ;
      RECT 108.8 -90.05 109.06 -48.96 ;
      RECT 107.84 -90.05 108.1 -48.96 ;
      RECT 106.88 -90.05 107.14 -48.96 ;
      RECT 105.92 -90.05 106.18 -48.96 ;
      RECT 104.96 -90.05 105.22 -48.96 ;
      RECT 104 -90.05 104.26 -48.96 ;
      RECT 103.04 -90.05 103.3 -48.96 ;
      RECT 102.08 -90.05 102.34 -48.96 ;
      RECT 101.12 -90.05 101.38 -66.25 ;
      RECT 100.16 -90.05 100.42 -66.25 ;
      RECT 99.2 -90.05 99.46 -66.25 ;
      RECT 98.24 -90.05 98.5 -66.25 ;
      RECT 97.28 -90.05 97.54 -66.25 ;
      RECT 96.32 -90.05 96.58 -66.25 ;
      RECT 95.36 -90.05 95.62 -66.25 ;
      RECT 94.4 -90.05 94.66 -66.25 ;
      RECT 93.44 -90.05 93.7 -66.25 ;
      RECT 92.48 -90.05 92.74 -66.25 ;
      RECT 91.52 -90.05 91.78 -66.25 ;
      RECT 90.56 -90.05 90.82 -66.25 ;
      RECT 89.6 -90.05 89.86 -66.25 ;
      RECT 88.64 -90.05 88.9 -66.25 ;
      RECT 87.68 -90.05 87.94 -66.25 ;
      RECT 86.72 -90.05 86.98 -66.25 ;
      RECT 85.76 -90.05 86.02 -48.96 ;
      RECT 84.8 -90.05 85.06 -48.96 ;
      RECT 83.84 -90.05 84.1 -48.96 ;
      RECT 82.88 -90.05 83.14 -48.96 ;
      RECT 81.92 -90.05 82.18 -48.96 ;
      RECT 80.96 -90.05 81.22 -48.96 ;
      RECT 80 -90.05 80.26 -48.96 ;
      RECT 79.04 -90.05 79.3 -48.96 ;
      RECT 78.08 -90.05 78.34 -48.96 ;
      RECT 77.12 -90.05 77.38 -48.96 ;
      RECT 76.16 -90.05 76.42 -48.96 ;
      RECT 75.2 -90.05 75.46 -48.96 ;
      RECT 74.24 -90.05 74.5 -48.96 ;
      RECT 73.28 -90.05 73.54 -48.96 ;
      RECT 72.32 -90.05 72.58 -48.96 ;
      RECT 71.36 -90.05 71.62 -48.96 ;
      RECT 70.4 -90.05 70.66 -48.96 ;
      RECT 69.44 -90.05 69.7 -48.96 ;
      RECT 68.48 -90.05 68.74 -48.96 ;
      RECT 67.52 -90.05 67.78 -48.96 ;
      RECT 66.56 -90.05 66.82 -48.96 ;
      RECT 65.6 -90.05 65.86 -48.96 ;
      RECT 46.06 -90.47 47.27 -70.53 ;
      RECT 21.87 -70.86 32.63 -70.19 ;
      RECT 60.24 -91.43 64.82 -69.95 ;
      RECT 48.1 -71.56 49.8 -69.07 ;
      RECT 50.67 -72.55 64.82 -70.4 ;
      RECT 47.26 -71.6 49.74 -69.89 ;
      RECT 21.87 -72.46 32.62 -70.19 ;
      RECT 118.88 -90.05 125.11 -71.31 ;
      RECT 122.72 -96.81 124.04 -71.31 ;
      RECT 117.92 -96.81 118.18 -71.31 ;
      RECT 116.96 -96.81 117.22 -71.31 ;
      RECT 116 -96.81 116.26 -71.31 ;
      RECT 115.04 -96.81 115.3 -71.31 ;
      RECT 114.08 -96.81 114.34 -71.31 ;
      RECT 113.12 -96.81 113.38 -71.31 ;
      RECT 112.16 -96.81 112.42 -71.31 ;
      RECT 111.2 -96.81 111.46 -71.31 ;
      RECT 110.24 -96.81 110.5 -71.31 ;
      RECT 109.28 -96.81 109.54 -71.31 ;
      RECT 108.32 -96.81 108.58 -71.31 ;
      RECT 107.36 -96.81 107.62 -71.31 ;
      RECT 106.4 -96.81 106.66 -71.31 ;
      RECT 105.44 -96.81 105.7 -71.31 ;
      RECT 104.48 -96.81 104.74 -71.31 ;
      RECT 103.52 -96.81 103.78 -71.31 ;
      RECT 102.56 -96.81 102.82 -71.31 ;
      RECT 101.6 -96.81 101.86 -71.31 ;
      RECT 100.64 -96.81 100.9 -71.31 ;
      RECT 99.68 -96.81 99.94 -71.31 ;
      RECT 98.72 -96.81 98.98 -71.31 ;
      RECT 97.76 -96.81 98.02 -71.31 ;
      RECT 96.8 -96.81 97.06 -71.31 ;
      RECT 95.84 -96.81 96.1 -71.31 ;
      RECT 94.88 -96.81 95.14 -71.31 ;
      RECT 93.92 -96.81 94.18 -71.31 ;
      RECT 92.96 -96.81 93.22 -71.31 ;
      RECT 92 -96.81 92.26 -71.31 ;
      RECT 91.04 -96.81 91.3 -71.31 ;
      RECT 90.08 -96.81 90.34 -71.31 ;
      RECT 89.12 -96.81 89.38 -71.31 ;
      RECT 88.16 -96.81 88.42 -71.31 ;
      RECT 87.2 -96.81 87.46 -71.31 ;
      RECT 86.24 -96.81 86.5 -71.31 ;
      RECT 85.28 -96.81 85.54 -71.31 ;
      RECT 84.32 -96.81 84.58 -71.31 ;
      RECT 83.36 -96.81 83.62 -71.31 ;
      RECT 82.4 -96.81 82.66 -71.31 ;
      RECT 81.44 -96.81 81.7 -71.31 ;
      RECT 80.48 -96.81 80.74 -71.31 ;
      RECT 79.52 -96.81 79.78 -71.31 ;
      RECT 78.56 -96.81 78.82 -71.31 ;
      RECT 77.6 -96.81 77.86 -71.31 ;
      RECT 76.64 -96.81 76.9 -71.31 ;
      RECT 75.68 -96.81 75.94 -71.31 ;
      RECT 74.72 -96.81 74.98 -71.31 ;
      RECT 73.76 -96.81 74.02 -71.31 ;
      RECT 72.8 -96.81 73.06 -71.31 ;
      RECT 71.84 -96.81 72.1 -71.31 ;
      RECT 70.88 -96.81 71.14 -71.31 ;
      RECT 69.92 -96.81 70.18 -71.31 ;
      RECT 68.96 -96.81 69.22 -71.31 ;
      RECT 68 -96.81 68.26 -71.31 ;
      RECT 67.04 -96.81 67.3 -71.31 ;
      RECT 66.08 -96.81 66.34 -71.31 ;
      RECT 64.5 -96.81 65.38 -71.31 ;
      RECT 60.24 -90.05 125.11 -71.33 ;
      RECT 33.62 -86.7 42.85 -70.51 ;
      RECT 50.66 -72.55 125.11 -71.86 ;
      RECT 33.55 -86.69 47.27 -71.86 ;
      RECT 21.87 -72.46 32.63 -71.86 ;
      RECT 48.52 -96.81 51.08 -72.02 ;
      RECT 31.58 -96.81 35.86 -72.05 ;
      RECT 28.98 -96.81 30.82 -70.19 ;
      RECT 21.87 -96.81 25.56 -70.1 ;
      RECT 51.84 -96.81 53.69 -70.4 ;
      RECT 47.12 -96.11 51.08 -72.94 ;
      RECT 21.87 -96.81 35.86 -73.22 ;
      RECT 48.52 -96.81 58.52 -73.31 ;
      RECT 48.52 -96.81 63.02 -78.26 ;
      RECT -0.34 -83.03 125.11 -78.91 ;
      RECT 43.61 -86.75 45.3 -69.36 ;
      RECT 39.07 -89.84 42.85 -48.96 ;
      RECT 36.62 -89.84 38.31 -70.51 ;
      RECT 43.61 -90.28 45.24 -69.36 ;
      RECT 39.12 -96.81 44.54 -87.43 ;
      RECT 21.87 -89.84 45.24 -87.44 ;
      RECT 21.87 -88.17 125.11 -87.75 ;
      RECT 45.51 -90.47 65.38 -89.17 ;
      RECT 39.12 -90.28 65.38 -89.17 ;
      RECT 21.87 -96.81 37.92 -87.44 ;
      RECT 121.76 -96.81 122.02 -71.31 ;
      RECT 120.8 -96.81 121.06 -71.31 ;
      RECT 119.84 -96.81 120.1 -71.31 ;
      RECT 118.88 -96.81 119.14 -71.31 ;
      RECT 64.5 -96.81 124.04 -90.91 ;
      RECT 21.87 -96.81 44.54 -91.04 ;
      RECT -0.34 -96.81 2.86 -48.96 ;
      RECT -0.34 -96.81 10.91 -92.52 ;
      RECT 48.52 -96.81 125.11 -92.91 ;
      RECT 21.87 -96.11 125.11 -93.07 ;
      RECT -0.34 -96.81 47.52 -93.97 ;
    LAYER M3 ;
      RECT 36.95 -53.02 56.55 -52.02 ;
      RECT 55.55 -96.34 56.55 -52.02 ;
      RECT 55.55 -96.34 92.71 -95.34 ;
      RECT 22.94 -59.87 23.14 -51.08 ;
      RECT 22.19 -56.2 22.39 -51.08 ;
      RECT 21.42 -52.49 21.62 -51.08 ;
    LAYER M3 SPACING 0.2 ;
      RECT 23.44 -50.65 125.11 -48.96 ;
      RECT 101.85 -68.47 125.11 -48.96 ;
      RECT -0.34 -54.11 21.12 -48.96 ;
      RECT 22.89 -61.49 23.78 -49.46 ;
      RECT -0.34 -51.72 86.25 -49.46 ;
      RECT 35.35 -67.73 86.25 -48.96 ;
      RECT 36.73 -68.47 86.25 -48.96 ;
      RECT -0.34 -52.24 33.75 -49.46 ;
      RECT 35.33 -53.02 86.25 -52.02 ;
      RECT 28.18 -70.79 33.75 -48.96 ;
      RECT 33.49 -70.86 33.75 -48.96 ;
      RECT -0.34 -54.11 26.98 -49.46 ;
      RECT 35.02 -67.73 86.25 -53.32 ;
      RECT 28.18 -70.79 34.12 -53.32 ;
      RECT 24.98 -59.46 34.12 -53.42 ;
      RECT 22.12 -56.24 34.12 -53.42 ;
      RECT -0.34 -58.87 20.92 -48.96 ;
      RECT 33.62 -96.81 35.83 -54.32 ;
      RECT -0.34 -57.82 23.78 -55.31 ;
      RECT 23.64 -63.04 26.98 -57.44 ;
      RECT 9.68 -64.95 21.69 -55.31 ;
      RECT -0.34 -96.81 7.08 -48.96 ;
      RECT 9.68 -61.49 26.98 -59.02 ;
      RECT 24.98 -96.81 32.62 -60.64 ;
      RECT 8.28 -64.95 22.44 -61.47 ;
      RECT -0.34 -96.81 10.91 -62.15 ;
      RECT 22.4 -67.87 23.78 -62.69 ;
      RECT 23.23 -96.81 32.62 -64.24 ;
      RECT -0.34 -67.97 19.8 -62.15 ;
      RECT 64.5 -70.47 123.6 -66.25 ;
      RECT -0.34 -67.87 35.83 -67.55 ;
      RECT -0.34 -67.97 21.63 -67.55 ;
      RECT 36.73 -68.5 63.02 -48.96 ;
      RECT 44.29 -68.95 63.02 -48.96 ;
      RECT 51.91 -76.6 63.02 -48.96 ;
      RECT 39.28 -96.81 43.51 -48.96 ;
      RECT 36.73 -89.84 38.08 -48.96 ;
      RECT 23.23 -70.79 38.08 -68.63 ;
      RECT 44.29 -70.76 51.01 -48.96 ;
      RECT 39.12 -96.81 47.52 -69.3 ;
      RECT 21.87 -96.81 32.62 -69.47 ;
      RECT 50.67 -96.81 58.58 -69.85 ;
      RECT 123.28 -96.81 125.11 -69.95 ;
      RECT 50.6 -70.86 64.82 -69.95 ;
      RECT 60.18 -96.81 64.82 -69.95 ;
      RECT 44.29 -96.11 49.8 -48.96 ;
      RECT 21.87 -70.86 32.69 -69.47 ;
      RECT 33.62 -89.84 49.8 -69.3 ;
      RECT 122.8 -96.81 125.11 -71.31 ;
      RECT 50.6 -76.6 125.11 -71.86 ;
      RECT 33.49 -89.84 49.8 -71.86 ;
      RECT 21.87 -96.81 32.69 -71.86 ;
      RECT 48.52 -96.81 58.58 -71.96 ;
      RECT 21.87 -96.81 37.92 -71.99 ;
      RECT 60.18 -90.05 125.11 -71.31 ;
      RECT 48.52 -96.81 65.3 -78.2 ;
      RECT -0.34 -83.03 125.11 -78.91 ;
      RECT 39.12 -95.04 125.11 -90.91 ;
      RECT 95.91 -96.81 125.11 -90.91 ;
      RECT 21.87 -96.81 38.22 -91.04 ;
      RECT 21.87 -95.04 125.11 -91.1 ;
      RECT -0.34 -96.81 47.52 -93.97 ;
      RECT 48.52 -96.81 94.33 -90.91 ;
    LAYER M4 SPACING 0.2 ;
      RECT 23.44 -51.72 125.11 -48.96 ;
      RECT 95.91 -96.81 125.11 -48.96 ;
      RECT -0.34 -54.11 21.12 -48.96 ;
      RECT 22.89 -61.49 33.75 -49.46 ;
      RECT 35.33 -76.6 125.11 -48.96 ;
      RECT 60.18 -95.04 125.11 -48.96 ;
      RECT -0.34 -54.11 33.75 -49.46 ;
      RECT 22.12 -57.82 33.75 -49.46 ;
      RECT 23.64 -96.81 37.92 -53.32 ;
      RECT -0.34 -67.97 20.92 -48.96 ;
      RECT -0.34 -57.82 125.11 -55.31 ;
      RECT -0.34 -67.87 21.69 -55.31 ;
      RECT -0.34 -61.49 125.11 -59.02 ;
      RECT -0.34 -67.87 22.44 -59.02 ;
      RECT -0.34 -67.87 125.11 -62.69 ;
      RECT 23.23 -96.81 37.92 -62.69 ;
      RECT -0.34 -67.97 21.63 -55.31 ;
      RECT -0.34 -96.81 10.91 -48.96 ;
      RECT 23.21 -69.17 125.11 -68.17 ;
      RECT 21.87 -96.81 37.92 -69.47 ;
      RECT 58.88 -76.62 59.88 -48.96 ;
      RECT 21.87 -89.84 58.58 -69.47 ;
      RECT 39.12 -96.81 94.33 -78.2 ;
      RECT -0.34 -83.03 125.11 -78.91 ;
      RECT 21.87 -96.81 38.22 -91.04 ;
      RECT 21.87 -95.04 125.11 -91.1 ;
      RECT -0.34 -96.81 94.33 -93.97 ;
  END
END LDO_Top_int

END LIBRARY
