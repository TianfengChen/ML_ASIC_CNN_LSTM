

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO writeback_controller 
  PIN clk 
    ANTENNAPARTIALMETALAREA 12.02 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1206 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2096 LAYER M4 ; 
    ANTENNAMAXAREACAR 92.9835 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.93879 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.38095 LAYER V4 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 3.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0336 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M4 ; 
    ANTENNAMAXAREACAR 122.578 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.23081 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.93633 LAYER V4 ;
  END reset
  PIN DRAM_in3_WEN 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 14.46 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1446 LAYER M4 ;
  END DRAM_in3_WEN
  PIN DRAM_in3_Data[7] 
    ANTENNADIFFAREA 3.348 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1526 LAYER M4 ;
  END DRAM_in3_Data[7]
  PIN DRAM_in3_Data[6] 
    ANTENNADIFFAREA 3.348 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 14.94 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1494 LAYER M4 ;
  END DRAM_in3_Data[6]
  PIN DRAM_in3_Data[5] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1126 LAYER M4 ;
  END DRAM_in3_Data[5]
  PIN DRAM_in3_Data[4] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M4 ;
  END DRAM_in3_Data[4]
  PIN DRAM_in3_Data[3] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0646 LAYER M4 ;
  END DRAM_in3_Data[3]
  PIN DRAM_in3_Data[2] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1112 LAYER M4 ;
  END DRAM_in3_Data[2]
  PIN DRAM_in3_Data[1] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 14.54 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1454 LAYER M4 ;
  END DRAM_in3_Data[1]
  PIN DRAM_in3_Data[0] 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 14.94 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1494 LAYER M4 ;
  END DRAM_in3_Data[0]
  PIN pk_out_3__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 91.4599 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.930128 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pk_out_3__PE_state__2_
  PIN pk_out_3__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.9412 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.225613 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_3__PE_state__1_
  PIN pk_out_3__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 26.7126 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.272794 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_3__PE_state__0_
  PIN pk_out_3__data__7_ 
  END pk_out_3__data__7_
  PIN pk_out_3__data__6_ 
  END pk_out_3__data__6_
  PIN pk_out_3__data__5_ 
  END pk_out_3__data__5_
  PIN pk_out_3__data__4_ 
  END pk_out_3__data__4_
  PIN pk_out_3__data__3_ 
  END pk_out_3__data__3_
  PIN pk_out_3__data__2_ 
  END pk_out_3__data__2_
  PIN pk_out_3__data__1_ 
  END pk_out_3__data__1_
  PIN pk_out_3__data__0_ 
  END pk_out_3__data__0_
  PIN pk_out_2__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 105.562 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.07115 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pk_out_2__PE_state__2_
  PIN pk_out_2__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 24.3922 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.250123 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_2__PE_state__1_
  PIN pk_out_2__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.2028 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.277696 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_2__PE_state__0_
  PIN pk_out_2__data__7_ 
  END pk_out_2__data__7_
  PIN pk_out_2__data__6_ 
  END pk_out_2__data__6_
  PIN pk_out_2__data__5_ 
  END pk_out_2__data__5_
  PIN pk_out_2__data__4_ 
  END pk_out_2__data__4_
  PIN pk_out_2__data__3_ 
  END pk_out_2__data__3_
  PIN pk_out_2__data__2_ 
  END pk_out_2__data__2_
  PIN pk_out_2__data__1_ 
  END pk_out_2__data__1_
  PIN pk_out_2__data__0_ 
  END pk_out_2__data__0_
  PIN pk_out_1__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 69.6651 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.712179 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pk_out_1__PE_state__2_
  PIN pk_out_1__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.451 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.220711 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_1__PE_state__1_
  PIN pk_out_1__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 LAYER M4 ; 
    ANTENNAMAXAREACAR 34.5558 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.351225 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22549 LAYER V4 ;
  END pk_out_1__PE_state__0_
  PIN pk_out_1__data__7_ 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.7072 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.403829 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__7_
  PIN pk_out_1__data__6_ 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.2117 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.448874 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__6_
  PIN pk_out_1__data__5_ 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.4099 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.430856 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__5_
  PIN pk_out_1__data__4_ 
    ANTENNAPARTIALMETALAREA 2.26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.4099 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.430856 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__4_
  PIN pk_out_1__data__3_ 
    ANTENNAPARTIALMETALAREA 2.42 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 42.3108 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.439865 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__3_
  PIN pk_out_1__data__2_ 
    ANTENNAPARTIALMETALAREA 1.62 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.5 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.331757 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__2_
  PIN pk_out_1__data__1_ 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 67.536 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.692117 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__1_
  PIN pk_out_1__data__0_ 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.5 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.331757 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pk_out_1__data__0_
  PIN pk_out_0__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6168 LAYER M4 ; 
    ANTENNAMAXAREACAR 6.89559 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.070655 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.259403 LAYER V4 ;
  END pk_out_0__PE_state__2_
  PIN pk_out_0__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 23.369 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.238038 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V4 ;
  END pk_out_0__PE_state__1_
  PIN pk_out_0__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.5316 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.321237 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V4 ;
  END pk_out_0__PE_state__0_
  PIN pk_out_0__data__7_ 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.047 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 91.4722 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.920718 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__7_
  PIN pk_out_0__data__6_ 
    ANTENNAPARTIALMETALAREA 1.7 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 15.7778 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.166088 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__6_
  PIN pk_out_0__data__5_ 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 97.0278 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.976273 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__5_
  PIN pk_out_0__data__4_ 
    ANTENNAPARTIALMETALAREA 4.3 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.043 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 132.676 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.33275 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__4_
  PIN pk_out_0__data__3_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 120.639 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.21238 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__3_
  PIN pk_out_0__data__2_ 
    ANTENNAPARTIALMETALAREA 3.82 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0382 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 141.935 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.42535 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__2_
  PIN pk_out_0__data__1_ 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 136.843 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.37442 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__1_
  PIN pk_out_0__data__0_ 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0318 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 142.861 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.43461 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END pk_out_0__data__0_
END writeback_controller

END LIBRARY
