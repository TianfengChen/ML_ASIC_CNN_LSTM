#Confidential Information of Artisan Components, Inc.
#Use subject to Artisan Components license.
#Copyright(c) 2003 Artisan Components, Inc.

#RDB genLef Version 2003Q1

NAMESCASESENSITIVE	ON ;

SITE	iosite
	SYMMETRY Y ;
	CLASS PAD ;
	SIZE 1.000 BY 247.000 ;
END	iosite

SITE	iocornersite
	SYMMETRY Y ;
	CLASS PAD ;
	SIZE 247.000 BY 247.000 ;
END	iocornersite

MACRO POSC4
	CLASS PAD INOUT ;
	FOREIGN POSC4 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN E0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER MQ ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M6 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M5 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M4 ;
			RECT 49.870 245.620 52.540 247.000 ;
		END
	END E0
	PIN E1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER MQ ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M6 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M5 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M4 ;
			RECT 53.140 245.620 55.810 247.000 ;
		END
	END E1
	PIN CK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER M5 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER LM ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER MQ ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M6 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M4 ;
			RECT 56.410 245.620 59.080 247.000 ;
		END
	END CK
	PIN PO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER MQ ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER M6 ;
			RECT 76.000 104.500 134.000 114.000 ;
		END
	END PO
	PIN PI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END PI
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POSC4

MACRO POSC3
	CLASS PAD INOUT ;
	FOREIGN POSC3 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN E0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER MQ ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M6 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M5 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M4 ;
			RECT 49.870 245.620 52.540 247.000 ;
		END
	END E0
	PIN E1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER MQ ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M6 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M5 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M4 ;
			RECT 53.140 245.620 55.810 247.000 ;
		END
	END E1
	PIN CK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER M5 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER LM ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER MQ ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M6 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M4 ;
			RECT 56.410 245.620 59.080 247.000 ;
		END
	END CK
	PIN PO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER MQ ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER M6 ;
			RECT 76.000 104.500 134.000 114.000 ;
		END
	END PO
	PIN PI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END PI
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POSC3

MACRO POSC2
	CLASS PAD INOUT ;
	FOREIGN POSC2 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN E0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER MQ ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M6 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M5 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M4 ;
			RECT 49.870 245.620 52.540 247.000 ;
		END
	END E0
	PIN E1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER MQ ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M6 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M5 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M4 ;
			RECT 53.140 245.620 55.810 247.000 ;
		END
	END E1
	PIN CK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER M5 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER LM ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER MQ ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M6 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M4 ;
			RECT 56.410 245.620 59.080 247.000 ;
		END
	END CK
	PIN PO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER MQ ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER M6 ;
			RECT 76.000 104.500 134.000 114.000 ;
		END
	END PO
	PIN PI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END PI
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POSC2

MACRO POSC1
	CLASS PAD INOUT ;
	FOREIGN POSC1 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN E0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER MQ ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M6 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M5 ;
			RECT 49.870 245.620 52.540 247.000 ;
			LAYER M4 ;
			RECT 49.870 245.620 52.540 247.000 ;
		END
	END E0
	PIN E1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER MQ ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M6 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M5 ;
			RECT 53.140 245.620 55.810 247.000 ;
			LAYER M4 ;
			RECT 53.140 245.620 55.810 247.000 ;
		END
	END E1
	PIN CK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER M5 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER LM ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER MQ ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M6 ;
			RECT 56.410 245.620 59.080 247.000 ;
			LAYER M4 ;
			RECT 56.410 245.620 59.080 247.000 ;
		END
	END CK
	PIN PO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER MQ ;
			RECT 76.000 104.500 134.000 114.000 ;
			LAYER M6 ;
			RECT 76.000 104.500 134.000 114.000 ;
		END
	END PO
	PIN PI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END PI
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			59.280 247.000
			59.280 245.420
			49.670 245.420 49.670 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			59.480 247.000
			59.480 245.220
			49.470 245.220 49.470 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POSC1

MACRO PBAREWIRE
	CLASS PAD INOUT ;
	FOREIGN PBAREWIRE 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER MQ ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M6 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M5 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M4 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M3 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M2 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M1 ;
			RECT 29.590 246.500 52.460 247.000 ;
		END
		PORT
			LAYER LM ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER MQ ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M6 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M5 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M4 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M3 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M2 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M1 ;
			RECT 4.720 246.500 27.590 247.000 ;
		END
	END P
	PIN PADR1
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER MQ ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M6 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M5 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M4 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M3 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M2 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M1 ;
			RECT 59.850 246.500 65.450 247.000 ;
		END
	END PADR1
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			65.610 247.000
			65.610 246.340
			59.690 246.340 59.690 247.000
			52.620 247.000 52.620 246.340
			29.430 246.340 29.430 247.000
			27.750 247.000 27.750 246.340
			4.560 246.340 4.560 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.850 247.000
			65.850 246.100
			59.450 246.100 59.450 247.000
			52.860 247.000 52.860 246.100
			29.190 246.100 29.190 247.000
			27.990 247.000 27.990 246.100
			4.320 246.100 4.320 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.850 247.000
			65.850 246.100
			59.450 246.100 59.450 247.000
			52.860 247.000 52.860 246.100
			29.190 246.100 29.190 247.000
			27.990 247.000 27.990 246.100
			4.320 246.100 4.320 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBAREWIRE

MACRO PANALOG
	CLASS PAD INOUT ;
	FOREIGN PANALOG 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER MQ ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M6 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M5 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M4 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M3 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M2 ;
			RECT 29.590 246.500 52.460 247.000 ;
			LAYER M1 ;
			RECT 29.590 246.500 52.460 247.000 ;
		END
		PORT
			LAYER LM ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER MQ ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M6 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M5 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M4 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M3 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M2 ;
			RECT 4.720 246.500 27.590 247.000 ;
			LAYER M1 ;
			RECT 4.720 246.500 27.590 247.000 ;
		END
	END P
	PIN PADR1
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER MQ ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M6 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M5 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M4 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M3 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M2 ;
			RECT 59.850 246.500 65.450 247.000 ;
			LAYER M1 ;
			RECT 59.850 246.500 65.450 247.000 ;
		END
	END PADR1
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			65.610 247.000
			65.610 246.340
			59.690 246.340 59.690 247.000
			52.620 247.000 52.620 246.340
			29.430 246.340 29.430 247.000
			27.750 247.000 27.750 246.340
			4.560 246.340 4.560 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.650 247.000
			65.650 246.300
			59.650 246.300 59.650 247.000
			52.660 247.000 52.660 246.300
			29.390 246.300 29.390 247.000
			27.790 247.000 27.790 246.300
			4.520 246.300 4.520 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.850 247.000
			65.850 246.100
			59.450 246.100 59.450 247.000
			52.860 247.000 52.860 246.100
			29.190 246.100 29.190 247.000
			27.990 247.000 27.990 246.100
			4.320 246.100 4.320 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.850 247.000
			65.850 246.100
			59.450 246.100 59.450 247.000
			52.860 247.000 52.860 246.100
			29.190 246.100 29.190 247.000
			27.990 247.000 27.990 246.100
			4.320 246.100 4.320 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PANALOG

MACRO PAVSS
	CLASS PAD POWER ;
	FOREIGN PAVSS 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN AVSS
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER MQ ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M6 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M5 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M4 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M3 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M2 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M1 ;
			RECT 35.990 246.500 65.170 247.000 ;
		END
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER MQ ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M6 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M5 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M4 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M3 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M2 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M1 ;
			RECT 4.830 246.500 34.070 247.000 ;
		END
	END AVSS
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			65.330 247.000
			65.330 246.340
			35.830 246.340 35.830 247.000
			34.230 247.000 34.230 246.340
			4.670 246.340 4.670 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.570 247.000
			65.570 246.100
			35.590 246.100 35.590 247.000
			34.470 247.000 34.470 246.100
			4.430 246.100 4.430 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.570 247.000
			65.570 246.100
			35.590 246.100 35.590 247.000
			34.470 247.000 34.470 246.100
			4.430 246.100 4.430 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PAVSS

MACRO PAVDD
	CLASS PAD POWER ;
	FOREIGN PAVDD 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN AVDD
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER MQ ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M6 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M5 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M5 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M4 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M3 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M2 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M1 ;
			RECT 35.960 246.500 63.100 247.000 ;
		END
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER MQ ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M6 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M5 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M5 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M4 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M3 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M2 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M1 ;
			RECT 6.900 246.500 34.040 247.000 ;
		END
	END AVDD
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			63.260 247.000
			63.260 246.340
			35.800 246.340 35.800 247.000
			34.200 247.000 34.200 246.340
			6.740 246.340 6.740 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			63.500 247.000
			63.500 246.100
			35.560 246.100 35.560 247.000
			34.440 247.000 34.440 246.100
			6.500 246.100 6.500 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			63.500 247.000
			63.500 246.100
			35.560 246.100 35.560 247.000
			34.440 247.000 34.440 246.100
			6.500 246.100 6.500 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PAVDD

MACRO PVDD
	CLASS PAD POWER ;
	FOREIGN PVDD 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER MQ ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M6 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M5 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M5 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M4 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M3 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M2 ;
			RECT 35.960 246.500 63.100 247.000 ;
			LAYER M1 ;
			RECT 35.960 246.500 63.100 247.000 ;
		END
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER MQ ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M6 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M5 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M5 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M4 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M3 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M2 ;
			RECT 6.900 246.500 34.040 247.000 ;
			LAYER M1 ;
			RECT 6.900 246.500 34.040 247.000 ;
		END
	END VDD
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			63.260 247.000
			63.260 246.340
			35.800 246.340 35.800 247.000
			34.200 247.000 34.200 246.340
			6.740 246.340 6.740 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			63.300 247.000
			63.300 246.300
			35.760 246.300 35.760 247.000
			34.240 247.000 34.240 246.300
			6.700 246.300 6.700 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			63.500 247.000
			63.500 246.100
			35.560 246.100 35.560 247.000
			34.440 247.000 34.440 246.100
			6.500 246.100 6.500 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			63.500 247.000
			63.500 246.100
			35.560 246.100 35.560 247.000
			34.440 247.000 34.440 246.100
			6.500 246.100 6.500 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PVDD

MACRO PVSS
	CLASS PAD POWER ;
	FOREIGN PVSS 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER MQ ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M6 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M5 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M4 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M2 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M1 ;
			RECT 35.990 246.500 65.170 247.000 ;
			LAYER M3 ;
			RECT 35.990 246.500 65.170 247.000 ;
		END
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER MQ ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M6 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M5 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M4 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M2 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M1 ;
			RECT 4.830 246.500 34.070 247.000 ;
			LAYER M3 ;
			RECT 4.830 246.500 34.070 247.000 ;
		END
	END VSS
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			65.330 247.000
			65.330 246.340
			35.830 246.340 35.830 247.000
			34.230 247.000 34.230 246.340
			4.670 246.340 4.670 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			65.370 247.000
			65.370 246.300
			35.790 246.300 35.790 247.000
			34.270 247.000 34.270 246.300
			4.630 246.300 4.630 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.570 247.000
			65.570 246.100
			35.590 246.100 35.590 247.000
			34.470 247.000 34.470 246.100
			4.430 246.100 4.430 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			65.570 247.000
			65.570 246.100
			35.590 246.100 35.590 247.000
			34.470 247.000 34.470 246.100
			4.430 246.100 4.430 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PVSS

MACRO PDVDD
	CLASS PAD POWER ;
	FOREIGN PDVDD 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN DVDD
		DIRECTION INOUT ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END DVDD
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PDVDD

MACRO PDVSS
	CLASS PAD POWER ;
	FOREIGN PDVSS 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN DVSS
		DIRECTION INOUT ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END DVSS
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PDVSS

MACRO PFILLQ
	CLASS PAD SPACER ;
	FOREIGN PFILLQ 0 0 ;
	ORIGIN 0 0 ;
	SIZE 17.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 16.920 0.000 16.920 246.840
			16.840 246.840 
			16.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 
			16.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 16.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 
			16.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 16.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 
			16.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 16.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 
			16.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 16.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 
			16.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 16.900 0.000 16.900 246.800
			16.800 246.800 16.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 16.800 0.000 16.800 246.600
			16.600 246.600 
			16.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 16.800 0.000 16.800 246.600
			16.600 246.600 16.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 16.800 0.000 16.800 246.600
			16.600 246.600 
			16.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 16.800 0.000 16.800 246.600
			16.600 246.600 16.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PFILLQ

MACRO PFILLH
	CLASS PAD SPACER ;
	FOREIGN PFILLH 0 0 ;
	ORIGIN 0 0 ;
	SIZE 34.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 33.920 0.000 33.920 246.840
			33.840 246.840 
			33.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 
			33.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 33.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 
			33.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 33.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 
			33.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 33.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 
			33.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 33.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 
			33.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 33.900 0.000 33.900 246.800
			33.800 246.800 33.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 33.800 0.000 33.800 246.600
			33.600 246.600 
			33.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 33.800 0.000 33.800 246.600
			33.600 246.600 33.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 33.800 0.000 33.800 246.600
			33.600 246.600 
			33.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 33.800 0.000 33.800 246.600
			33.600 246.600 33.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PFILLH

MACRO PFILL1
	CLASS PAD SPACER ;
	FOREIGN PFILL1 0 0 ;
	ORIGIN 0 0 ;
	SIZE 1.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
                LAYER M1 ;
                POLYGON 0.080 0.000 0.920 0.000 0.920 246.840
                        0.840 246.840
                        0.840 247.000
                        0.160 247.000 0.160 246.840 0.080 246.840
                        0.080 0.000 ;
                LAYER M2 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800
                        0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER V1 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800 0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER M3 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800
                        0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER V2 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800 0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER M4 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800
                        0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER V3 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800 0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER M5 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800
                        0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER V4 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800 0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER M6 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800
                        0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER V5 ;
                POLYGON 0.100 0.000 0.900 0.000 0.900 246.800
                        0.800 246.800 0.800 247.000
                        0.200 247.000 0.200 246.800 0.100 246.800
                        0.100 0.000 ;
                LAYER MQ ;
                POLYGON 0.200 0.000 0.800 0.000 0.800 246.600
                        0.200 246.600
                        0.200 0.000 ;
                LAYER VL ;
                POLYGON 0.200 0.000 0.800 0.000 0.800 246.600
                        0.200 246.600
                        0.200 0.000 ;
                LAYER LM ;
                POLYGON 0.200 0.000 0.800 0.000 0.800 246.600
                        0.200 246.600
                        0.200 0.000 ;
                LAYER VQ ;
                POLYGON 0.200 0.000 0.800 0.000 0.800 246.600
                        0.200 246.600
                        0.200 0.000 ;
END
END PFILL1

MACRO PCORNER
	CLASS ENDCAP BOTTOMLEFT ;
	FOREIGN PCORNER 0 0 ;
	ORIGIN 0 0 ;
	SIZE 247.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iocornersite ;
	OBS
		LAYER M1 ;
		POLYGON 0.000 0.000 246.920 0.000 246.920 246.840
			246.840 246.840 
			246.840 246.920 
			0.000 246.920
			0.000 0.000 ;
		LAYER M2 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 
			246.800 246.900 
			0.000 246.900
			0.000 0.000 ;
		LAYER V1 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 246.800 246.900
			0.000 246.900
			0.000 0.000 ;
		LAYER M3 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 
			246.800 246.900 
			0.000 246.900
			0.000 0.000 ;
		LAYER V2 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 246.800 246.900
			0.000 246.900
			0.000 0.000 ;
		LAYER M4 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 
			246.800 246.900 
			0.000 246.900
			0.000 0.000 ;
		LAYER V3 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 246.800 246.900
			0.000 246.900
			0.000 0.000 ;
		LAYER M5 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 
			246.800 246.900 
			0.000 246.900
			0.000 0.000 ;
		LAYER V4 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 246.800 246.900
			0.000 246.900
			0.000 0.000 ;
		LAYER M6 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 
			246.800 246.900 
			0.000 246.900
			0.000 0.000 ;
		LAYER V5 ;
		POLYGON 0.000 0.000 246.900 0.000 246.900 246.800
			246.800 246.800 246.800 246.900
			0.000 246.900
			0.000 0.000 ;
		LAYER MQ ;
		POLYGON 0.000 0.000 246.800 0.000 246.800 246.600
			246.600 246.600 
			246.600 246.800 
			0.000 246.800
			0.000 0.000 ;
		LAYER VL ;
		POLYGON 0.000 0.000 246.800 0.000 246.800 246.600
			246.600 246.600 246.600 246.800
			0.000 246.800
			0.000 0.000 ;
		LAYER LM ;
		POLYGON 0.000 0.000 246.800 0.000 246.800 246.600
			246.600 246.600 
			246.600 246.800 
			0.000 246.800
			0.000 0.000 ;
		LAYER VQ ;
		POLYGON 0.000 0.000 246.800 0.000 246.800 246.600
			246.600 246.600 246.600 246.800
			0.000 246.800
			0.000 0.000 ;
END
END PCORNER

MACRO PBREAKBFDVDDR
	CLASS PAD SPACER ;
	FOREIGN PBREAKBFDVDDR 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBREAKBFDVDDR

MACRO PBREAKDVDDR
	CLASS PAD SPACER ;
	FOREIGN PBREAKDVDDR 0 0 ;
	ORIGIN 0 0 ;
	SIZE 140.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 139.920 0.000 139.920 246.840
			139.840 246.840 
			139.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 
			139.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 139.900 0.000 139.900 246.800
			139.800 246.800 139.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 
			139.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 139.800 0.000 139.800 246.600
			139.600 246.600 139.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBREAKDVDDR

MACRO PBREAKBF
	CLASS PAD SPACER ;
	FOREIGN PBREAKBF 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBREAKBF

MACRO PBREAK
	CLASS PAD SPACER ;
	FOREIGN PBREAK 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBREAK

MACRO POCT8C
	CLASS PAD OUTPUT ;
	FOREIGN POCT8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT8C

MACRO POCT8B
	CLASS PAD OUTPUT ;
	FOREIGN POCT8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT8B

MACRO POCT8A
	CLASS PAD OUTPUT ;
	FOREIGN POCT8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT8A

MACRO POCT4C
	CLASS PAD OUTPUT ;
	FOREIGN POCT4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT4C

MACRO POCT4A
	CLASS PAD OUTPUT ;
	FOREIGN POCT4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT4A

MACRO POCT2C
	CLASS PAD OUTPUT ;
	FOREIGN POCT2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT2C

MACRO POCT2A
	CLASS PAD OUTPUT ;
	FOREIGN POCT2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT2A

MACRO POCT24C
	CLASS PAD OUTPUT ;
	FOREIGN POCT24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT24C

MACRO POCT24B
	CLASS PAD OUTPUT ;
	FOREIGN POCT24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT24B

MACRO POCT24A
	CLASS PAD OUTPUT ;
	FOREIGN POCT24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT24A

MACRO POCT16C
	CLASS PAD OUTPUT ;
	FOREIGN POCT16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT16C

MACRO POCT16B
	CLASS PAD OUTPUT ;
	FOREIGN POCT16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT16B

MACRO POCT16A
	CLASS PAD OUTPUT ;
	FOREIGN POCT16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT16A

MACRO POCT12C
	CLASS PAD OUTPUT ;
	FOREIGN POCT12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT12C

MACRO POCT12B
	CLASS PAD OUTPUT ;
	FOREIGN POCT12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT12B

MACRO POCT12A
	CLASS PAD OUTPUT ;
	FOREIGN POCT12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POCT12A

MACRO POOD8C
	CLASS PAD OUTPUT ;
	FOREIGN POOD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD8C

MACRO POOD8B
	CLASS PAD OUTPUT ;
	FOREIGN POOD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD8B

MACRO POOD8A
	CLASS PAD OUTPUT ;
	FOREIGN POOD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD8A

MACRO POOD4C
	CLASS PAD OUTPUT ;
	FOREIGN POOD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD4C

MACRO POOD4A
	CLASS PAD OUTPUT ;
	FOREIGN POOD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD4A

MACRO POOD2C
	CLASS PAD OUTPUT ;
	FOREIGN POOD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD2C

MACRO POOD2A
	CLASS PAD OUTPUT ;
	FOREIGN POOD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD2A

MACRO POOD24C
	CLASS PAD OUTPUT ;
	FOREIGN POOD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD24C

MACRO POOD24B
	CLASS PAD OUTPUT ;
	FOREIGN POOD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD24B

MACRO POOD24A
	CLASS PAD OUTPUT ;
	FOREIGN POOD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD24A

MACRO POOD16C
	CLASS PAD OUTPUT ;
	FOREIGN POOD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD16C

MACRO POOD16B
	CLASS PAD OUTPUT ;
	FOREIGN POOD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD16B

MACRO POOD16A
	CLASS PAD OUTPUT ;
	FOREIGN POOD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD16A

MACRO POOD12C
	CLASS PAD OUTPUT ;
	FOREIGN POOD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD12C

MACRO POOD12B
	CLASS PAD OUTPUT ;
	FOREIGN POOD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD12B

MACRO POOD12A
	CLASS PAD OUTPUT ;
	FOREIGN POOD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOD12A

MACRO POOC8C
	CLASS PAD OUTPUT ;
	FOREIGN POOC8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC8C

MACRO POOC8B
	CLASS PAD OUTPUT ;
	FOREIGN POOC8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC8B

MACRO POOC8A
	CLASS PAD OUTPUT ;
	FOREIGN POOC8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC8A

MACRO POOC4C
	CLASS PAD OUTPUT ;
	FOREIGN POOC4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC4C

MACRO POOC4A
	CLASS PAD OUTPUT ;
	FOREIGN POOC4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC4A

MACRO POOC2C
	CLASS PAD OUTPUT ;
	FOREIGN POOC2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC2C

MACRO POOC2A
	CLASS PAD OUTPUT ;
	FOREIGN POOC2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC2A

MACRO POOC24C
	CLASS PAD OUTPUT ;
	FOREIGN POOC24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC24C

MACRO POOC24B
	CLASS PAD OUTPUT ;
	FOREIGN POOC24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC24B

MACRO POOC24A
	CLASS PAD OUTPUT ;
	FOREIGN POOC24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC24A

MACRO POOC16C
	CLASS PAD OUTPUT ;
	FOREIGN POOC16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC16C

MACRO POOC16B
	CLASS PAD OUTPUT ;
	FOREIGN POOC16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC16B

MACRO POOC16A
	CLASS PAD OUTPUT ;
	FOREIGN POOC16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC16A

MACRO POOC12C
	CLASS PAD OUTPUT ;
	FOREIGN POOC12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC12C

MACRO POOC12B
	CLASS PAD OUTPUT ;
	FOREIGN POOC12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC12B

MACRO POOC12A
	CLASS PAD OUTPUT ;
	FOREIGN POOC12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			54.650 245.420 54.650 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			54.450 245.220 54.450 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POOC12A

MACRO POC8C
	CLASS PAD OUTPUT ;
	FOREIGN POC8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC8C

MACRO POC8B
	CLASS PAD OUTPUT ;
	FOREIGN POC8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC8B

MACRO POC8A
	CLASS PAD OUTPUT ;
	FOREIGN POC8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC8A

MACRO POC4C
	CLASS PAD OUTPUT ;
	FOREIGN POC4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC4C

MACRO POC4A
	CLASS PAD OUTPUT ;
	FOREIGN POC4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC4A

MACRO POC2C
	CLASS PAD OUTPUT ;
	FOREIGN POC2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC2C

MACRO POC2A
	CLASS PAD OUTPUT ;
	FOREIGN POC2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC2A

MACRO POC24C
	CLASS PAD OUTPUT ;
	FOREIGN POC24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC24C

MACRO POC24B
	CLASS PAD OUTPUT ;
	FOREIGN POC24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC24B

MACRO POC24A
	CLASS PAD OUTPUT ;
	FOREIGN POC24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC24A

MACRO POC16C
	CLASS PAD OUTPUT ;
	FOREIGN POC16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC16C

MACRO POC16B
	CLASS PAD OUTPUT ;
	FOREIGN POC16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC16B

MACRO POC16A
	CLASS PAD OUTPUT ;
	FOREIGN POC16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC16A

MACRO POC12C
	CLASS PAD OUTPUT ;
	FOREIGN POC12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC12C

MACRO POC12B
	CLASS PAD OUTPUT ;
	FOREIGN POC12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC12B

MACRO POC12A
	CLASS PAD OUTPUT ;
	FOREIGN POC12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			60.950 247.000
			60.950 245.460
			57.960 245.460 57.960 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			60.990 247.000
			60.990 245.420
			57.920 245.420 57.920 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			61.190 247.000
			61.190 245.220
			57.720 245.220 57.720 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END POC12A

MACRO PICU
	CLASS PAD INPUT ;
	FOREIGN PICU 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PICU

MACRO PICSU
	CLASS PAD INPUT ;
	FOREIGN PICSU 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PICSU

MACRO PICSD
	CLASS PAD INPUT ;
	FOREIGN PICSD 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PICSD

MACRO PICD
	CLASS PAD INPUT ;
	FOREIGN PICD 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PICD

MACRO PICS
	CLASS PAD INPUT ;
	FOREIGN PICS 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PICS

MACRO PIC
	CLASS PAD INPUT ;
	FOREIGN PIC 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN P
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			61.190 245.420 61.190 247.000
			54.450 247.000 54.450 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			60.990 245.220 60.990 247.000
			54.650 247.000 54.650 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PIC

MACRO PBCSCTU8C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU8C

MACRO PBCSCTU8B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU8B

MACRO PBCSCTU8A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU8A

MACRO PBCSCTU4C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU4C

MACRO PBCSCTU4A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU4A

MACRO PBCSCTU2C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU2C

MACRO PBCSCTU2A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU2A

MACRO PBCSCTU24C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU24C

MACRO PBCSCTU24B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU24B

MACRO PBCSCTU24A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU24A

MACRO PBCSCTU16C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU16C

MACRO PBCSCTU16B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU16B

MACRO PBCSCTU16A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU16A

MACRO PBCSCTU12C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU12C

MACRO PBCSCTU12B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU12B

MACRO PBCSCTU12A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTU12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTU12A

MACRO PBCCTU8C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU8C

MACRO PBCCTU8B
	CLASS PAD INOUT ;
	FOREIGN PBCCTU8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU8B

MACRO PBCCTU8A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU8A

MACRO PBCCTU4C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU4C

MACRO PBCCTU4A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU4A

MACRO PBCCTU2C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU2C

MACRO PBCCTU2A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU2A

MACRO PBCCTU24C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU24C

MACRO PBCCTU24B
	CLASS PAD INOUT ;
	FOREIGN PBCCTU24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU24B

MACRO PBCCTU24A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU24A

MACRO PBCCTU16C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU16C

MACRO PBCCTU16B
	CLASS PAD INOUT ;
	FOREIGN PBCCTU16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU16B

MACRO PBCCTU16A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU16A

MACRO PBCCTU12C
	CLASS PAD INOUT ;
	FOREIGN PBCCTU12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU12C

MACRO PBCCTU12B
	CLASS PAD INOUT ;
	FOREIGN PBCCTU12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU12B

MACRO PBCCTU12A
	CLASS PAD INOUT ;
	FOREIGN PBCCTU12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTU12A

MACRO PBCSOCU8C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU8C

MACRO PBCSOCU8B
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU8B

MACRO PBCSOCU8A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU8A

MACRO PBCSOCU4C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU4C

MACRO PBCSOCU4A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU4A

MACRO PBCSOCU2C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU2C

MACRO PBCSOCU2A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU2A

MACRO PBCSOCU24C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU24C

MACRO PBCSOCU24B
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU24B

MACRO PBCSOCU24A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU24A

MACRO PBCSOCU16C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU16C

MACRO PBCSOCU16B
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU16B

MACRO PBCSOCU16A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU16A

MACRO PBCSOCU12C
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU12C

MACRO PBCSOCU12B
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU12B

MACRO PBCSOCU12A
	CLASS PAD INOUT ;
	FOREIGN PBCSOCU12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOCU12A

MACRO PBCOCU8C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU8C

MACRO PBCOCU8B
	CLASS PAD INOUT ;
	FOREIGN PBCOCU8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU8B

MACRO PBCOCU8A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU8A

MACRO PBCOCU4C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU4C

MACRO PBCOCU4A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU4A

MACRO PBCOCU2C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU2C

MACRO PBCOCU2A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU2A

MACRO PBCOCU24C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU24C

MACRO PBCOCU24B
	CLASS PAD INOUT ;
	FOREIGN PBCOCU24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU24B

MACRO PBCOCU24A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU24A

MACRO PBCOCU16C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU16C

MACRO PBCOCU16B
	CLASS PAD INOUT ;
	FOREIGN PBCOCU16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU16B

MACRO PBCOCU16A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU16A

MACRO PBCOCU12C
	CLASS PAD INOUT ;
	FOREIGN PBCOCU12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU12C

MACRO PBCOCU12B
	CLASS PAD INOUT ;
	FOREIGN PBCOCU12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU12B

MACRO PBCOCU12A
	CLASS PAD INOUT ;
	FOREIGN PBCOCU12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN PU
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER MQ ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M6 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M5 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M4 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M3 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M2 ;
			RECT 45.040 245.620 47.710 247.000 ;
			LAYER M1 ;
			RECT 45.040 245.620 47.710 247.000 ;
		END
	END PU
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			47.870 247.000 47.870 245.460
			44.880 245.460 44.880 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			47.910 247.000 47.910 245.420
			44.840 245.420 44.840 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			48.110 247.000 48.110 245.220
			44.640 245.220 44.640 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOCU12A

MACRO PBCSCTD8C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD8C

MACRO PBCSCTD8B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD8B

MACRO PBCSCTD8A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD8A

MACRO PBCSCTD4C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD4C

MACRO PBCSCTD4A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD4A

MACRO PBCSCTD2C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD2C

MACRO PBCSCTD2A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD2A

MACRO PBCSCTD24C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD24C

MACRO PBCSCTD24B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD24B

MACRO PBCSCTD24A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD24A

MACRO PBCSCTD16C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD16C

MACRO PBCSCTD16B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD16B

MACRO PBCSCTD16A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD16A

MACRO PBCSCTD12C
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD12C

MACRO PBCSCTD12B
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD12B

MACRO PBCSCTD12A
	CLASS PAD INOUT ;
	FOREIGN PBCSCTD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCTD12A

MACRO PBCCTD8C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD8C

MACRO PBCCTD8B
	CLASS PAD INOUT ;
	FOREIGN PBCCTD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD8B

MACRO PBCCTD8A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD8A

MACRO PBCCTD4C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD4C

MACRO PBCCTD4A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD4A

MACRO PBCCTD2C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD2C

MACRO PBCCTD2A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD2A

MACRO PBCCTD24C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD24C

MACRO PBCCTD24B
	CLASS PAD INOUT ;
	FOREIGN PBCCTD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD24B

MACRO PBCCTD24A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD24A

MACRO PBCCTD16C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD16C

MACRO PBCCTD16B
	CLASS PAD INOUT ;
	FOREIGN PBCCTD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD16B

MACRO PBCCTD16A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD16A

MACRO PBCCTD12C
	CLASS PAD INOUT ;
	FOREIGN PBCCTD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD12C

MACRO PBCCTD12B
	CLASS PAD INOUT ;
	FOREIGN PBCCTD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD12B

MACRO PBCCTD12A
	CLASS PAD INOUT ;
	FOREIGN PBCCTD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCTD12A

MACRO PBCSODD8C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD8C

MACRO PBCSODD8B
	CLASS PAD INOUT ;
	FOREIGN PBCSODD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD8B

MACRO PBCSODD8A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD8A

MACRO PBCSODD4C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD4C

MACRO PBCSODD4A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD4A

MACRO PBCSODD2C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD2C

MACRO PBCSODD2A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD2A

MACRO PBCSODD24C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD24C

MACRO PBCSODD24B
	CLASS PAD INOUT ;
	FOREIGN PBCSODD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD24B

MACRO PBCSODD24A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD24A

MACRO PBCSODD16C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD16C

MACRO PBCSODD16B
	CLASS PAD INOUT ;
	FOREIGN PBCSODD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD16B

MACRO PBCSODD16A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD16A

MACRO PBCSODD12C
	CLASS PAD INOUT ;
	FOREIGN PBCSODD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD12C

MACRO PBCSODD12B
	CLASS PAD INOUT ;
	FOREIGN PBCSODD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD12B

MACRO PBCSODD12A
	CLASS PAD INOUT ;
	FOREIGN PBCSODD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSODD12A

MACRO PBCODD8C
	CLASS PAD INOUT ;
	FOREIGN PBCODD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD8C

MACRO PBCODD8B
	CLASS PAD INOUT ;
	FOREIGN PBCODD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD8B

MACRO PBCODD8A
	CLASS PAD INOUT ;
	FOREIGN PBCODD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD8A

MACRO PBCODD4C
	CLASS PAD INOUT ;
	FOREIGN PBCODD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD4C

MACRO PBCODD4A
	CLASS PAD INOUT ;
	FOREIGN PBCODD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD4A

MACRO PBCODD2C
	CLASS PAD INOUT ;
	FOREIGN PBCODD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD2C

MACRO PBCODD2A
	CLASS PAD INOUT ;
	FOREIGN PBCODD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD2A

MACRO PBCODD24C
	CLASS PAD INOUT ;
	FOREIGN PBCODD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD24C

MACRO PBCODD24B
	CLASS PAD INOUT ;
	FOREIGN PBCODD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD24B

MACRO PBCODD24A
	CLASS PAD INOUT ;
	FOREIGN PBCODD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD24A

MACRO PBCODD16C
	CLASS PAD INOUT ;
	FOREIGN PBCODD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD16C

MACRO PBCODD16B
	CLASS PAD INOUT ;
	FOREIGN PBCODD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD16B

MACRO PBCODD16A
	CLASS PAD INOUT ;
	FOREIGN PBCODD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD16A

MACRO PBCODD12C
	CLASS PAD INOUT ;
	FOREIGN PBCODD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD12C

MACRO PBCODD12B
	CLASS PAD INOUT ;
	FOREIGN PBCODD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD12B

MACRO PBCODD12A
	CLASS PAD INOUT ;
	FOREIGN PBCODD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN PD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER MQ ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M6 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M5 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M4 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M3 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M2 ;
			RECT 48.310 245.620 50.980 247.000 ;
			LAYER M1 ;
			RECT 48.310 245.620 50.980 247.000 ;
		END
	END PD
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			51.140 247.000 51.140 245.460
			48.150 245.460 48.150 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			48.110 245.420 48.110 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			47.910 245.220 47.910 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCODD12A

MACRO PBCSCT8C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT8C

MACRO PBCSCT8B
	CLASS PAD INOUT ;
	FOREIGN PBCSCT8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT8B

MACRO PBCSCT8A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT8A

MACRO PBCSCT4C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT4C

MACRO PBCSCT4A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT4A

MACRO PBCSCT2C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT2C

MACRO PBCSCT2A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT2A

MACRO PBCSCT24C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT24C

MACRO PBCSCT24B
	CLASS PAD INOUT ;
	FOREIGN PBCSCT24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT24B

MACRO PBCSCT24A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT24A

MACRO PBCSCT16C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT16C

MACRO PBCSCT16B
	CLASS PAD INOUT ;
	FOREIGN PBCSCT16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT16B

MACRO PBCSCT16A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT16A

MACRO PBCSCT12C
	CLASS PAD INOUT ;
	FOREIGN PBCSCT12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT12C

MACRO PBCSCT12B
	CLASS PAD INOUT ;
	FOREIGN PBCSCT12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT12B

MACRO PBCSCT12A
	CLASS PAD INOUT ;
	FOREIGN PBCSCT12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSCT12A

MACRO PBCCT8C
	CLASS PAD INOUT ;
	FOREIGN PBCCT8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT8C

MACRO PBCCT8B
	CLASS PAD INOUT ;
	FOREIGN PBCCT8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT8B

MACRO PBCCT8A
	CLASS PAD INOUT ;
	FOREIGN PBCCT8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT8A

MACRO PBCCT4C
	CLASS PAD INOUT ;
	FOREIGN PBCCT4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT4C

MACRO PBCCT4A
	CLASS PAD INOUT ;
	FOREIGN PBCCT4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT4A

MACRO PBCCT2C
	CLASS PAD INOUT ;
	FOREIGN PBCCT2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT2C

MACRO PBCCT2A
	CLASS PAD INOUT ;
	FOREIGN PBCCT2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT2A

MACRO PBCCT24C
	CLASS PAD INOUT ;
	FOREIGN PBCCT24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT24C

MACRO PBCCT24B
	CLASS PAD INOUT ;
	FOREIGN PBCCT24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT24B

MACRO PBCCT24A
	CLASS PAD INOUT ;
	FOREIGN PBCCT24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT24A

MACRO PBCCT16C
	CLASS PAD INOUT ;
	FOREIGN PBCCT16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT16C

MACRO PBCCT16B
	CLASS PAD INOUT ;
	FOREIGN PBCCT16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT16B

MACRO PBCCT16A
	CLASS PAD INOUT ;
	FOREIGN PBCCT16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT16A

MACRO PBCCT12C
	CLASS PAD INOUT ;
	FOREIGN PBCCT12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT12C

MACRO PBCCT12B
	CLASS PAD INOUT ;
	FOREIGN PBCCT12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT12B

MACRO PBCCT12A
	CLASS PAD INOUT ;
	FOREIGN PBCCT12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCCT12A

MACRO PBCSOD8C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD8C

MACRO PBCSOD8B
	CLASS PAD INOUT ;
	FOREIGN PBCSOD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD8B

MACRO PBCSOD8A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD8A

MACRO PBCSOD4C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD4C

MACRO PBCSOD4A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD4A

MACRO PBCSOD2C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD2C

MACRO PBCSOD2A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD2A

MACRO PBCSOD24C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD24C

MACRO PBCSOD24B
	CLASS PAD INOUT ;
	FOREIGN PBCSOD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD24B

MACRO PBCSOD24A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD24A

MACRO PBCSOD16C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD16C

MACRO PBCSOD16B
	CLASS PAD INOUT ;
	FOREIGN PBCSOD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD16B

MACRO PBCSOD16A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD16A

MACRO PBCSOD12C
	CLASS PAD INOUT ;
	FOREIGN PBCSOD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD12C

MACRO PBCSOD12B
	CLASS PAD INOUT ;
	FOREIGN PBCSOD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD12B

MACRO PBCSOD12A
	CLASS PAD INOUT ;
	FOREIGN PBCSOD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOD12A

MACRO PBCOD8C
	CLASS PAD INOUT ;
	FOREIGN PBCOD8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD8C

MACRO PBCOD8B
	CLASS PAD INOUT ;
	FOREIGN PBCOD8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD8B

MACRO PBCOD8A
	CLASS PAD INOUT ;
	FOREIGN PBCOD8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD8A

MACRO PBCOD4C
	CLASS PAD INOUT ;
	FOREIGN PBCOD4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD4C

MACRO PBCOD4A
	CLASS PAD INOUT ;
	FOREIGN PBCOD4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD4A

MACRO PBCOD2C
	CLASS PAD INOUT ;
	FOREIGN PBCOD2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD2C

MACRO PBCOD2A
	CLASS PAD INOUT ;
	FOREIGN PBCOD2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD2A

MACRO PBCOD24C
	CLASS PAD INOUT ;
	FOREIGN PBCOD24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD24C

MACRO PBCOD24B
	CLASS PAD INOUT ;
	FOREIGN PBCOD24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD24B

MACRO PBCOD24A
	CLASS PAD INOUT ;
	FOREIGN PBCOD24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD24A

MACRO PBCOD16C
	CLASS PAD INOUT ;
	FOREIGN PBCOD16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD16C

MACRO PBCOD16B
	CLASS PAD INOUT ;
	FOREIGN PBCOD16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD16B

MACRO PBCOD16A
	CLASS PAD INOUT ;
	FOREIGN PBCOD16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD16A

MACRO PBCOD12C
	CLASS PAD INOUT ;
	FOREIGN PBCOD12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD12C

MACRO PBCOD12B
	CLASS PAD INOUT ;
	FOREIGN PBCOD12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD12B

MACRO PBCOD12A
	CLASS PAD INOUT ;
	FOREIGN PBCOD12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOD12A

MACRO PBCSOC8C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC8C

MACRO PBCSOC8B
	CLASS PAD INOUT ;
	FOREIGN PBCSOC8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC8B

MACRO PBCSOC8A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC8A

MACRO PBCSOC4C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC4C

MACRO PBCSOC4A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC4A

MACRO PBCSOC2C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC2C

MACRO PBCSOC2A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC2A

MACRO PBCSOC24C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC24C

MACRO PBCSOC24B
	CLASS PAD INOUT ;
	FOREIGN PBCSOC24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC24B

MACRO PBCSOC24A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC24A

MACRO PBCSOC16C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC16C

MACRO PBCSOC16B
	CLASS PAD INOUT ;
	FOREIGN PBCSOC16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC16B

MACRO PBCSOC16A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC16A

MACRO PBCSOC12C
	CLASS PAD INOUT ;
	FOREIGN PBCSOC12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC12C

MACRO PBCSOC12B
	CLASS PAD INOUT ;
	FOREIGN PBCSOC12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC12B

MACRO PBCSOC12A
	CLASS PAD INOUT ;
	FOREIGN PBCSOC12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCSOC12A

MACRO PBCOC8C
	CLASS PAD INOUT ;
	FOREIGN PBCOC8C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC8C

MACRO PBCOC8B
	CLASS PAD INOUT ;
	FOREIGN PBCOC8B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC8B

MACRO PBCOC8A
	CLASS PAD INOUT ;
	FOREIGN PBCOC8A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC8A

MACRO PBCOC4C
	CLASS PAD INOUT ;
	FOREIGN PBCOC4C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC4C

MACRO PBCOC4A
	CLASS PAD INOUT ;
	FOREIGN PBCOC4A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC4A

MACRO PBCOC2C
	CLASS PAD INOUT ;
	FOREIGN PBCOC2C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC2C

MACRO PBCOC2A
	CLASS PAD INOUT ;
	FOREIGN PBCOC2A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC2A

MACRO PBCOC24C
	CLASS PAD INOUT ;
	FOREIGN PBCOC24C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC24C

MACRO PBCOC24B
	CLASS PAD INOUT ;
	FOREIGN PBCOC24B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC24B

MACRO PBCOC24A
	CLASS PAD INOUT ;
	FOREIGN PBCOC24A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC24A

MACRO PBCOC16C
	CLASS PAD INOUT ;
	FOREIGN PBCOC16C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC16C

MACRO PBCOC16B
	CLASS PAD INOUT ;
	FOREIGN PBCOC16B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC16B

MACRO PBCOC16A
	CLASS PAD INOUT ;
	FOREIGN PBCOC16A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC16A

MACRO PBCOC12C
	CLASS PAD INOUT ;
	FOREIGN PBCOC12C 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC12C

MACRO PBCOC12B
	CLASS PAD INOUT ;
	FOREIGN PBCOC12B 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC12B

MACRO PBCOC12A
	CLASS PAD INOUT ;
	FOREIGN PBCOC12A 0 0 ;
	ORIGIN 0 0 ;
	SIZE 70.000 BY 247.000 ;
	SYMMETRY X Y R90 ;
	SITE iosite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER MQ ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M6 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M5 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M4 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M3 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M2 ;
			RECT 61.390 245.620 64.060 247.000 ;
			LAYER M1 ;
			RECT 61.390 245.620 64.060 247.000 ;
		END
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER MQ ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M6 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M5 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M4 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M3 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M2 ;
			RECT 58.120 245.620 60.790 247.000 ;
			LAYER M1 ;
			RECT 58.120 245.620 60.790 247.000 ;
		END
	END A
	PIN P
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER LM ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER MQ ;
			RECT 6.000 104.500 64.000 114.000 ;
			LAYER M6 ;
			RECT 6.000 104.500 64.000 114.000 ;
		END
	END P
	PIN IE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER MQ ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M6 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M5 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M4 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M3 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M2 ;
			RECT 51.580 245.620 54.250 247.000 ;
			LAYER M1 ;
			RECT 51.580 245.620 54.250 247.000 ;
		END
	END IE
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			CLASS CORE ;
			LAYER LM ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER MQ ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M6 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M5 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M4 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M3 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M2 ;
			RECT 54.850 245.620 57.520 247.000 ;
			LAYER M1 ;
			RECT 54.850 245.620 57.520 247.000 ;
		END
	END OE
	OBS
		LAYER M1 ;
		POLYGON 0.080 0.000 69.920 0.000 69.920 246.840
			69.840 246.840 
			69.840 247.000 
			64.220 247.000
			64.220 245.460
			61.230 245.460 61.230 247.000
			60.950 247.000 60.950 245.460
			57.960 245.460 57.960 247.000
			57.680 247.000 57.680 245.460
			54.690 245.460 54.690 247.000
			54.410 247.000 54.410 245.460
			51.420 245.460 51.420 247.000
			0.160 247.000 0.160 246.840 0.080 246.840
			0.080 0.000 ;
		LAYER M2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V1 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V2 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V3 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V4 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER M6 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 
			69.800 247.000 
			64.260 247.000
			64.260 245.420
			51.380 245.420 51.380 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER V5 ;
		POLYGON 0.100 0.000 69.900 0.000 69.900 246.800
			69.800 246.800 69.800 247.000
			0.200 247.000 0.200 246.800 0.100 246.800
			0.100 0.000 ;
		LAYER MQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VL ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER LM ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 
			69.600 247.000 
			64.460 247.000
			64.460 245.220
			51.180 245.220 51.180 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
		LAYER VQ ;
		POLYGON 0.200 0.000 69.800 0.000 69.800 246.600
			69.600 246.600 69.600 247.000
			0.400 247.000 0.400 246.600 0.200 246.600
			0.200 0.000 ;
END
END PBCOC12A

END LIBRARY
