
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.3.58
#
# REF LIBS: lab3 
# TECH LIB NAME: cmrf8sf
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.010000 ;

MACRO reset_driver
    CLASS BLOCK ;
    FOREIGN reset_driver 0 -0.28 ;
    ORIGIN 0.000 0.280 ;
    SIZE 11.190 BY 4.160 ;
    SYMMETRY X Y R90 ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.470 0.680 1.750 ;
        RECT  0.080 1.240 0.400 1.750 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.830 1.240 10.550 1.960 ;
        RECT  9.990 0.440 10.270 3.080 ;
        RECT  9.830 1.240 10.270 1.970 ;
        RECT  9.030 0.440 9.310 0.720 ;
        RECT  9.030 2.800 9.310 3.080 ;
        RECT  8.070 0.440 8.350 0.720 ;
        RECT  8.070 2.800 8.350 3.080 ;
        RECT  7.110 0.650 7.390 0.930 ;
        RECT  7.110 2.800 7.390 3.080 ;
        END
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 11.190 0.280 ;
        RECT  10.470 -0.280 10.750 0.680 ;
        RECT  9.510 -0.280 9.790 0.670 ;
        RECT  8.550 -0.280 8.830 0.670 ;
        RECT  7.590 -0.280 7.870 0.670 ;
        RECT  6.630 -0.280 7.870 0.340 ;
        RECT  6.630 -0.280 6.910 0.990 ;
        RECT  5.540 -0.280 5.820 0.870 ;
        RECT  4.540 -0.280 5.820 0.340 ;
        RECT  4.540 -0.280 4.820 0.400 ;
        RECT  3.540 -0.280 3.820 1.030 ;
        RECT  2.590 -0.280 2.870 0.860 ;
        RECT  1.630 -0.280 1.910 0.920 ;
        RECT  0.160 -0.280 0.440 0.990 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 11.190 3.880 ;
        RECT  10.470 2.310 10.750 3.880 ;
        RECT  9.510 2.340 9.790 3.880 ;
        RECT  8.550 2.340 8.830 3.880 ;
        RECT  7.590 2.330 7.870 3.880 ;
        RECT  6.630 1.910 6.910 3.880 ;
        RECT  5.460 1.970 5.740 3.880 ;
        RECT  4.500 2.520 4.780 3.880 ;
        RECT  3.540 2.240 3.820 3.880 ;
        RECT  2.680 2.420 2.960 3.880 ;
        RECT  1.630 2.530 1.910 3.880 ;
        RECT  0.160 2.750 0.440 3.880 ;
        END
    END VDD
    OBS
        LAYER PC ;
        RECT  0.440 1.510 0.640 1.710 ;
        RECT  0.520 0.160 0.640 3.420 ;
        RECT  1.950 1.510 2.550 1.710 ;
        RECT  2.430 0.270 2.550 3.310 ;
        RECT  1.950 0.270 2.070 3.440 ;
        RECT  4.900 0.160 5.020 1.540 ;
        RECT  5.380 0.420 5.500 1.540 ;
        RECT  3.860 1.420 5.500 1.540 ;
        RECT  3.860 1.400 4.940 1.600 ;
        RECT  5.300 1.420 5.420 3.260 ;
        RECT  3.860 0.160 3.980 3.440 ;
        RECT  4.340 0.160 4.460 3.440 ;
        RECT  4.820 1.400 4.940 3.440 ;
        RECT  6.360 1.420 10.430 1.540 ;
        RECT  6.360 1.400 9.470 1.600 ;
        RECT  6.950 0.420 7.070 3.310 ;
        RECT  7.430 0.160 7.550 3.430 ;
        RECT  7.910 0.160 8.030 3.430 ;
        RECT  8.390 0.160 8.510 3.430 ;
        RECT  8.870 0.160 8.990 3.430 ;
        RECT  9.350 0.160 9.470 3.430 ;
        RECT  9.830 0.160 9.950 3.430 ;
        RECT  10.310 0.160 10.430 3.430 ;
        LAYER M1 ;
        RECT  0.680 0.440 1.000 1.310 ;
        RECT  0.840 1.470 2.190 1.750 ;
        RECT  0.840 1.240 1.120 2.360 ;
        RECT  1.620 1.470 1.900 2.360 ;
        RECT  0.680 1.910 0.960 3.160 ;
        RECT  2.110 0.650 2.390 1.310 ;
        RECT  2.110 1.120 2.660 1.310 ;
        RECT  2.420 1.240 4.610 1.550 ;
        RECT  3.530 1.240 4.610 1.640 ;
        RECT  3.530 1.240 3.770 1.960 ;
        RECT  2.420 1.120 2.660 2.170 ;
        RECT  2.110 1.910 2.660 2.170 ;
        RECT  2.110 1.910 2.390 3.080 ;
        RECT  4.020 0.600 5.340 1.080 ;
        RECT  6.660 1.240 6.950 1.640 ;
        RECT  4.930 1.390 6.950 1.640 ;
        RECT  4.930 1.040 5.570 1.810 ;
        RECT  4.020 1.800 5.300 2.280 ;
        RECT  4.980 0.600 5.300 2.890 ;
        RECT  4.020 1.800 4.300 3.160 ;
    END
END reset_driver

END LIBRARY
