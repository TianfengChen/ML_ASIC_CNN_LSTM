

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO Main_controller 
  PIN clk 
    ANTENNAPARTIALMETALAREA 7.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.075 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8352 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.44732 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0952826 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0957854 LAYER V3 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 27.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 14.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1416 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.932 LAYER M4 ; 
    ANTENNAMAXAREACAR 25.2218 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.252442 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.01838 LAYER V4 ;
  END reset
  PIN wrb 
    ANTENNAPARTIALMETALAREA 10.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1078 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1616 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2088 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.9899 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.229167 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER V4 ;
  END wrb
  PIN PE_state[2] 
    ANTENNAPARTIALMETALAREA 14.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1422 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.172 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1128 LAYER M3 ;
  END PE_state[2]
  PIN PE_state[1] 
    ANTENNAPARTIALMETALAREA 12.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.196 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1456 LAYER M3 ;
  END PE_state[1]
  PIN PE_state[0] 
    ANTENNAPARTIALMETALAREA 13.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.378 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1552 LAYER M3 ;
  END PE_state[0]
  PIN wrb_addr[7] 
    ANTENNAPARTIALMETALAREA 4.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0414 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4824 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.5562 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.153255 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V3 ;
  END wrb_addr[7]
  PIN wrb_addr[6] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.42 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.979 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.121749 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.765189 LAYER V3 ;
  END wrb_addr[6]
  PIN wrb_addr[5] 
    ANTENNADIFFAREA 2.014 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.7051 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.208333 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.93633 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M3 ;
    ANTENNAGATEAREA 0.4464 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.1101 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.244176 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V3 ;
  END wrb_addr[5]
  PIN wrb_addr[4] 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.132 LAYER M2 ; 
    ANTENNAMAXAREACAR 15.0939 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.151364 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.909091 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0256 LAYER M3 ;
    ANTENNAGATEAREA 0.2952 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.495 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.238085 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.49649 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0128 LAYER M4 ;
    ANTENNAGATEAREA 0.5208 LAYER M4 ; 
    ANTENNAMAXAREACAR 25.876 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.262662 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.63854 LAYER V4 ;
  END wrb_addr[4]
  PIN wrb_addr[3] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M2 ; 
    ANTENNAMAXAREACAR 53.6782 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.537069 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0208 LAYER M3 ;
    ANTENNAGATEAREA 0.4152 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.5915 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.587165 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.91682 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0248 LAYER M4 ;
    ANTENNAGATEAREA 0.684 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.1587 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.623423 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.91682 LAYER V4 ;
  END wrb_addr[3]
  PIN wrb_addr[2] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.0163 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.144202 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.857199 LAYER V3 ;
  END wrb_addr[2]
  PIN wrb_addr[1] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.027 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3336 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.3925 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.137809 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.814521 LAYER V3 ;
  END wrb_addr[1]
  PIN wrb_addr[0] 
    ANTENNAPARTIALMETALAREA 4.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2256 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.2724 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.532477 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.65346 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M4 ;
    ANTENNAGATEAREA 0.5616 LAYER M4 ; 
    ANTENNAMAXAREACAR 53.9106 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.549571 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.65346 LAYER V4 ;
  END wrb_addr[0]
  PIN rdB_addr[3] 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.75 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0808 LAYER M3 ;
  END rdB_addr[3]
  PIN rdB_addr[2] 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.56 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0552 LAYER M3 ;
  END rdB_addr[2]
  PIN rdB_addr[1] 
    ANTENNAPARTIALMETALAREA 8.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.083 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 8.58 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4848 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.087 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.209418 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.632911 LAYER V3 ;
  END rdB_addr[1]
  PIN rdB_addr[0] 
    ANTENNAPARTIALMETALAREA 8.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.112 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.7611 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.47298 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V3 ;
  END rdB_addr[0]
  PIN mem_addr[12] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.3303 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.209715 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.94308 LAYER V3 ;
  END mem_addr[12]
  PIN mem_addr[11] 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0494 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 LAYER M2 ; 
    ANTENNAMAXAREACAR 28.366 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.28412 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.54625 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M3 ;
    ANTENNAGATEAREA 0.2016 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.323803 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.54625 LAYER V3 ;
  END mem_addr[11]
  PIN mem_addr[10] 
    ANTENNAPARTIALMETALAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0296 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 LAYER M2 ; 
    ANTENNAMAXAREACAR 12.5393 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.124365 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.822535 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.4884 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.273374 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[10]
  PIN mem_addr[9] 
    ANTENNAPARTIALMETALAREA 4.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.043 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 LAYER M2 ; 
    ANTENNAMAXAREACAR 17.3114 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.172086 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.822535 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.8416 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.346906 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[9]
  PIN mem_addr[8] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0224 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5808 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.1148 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.224186 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END mem_addr[8]
  PIN mem_addr[7] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.6908 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.176539 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[7]
  PIN mem_addr[6] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.4567 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.20882 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END mem_addr[6]
  PIN mem_addr[5] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0198 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M2 ; 
    ANTENNAMAXAREACAR 15.3044 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.152016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0352 LAYER M3 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.5875 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.484365 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[5]
  PIN mem_addr[4] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0304 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.432 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.393 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.34994 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END mem_addr[4]
  PIN mem_addr[3] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.0441 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.183121 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END mem_addr[3]
  PIN mem_addr[2] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0198 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.7939 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.33655 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[2]
  PIN mem_addr[1] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M2 ; 
    ANTENNAMAXAREACAR 16.4778 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.165323 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.806452 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0216 LAYER M3 ;
    ANTENNAGATEAREA 0.3504 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.8096 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.376586 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END mem_addr[1]
  PIN mem_addr[0] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.5894 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.180242 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0352 LAYER M4 ;
    ANTENNAGATEAREA 0.504 LAYER M4 ; 
    ANTENNAMAXAREACAR 24.4941 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.250083 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.52408 LAYER V4 ;
  END mem_addr[0]
  PIN SRAM_in_A_addr[9] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0918 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6648 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.6225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.330814 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.12121 LAYER V3 ;
  END SRAM_in_A_addr[9]
  PIN SRAM_in_A_addr[8] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0934 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6144 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.3121 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.272852 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER V3 ;
  END SRAM_in_A_addr[8]
  PIN SRAM_in_A_addr[7] 
    ANTENNAPARTIALMETALAREA 12.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4752 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.8714 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.310374 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.24362 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0368 LAYER M4 ;
    ANTENNAGATEAREA 1.3176 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.634 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.338303 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.53568 LAYER V4 ;
  END SRAM_in_A_addr[7]
  PIN SRAM_in_A_addr[6] 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0494 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0344 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4304 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.6146 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.464998 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.9639 LAYER V4 ;
  END SRAM_in_A_addr[6]
  PIN SRAM_in_A_addr[5] 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0566 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1024 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0616 LAYER M4 ; 
    ANTENNAMAXAREACAR 29.8738 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.307735 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.96078 LAYER V4 ;
  END SRAM_in_A_addr[5]
  PIN SRAM_in_A_addr[4] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.119 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.54 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.4508 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.300543 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V3 ;
  END SRAM_in_A_addr[4]
  PIN SRAM_in_A_addr[3] 
    ANTENNADIFFAREA 4.168 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1438 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.3946 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.310621 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.85234 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M4 ;
    ANTENNAGATEAREA 0.7824 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.3659 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.320846 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.85234 LAYER V4 ;
  END SRAM_in_A_addr[3]
  PIN SRAM_in_A_addr[2] 
    ANTENNADIFFAREA 4.168 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1502 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9312 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1379 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.236171 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.00899 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M4 ;
    ANTENNAGATEAREA 1.2192 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.0447 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.315567 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.65873 LAYER V4 ;
  END SRAM_in_A_addr[2]
  PIN SRAM_in_A_addr[1] 
    ANTENNADIFFAREA 4.168 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.124 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3912 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5277 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.427609 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.983711 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0232 LAYER M4 ;
    ANTENNAGATEAREA 1.3512 LAYER M4 ; 
    ANTENNAMAXAREACAR 44.1855 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.444779 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.46248 LAYER V4 ;
  END SRAM_in_A_addr[1]
  PIN SRAM_in_A_addr[0] 
    ANTENNAPARTIALMETALAREA 8.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.083 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3216 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.8917 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316867 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.641952 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0528 LAYER M4 ;
    ANTENNAGATEAREA 1.2504 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.0823 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.359094 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.31444 LAYER V4 ;
  END SRAM_in_A_addr[0]
  PIN SRAM_in_B_addr[9] 
    ANTENNAPARTIALMETALAREA 4.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0494 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5208 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.2374 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.180612 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.69207 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M4 ;
    ANTENNAGATEAREA 0.8016 LAYER M4 ; 
    ANTENNAMAXAREACAR 19.9839 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.198576 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.69207 LAYER V4 ;
  END SRAM_in_B_addr[9]
  PIN SRAM_in_B_addr[8] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0486 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2328 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4328 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.276357 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.46248 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0224 LAYER M4 ;
    ANTENNAGATEAREA 0.5976 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.1142 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.31384 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.94344 LAYER V4 ;
  END SRAM_in_B_addr[8]
  PIN SRAM_in_B_addr[7] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0526 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6528 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.3543 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.208662 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.6377 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0104 LAYER M4 ;
    ANTENNAGATEAREA 0.7224 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.7386 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.223059 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V4 ;
  END SRAM_in_B_addr[7]
  PIN SRAM_in_B_addr[6] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.075 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6816 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.5212 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.202229 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END SRAM_in_B_addr[6]
  PIN SRAM_in_B_addr[5] 
    ANTENNAPARTIALMETALAREA 5.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0534 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5208 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6761 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.26982 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.03564 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M4 ;
    ANTENNAGATEAREA 0.6504 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.8446 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.28212 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.16049 LAYER V4 ;
  END SRAM_in_B_addr[5]
  PIN SRAM_in_B_addr[4] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.055 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.1858 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.239644 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END SRAM_in_B_addr[4]
  PIN SRAM_in_B_addr[3] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0614 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4272 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.921 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.21729 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V3 ;
  END SRAM_in_B_addr[3]
  PIN SRAM_in_B_addr[2] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0968 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.7034 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.30397 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.44828 LAYER V3 ;
  END SRAM_in_B_addr[2]
  PIN SRAM_in_B_addr[1] 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0606 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.056 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3212 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.185973 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.76671 LAYER V3 ;
  END SRAM_in_B_addr[1]
  PIN SRAM_in_B_addr[0] 
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1134 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2096 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.4371 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.452083 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V3 ;
  END SRAM_in_B_addr[0]
  PIN SRAM_WENB1 
    ANTENNAPARTIALMETALAREA 5.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0534 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.33125 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V3 ;
    ANTENNADIFFAREA 2.848 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0248 LAYER M4 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 46.7083 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.474769 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END SRAM_WENB1
  PIN SRAM_WENB2 
    ANTENNADIFFAREA 2.848 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.055 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3456 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.6412 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.226042 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END SRAM_WENB2
  PIN SRAM_WENB3 
    ANTENNADIFFAREA 2.848 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3456 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.1713 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.225926 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V3 ;
  END SRAM_WENB3
  PIN SRAM_WENB4 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.4213 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.327315 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V3 ;
    ANTENNADIFFAREA 2.848 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0752 LAYER M4 ;
    ANTENNAGATEAREA 0.42 LAYER M4 ; 
    ANTENNAMAXAREACAR 50.1356 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.506362 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.68817 LAYER V4 ;
  END SRAM_WENB4
END Main_controller

END LIBRARY
