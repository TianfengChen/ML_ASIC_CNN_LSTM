

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO CNN_controller 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0142 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8352 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.45498 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0253592 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.191571 LAYER V3 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 11.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1142 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.408 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.0493 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.309755 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.392157 LAYER V3 ;
  END reset
  PIN PE_state[2] 
    ANTENNAPARTIALMETALAREA 9.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0918 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.576 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.12 LAYER M3 ;
  END PE_state[2]
  PIN PE_state[1] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.047 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.172 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 11.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1168 LAYER M3 ;
  END PE_state[1]
  PIN PE_state[0] 
    ANTENNAPARTIALMETALAREA 6.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0686 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1432 LAYER M3 ;
  END PE_state[0]
  PIN wrb_addr[7] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5208 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.0546 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.234909 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V3 ;
  END wrb_addr[7]
  PIN wrb_addr[6] 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7968 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.3286 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.260826 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER V3 ;
  END wrb_addr[6]
  PIN wrb_addr[5] 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5592 LAYER M4 ; 
    ANTENNAMAXAREACAR 10.8714 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.112327 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.05215 LAYER V4 ;
  END wrb_addr[5]
  PIN wrb_addr[4] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1056 LAYER M2 ; 
    ANTENNAMAXAREACAR 30.8977 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.308902 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.89394 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M3 ;
    ANTENNAGATEAREA 0.1056 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.2917 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.460417 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.65152 LAYER V3 ;
    ANTENNADIFFAREA 3.488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0072 LAYER M4 ;
    ANTENNAGATEAREA 0.5568 LAYER M4 ; 
    ANTENNAMAXAREACAR 46.5129 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.473348 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.65152 LAYER V4 ;
  END wrb_addr[4]
  PIN wrb_addr[3] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.4368 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.364655 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAGATEAREA 0.3912 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6863 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.389195 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.25167 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M4 ;
    ANTENNAGATEAREA 0.564 LAYER M4 ; 
    ANTENNAMAXAREACAR 39.4664 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.397706 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.25167 LAYER V4 ;
  END wrb_addr[3]
  PIN wrb_addr[2] 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3216 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.39428 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0986526 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER V3 ;
  END wrb_addr[2]
  PIN wrb_addr[1] 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0334 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4272 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.67823 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.086064 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.490296 LAYER V3 ;
  END wrb_addr[1]
  PIN wrb_addr[0] 
    ANTENNAPARTIALMETALAREA 4.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0462 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4272 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.84898 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0997301 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.677462 LAYER V3 ;
  END wrb_addr[0]
  PIN wrb 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2056 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M4 ; 
    ANTENNAMAXAREACAR 19.0197 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.197097 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.93633 LAYER V4 ;
  END wrb
  PIN rdB_addr[3] 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.94 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0384 LAYER M3 ;
  END rdB_addr[3]
  PIN rdB_addr[2] 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.039 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 8.294 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.4722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.41713 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V3 ;
  END rdB_addr[2]
  PIN rdB_addr[1] 
    ANTENNAPARTIALMETALAREA 7.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0742 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 4.2 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3072 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.0685 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.375244 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.70068 LAYER V3 ;
  END rdB_addr[1]
  PIN rdB_addr[0] 
    ANTENNAPARTIALMETALAREA 6.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0662 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.816 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4224 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.2294 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.320169 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.70068 LAYER V3 ;
  END rdB_addr[0]
  PIN mem_addr1[15] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.612 LAYER M4 ; 
    ANTENNAMAXAREACAR 22.4982 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.228243 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.4328 LAYER V4 ;
  END mem_addr1[15]
  PIN mem_addr1[14] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 4.168 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 30.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4656 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.2021 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.736226 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.978273 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M4 ;
    ANTENNAGATEAREA 0.7752 LAYER M4 ; 
    ANTENNAMAXAREACAR 74.5953 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.750674 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.16749 LAYER V4 ;
  END mem_addr1[14]
  PIN mem_addr1[13] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 28.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5808 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.5926 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.591446 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.65289 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0176 LAYER M4 ;
    ANTENNAGATEAREA 0.8208 LAYER M4 ; 
    ANTENNAMAXAREACAR 60.6881 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.612889 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.71429 LAYER V4 ;
  END mem_addr1[13]
  PIN mem_addr1[12] 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2416 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7944 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.0474 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.466949 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.66667 LAYER V3 ;
  END mem_addr1[12]
  PIN mem_addr1[11] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 3.488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 22.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.84 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.3942 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.511321 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.66667 LAYER V3 ;
  END mem_addr1[11]
  PIN mem_addr1[10] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3696 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.602 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.541962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.43867 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0296 LAYER M4 ;
    ANTENNAGATEAREA 0.8784 LAYER M4 ; 
    ANTENNAMAXAREACAR 56.9262 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.57566 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.43867 LAYER V4 ;
  END mem_addr1[10]
  PIN mem_addr1[9] 
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.176 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1448 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9048 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.5729 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.228924 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER V3 ;
  END mem_addr1[9]
  PIN mem_addr1[8] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.176 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0008 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0562 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.361028 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.73993 LAYER V3 ;
  END mem_addr1[8]
  PIN mem_addr1[7] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 35.869 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.363038 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0344 LAYER M4 ;
    ANTENNAGATEAREA 1.1928 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.6523 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.391877 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.84615 LAYER V4 ;
  END mem_addr1[7]
  PIN mem_addr1[6] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M2 ; 
    ANTENNAMAXAREACAR 17.5531 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.176075 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.806452 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0576 LAYER M3 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.994 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.563172 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0104 LAYER M4 ;
    ANTENNAGATEAREA 0.852 LAYER M4 ; 
    ANTENNAMAXAREACAR 57.1677 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.575379 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V4 ;
  END mem_addr1[6]
  PIN mem_addr1[5] 
    ANTENNADIFFAREA 2.176 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.059 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER V2 ;
    ANTENNADIFFAREA 2.176 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9504 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.3666 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.179482 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.0202 LAYER V3 ;
  END mem_addr1[5]
  PIN mem_addr1[4] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0318 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.072 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.4667 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.458889 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 1.66667 LAYER V2 ;
    ANTENNADIFFAREA 2.176 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0448 LAYER M3 ;
    ANTENNAGATEAREA 0.4752 LAYER M3 ; 
    ANTENNAMAXAREACAR 54.6418 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.553165 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.06229 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0416 LAYER M4 ;
    ANTENNAGATEAREA 0.648 LAYER M4 ; 
    ANTENNAMAXAREACAR 60.9998 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.617363 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.06229 LAYER V4 ;
  END mem_addr1[4]
  PIN mem_addr1[3] 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7248 LAYER M4 ; 
    ANTENNAMAXAREACAR 32.3405 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.326721 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.72328 LAYER V4 ;
  END mem_addr1[3]
  PIN mem_addr1[2] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0808 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.66 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.4457 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.377935 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.73412 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0328 LAYER M4 ;
    ANTENNAGATEAREA 1.14 LAYER M4 ; 
    ANTENNAMAXAREACAR 40.2878 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.406707 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.73412 LAYER V4 ;
  END mem_addr1[2]
  PIN mem_addr1[1] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0608 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6858 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.390655 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.75535 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.044 LAYER M4 ;
    ANTENNAGATEAREA 0.9696 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.1412 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.436034 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.75535 LAYER V4 ;
  END mem_addr1[1]
  PIN mem_addr1[0] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 21.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2176 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7464 LAYER M4 ; 
    ANTENNAMAXAREACAR 59.4246 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.60234 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V4 ;
  END mem_addr1[0]
  PIN mem_addr2[15] 
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.3565 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.421875 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END mem_addr2[15]
  PIN mem_addr2[14] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0512 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0744 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 53.8565 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.546875 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END mem_addr2[14]
  PIN mem_addr2[13] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0504 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 46.6806 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.477431 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END mem_addr2[13]
  PIN mem_addr2[12] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.9861 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.468171 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END mem_addr2[12]
  PIN mem_addr2[11] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 24.4583 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.255208 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END mem_addr2[11]
  PIN mem_addr2[10] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0608 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.3807 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.660201 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V4 ;
  END mem_addr2[10]
  PIN mem_addr2[9] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.96 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 14.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1408 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.132 LAYER M4 ; 
    ANTENNAMAXAREACAR 152.162 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.52818 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.42424 LAYER V4 ;
  END mem_addr2[9]
  PIN mem_addr2[8] 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0424 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0704 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 61.4954 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.625579 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END mem_addr2[8]
  PIN mem_addr2[7] 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.17 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.658737 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V4 ;
  END mem_addr2[7]
  PIN mem_addr2[6] 
    ANTENNAPARTIALMETALAREA 7.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0774 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 93.6647 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.943683 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER V3 ;
  END mem_addr2[6]
  PIN mem_addr2[5] 
    ANTENNAPARTIALMETALAREA 6.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0654 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 17.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.457 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.12998 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER V3 ;
  END mem_addr2[5]
  PIN mem_addr2[4] 
    ANTENNAPARTIALMETALAREA 8.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0846 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1552 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.132 LAYER M4 ; 
    ANTENNAMAXAREACAR 18.8818 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.201364 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.21212 LAYER V4 ;
  END mem_addr2[4]
  PIN mem_addr2[3] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0416 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M4 ; 
    ANTENNAMAXAREACAR 93.1034 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.951724 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER V4 ;
  END mem_addr2[3]
  PIN mem_addr2[2] 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.132 LAYER M4 ; 
    ANTENNAMAXAREACAR 83.4273 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.843788 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.51515 LAYER V4 ;
  END mem_addr2[2]
  PIN mem_addr2[1] 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1912 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 17.3206 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.185618 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V4 ;
  END mem_addr2[1]
  PIN mem_addr2[0] 
    ANTENNAPARTIALMETALAREA 21.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.7097 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.471505 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER V4 ;
  END mem_addr2[0]
  PIN SRAM_in_A_addr[9] 
    ANTENNADIFFAREA 2.176 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0486 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8568 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.1214 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.24621 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.05128 LAYER V3 ;
  END SRAM_in_A_addr[9]
  PIN SRAM_in_A_addr[8] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0414 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5399 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.160283 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.1057 LAYER V3 ;
    ANTENNADIFFAREA 2.176 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0336 LAYER M4 ;
    ANTENNAGATEAREA 0.8304 LAYER M4 ; 
    ANTENNAMAXAREACAR 19.538 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.200745 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.90239 LAYER V4 ;
  END SRAM_in_A_addr[8]
  PIN SRAM_in_A_addr[7] 
    ANTENNAPARTIALMETALAREA 2.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.9655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.454598 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER V3 ;
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0328 LAYER M4 ;
    ANTENNAGATEAREA 1.4328 LAYER M4 ; 
    ANTENNAMAXAREACAR 46.1989 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.47749 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.03577 LAYER V4 ;
  END SRAM_in_A_addr[7]
  PIN SRAM_in_A_addr[6] 
    ANTENNAPARTIALMETALAREA 12.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.127 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.524 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.6279 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.176251 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.11506 LAYER V3 ;
    ANTENNADIFFAREA 7.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER M4 ;
    ANTENNAGATEAREA 2.1576 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.3571 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.292788 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.88172 LAYER V4 ;
  END SRAM_in_A_addr[6]
  PIN SRAM_in_A_addr[5] 
    ANTENNADIFFAREA 3.996 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1896 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.6435 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.389662 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.843882 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0104 LAYER M4 ;
    ANTENNAGATEAREA 1.824 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.1917 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.395364 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.843882 LAYER V4 ;
  END SRAM_in_A_addr[5]
  PIN SRAM_in_A_addr[4] 
    ANTENNADIFFAREA 3.348 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.075 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9504 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.4998 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.209343 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.26263 LAYER V3 ;
  END SRAM_in_A_addr[4]
  PIN SRAM_in_A_addr[3] 
    ANTENNADIFFAREA 7.362 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0846 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1736 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.4605 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.16886 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V3 ;
  END SRAM_in_A_addr[3]
  PIN SRAM_in_A_addr[2] 
    ANTENNADIFFAREA 13.772 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1238 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0848 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.1962 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.446572 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.33637 LAYER V3 ;
    ANTENNADIFFAREA 13.772 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAGATEAREA 1.5312 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.1628 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.456499 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.33637 LAYER V4 ;
  END SRAM_in_A_addr[2]
  PIN SRAM_in_A_addr[1] 
    ANTENNADIFFAREA 10.52 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3216 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.8477 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.374198 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.05521 LAYER V3 ;
    ANTENNADIFFAREA 10.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER M4 ;
    ANTENNAGATEAREA 1.9824 LAYER M4 ; 
    ANTENNAMAXAREACAR 40.4797 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.410921 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.05521 LAYER V4 ;
  END SRAM_in_A_addr[1]
  PIN SRAM_in_A_addr[0] 
    ANTENNADIFFAREA 13.772 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0758 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4248 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.3658 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.427468 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.869356 LAYER V3 ;
    ANTENNADIFFAREA 13.772 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER M4 ;
    ANTENNAGATEAREA 1.7952 LAYER M4 ; 
    ANTENNAMAXAREACAR 48.1145 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.4854 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.01228 LAYER V4 ;
  END SRAM_in_A_addr[0]
  PIN SRAM_in_B_addr[9] 
    ANTENNADIFFAREA 7.676 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 32.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.323 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8496 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.8993 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.515063 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.32558 LAYER V3 ;
  END SRAM_in_B_addr[9]
  PIN SRAM_in_B_addr[8] 
    ANTENNADIFFAREA 3.996 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 30.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3078 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3344 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.3755 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.323795 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.99794 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.68 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0472 LAYER M4 ;
    ANTENNAGATEAREA 1.6464 LAYER M4 ; 
    ANTENNAMAXAREACAR 35.218 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.352464 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.99794 LAYER V4 ;
  END SRAM_in_B_addr[8]
  PIN SRAM_in_B_addr[7] 
    ANTENNADIFFAREA 3.996 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 30.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.303 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.44 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.5384 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.370711 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.93798 LAYER V3 ;
  END SRAM_in_B_addr[7]
  PIN SRAM_in_B_addr[6] 
    ANTENNADIFFAREA 3.996 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 22.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2246 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5424 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.9567 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.523399 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.20234 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M4 ;
    ANTENNAGATEAREA 1.7304 LAYER M4 ; 
    ANTENNAMAXAREACAR 52.6271 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.530334 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.23013 LAYER V4 ;
  END SRAM_in_B_addr[6]
  PIN SRAM_in_B_addr[5] 
    ANTENNAPARTIALMETALAREA 14.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1462 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3784 LAYER M4 ; 
    ANTENNAMAXAREACAR 16.8437 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.174892 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.19053 LAYER V4 ;
  END SRAM_in_B_addr[5]
  PIN SRAM_in_B_addr[4] 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0198 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0904 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8144 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.1358 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.2839 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.65699 LAYER V4 ;
  END SRAM_in_B_addr[4]
  PIN SRAM_in_B_addr[3] 
    ANTENNAPARTIALMETALAREA 8.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0854 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 12.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1264 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2168 LAYER M4 ; 
    ANTENNAMAXAREACAR 71.952 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.72933 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.08495 LAYER V4 ;
  END SRAM_in_B_addr[3]
  PIN SRAM_in_B_addr[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 18.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.184 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5912 LAYER M4 ; 
    ANTENNAMAXAREACAR 42.4232 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.438004 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.61169 LAYER V4 ;
  END SRAM_in_B_addr[2]
  PIN SRAM_in_B_addr[1] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1544 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3464 LAYER M4 ; 
    ANTENNAMAXAREACAR 34.4434 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.345471 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.67232 LAYER V4 ;
  END SRAM_in_B_addr[1]
  PIN SRAM_in_B_addr[0] 
    ANTENNAPARTIALMETALAREA 12.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1262 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.762 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0824 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0176 LAYER M4 ; 
    ANTENNAMAXAREACAR 44.3633 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.447259 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38339 LAYER V4 ;
  END SRAM_in_B_addr[0]
  PIN SRAM_WENB12 
    ANTENNAPARTIALMETALAREA 13.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1374 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 12.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1592 LAYER M4 ; 
    ANTENNAMAXAREACAR 53.1084 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.536859 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.4311 LAYER V4 ;
  END SRAM_WENB12
  PIN SRAM_WENB34 
    ANTENNAPARTIALMETALAREA 13.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1366 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5288 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.7448 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.333261 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.00148 LAYER V4 ;
  END SRAM_WENB34
END CNN_controller

END LIBRARY
