VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PLL_integerN_top_lef
  CLASS BLOCK ;
  ORIGIN 6.07 0 ;
  FOREIGN PLL_integerN_top_lef -6.07 0 ;
  SIZE 57.31 BY 72.3 ;
  SYMMETRY X Y R90 ;
  PIN avdd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -4.72 0.73 -4.07 1.38 ;
    END
  END avdd
  PIN agnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 42.85 0 43.65 0.78 ;
    END
  END agnd
  PIN divide_num[0]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 24.95 0.16 25.15 0.36 ;
    END
  END divide_num[0]
  PIN divide_num[1]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 19.75 0.16 19.95 0.36 ;
    END
  END divide_num[1]
  PIN divide_num[2]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 14.55 0.17 14.75 0.37 ;
    END
  END divide_num[2]
  PIN fout
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.04 67.83 51.24 68.03 ;
    END
  END fout
  PIN Iref
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 50.6 58.2 50.8 58.4 ;
    END
  END Iref
  PIN Vctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 50.6 56.7 50.8 56.9 ;
    END
  END Vctrl
  PIN fref
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT -6.07 61.8 -5.87 62 ;
    END
  END fref
  OBS
    LAYER M1 ;
      RECT -2.73 71.36 50.28 72.3 ;
      RECT -4.72 3.3 -2.5 72.29 ;
      RECT 48.73 70.15 48.89 72.3 ;
      RECT 47.01 68.87 47.17 72.3 ;
      RECT 40.04 70.15 40.2 72.3 ;
      RECT 38.32 68.87 38.48 72.3 ;
      RECT 5.05 70.4 5.5 72.3 ;
      RECT 2.93 70.4 3.09 72.3 ;
      RECT 1.24 70.4 1.4 72.3 ;
      RECT -4.72 53.39 -1.3 72.29 ;
      RECT 49.32 65.92 49.52 70.44 ;
      RECT 49.32 67.77 49.64 68.09 ;
      RECT -0.35 0.73 0.45 2.58 ;
      RECT 44.05 0.73 44.85 2.36 ;
      RECT -2.15 0.73 44.85 1.38 ;
      RECT 3.57 69.03 3.73 70.8 ;
      RECT 3.36 69.03 3.73 70.78 ;
      RECT 0.3 69.78 0.76 70.82 ;
      RECT 0.3 66.27 0.46 70.82 ;
      RECT 0.28 64.19 50.29 65.06 ;
      RECT 4.31 70.09 4.47 70.8 ;
      RECT 1.88 69.91 2.04 70.8 ;
    LAYER M1 SPACING 0.16 ;
      RECT -6.07 1.7 51.24 72.3 ;
      RECT -3.75 0 51.24 72.3 ;
      RECT -6.07 0 -5.04 72.3 ;
      RECT -6.07 0 51.24 0.41 ;
    LAYER M2 ;
      RECT 42.85 2.7 43.65 35.9 ;
      RECT 41.15 2.62 42.15 4.6 ;
      RECT 24.95 2.28 25.15 5.4 ;
      RECT 19.75 2.28 19.95 5.4 ;
      RECT 14.55 2.29 14.75 9.8 ;
      RECT -4.72 53.39 -1.38 72.29 ;
    LAYER M2 SPACING 0.2 ;
      RECT -6.07 68.33 51.24 72.3 ;
      RECT -6.07 1.68 50.74 72.3 ;
      RECT 43.95 0 51.24 67.53 ;
      RECT -3.77 1.08 51.24 67.53 ;
      RECT -6.07 0 -5.02 72.3 ;
      RECT -3.77 0.67 42.55 72.3 ;
      RECT 25.45 0 42.55 72.3 ;
      RECT 15.05 0.66 42.55 72.3 ;
      RECT -3.77 0 14.25 72.3 ;
      RECT 20.25 0 24.65 72.3 ;
      RECT 15.05 0 19.45 72.3 ;
      RECT -6.07 0 14.25 0.43 ;
    LAYER M3 ;
      RECT 41.75 6.8 41.95 7.4 ;
      RECT 41.35 6.8 41.95 7 ;
      RECT 41.35 30.8 41.55 31.8 ;
      RECT 40.95 31.2 41.55 31.4 ;
      RECT 2.95 6.8 39.55 7 ;
      RECT 2.95 6.4 3.15 7 ;
      RECT 38.55 7.2 38.75 7.8 ;
      RECT 38.15 7.2 38.75 7.4 ;
      RECT 22.55 14.4 22.75 15 ;
      RECT 21.75 14.4 21.95 15 ;
      RECT 21.75 14.4 38.35 14.6 ;
      RECT 38.15 14 38.35 14.6 ;
      RECT 26.55 16.8 26.75 17.4 ;
      RECT 32.15 16.8 38.35 17 ;
      RECT 26.55 16.8 27.95 17 ;
      RECT 27.75 16.4 27.95 17 ;
      RECT 32.15 16.4 32.35 17 ;
      RECT 27.75 16.4 32.35 16.6 ;
      RECT 32.15 17.6 32.35 18.2 ;
      RECT 32.15 17.6 37.15 17.8 ;
      RECT 12.15 7.2 12.35 7.8 ;
      RECT 12.15 7.2 35.95 7.4 ;
      RECT 26.95 19.2 35.95 19.4 ;
      RECT 35.75 18.8 35.95 19.4 ;
      RECT 26.95 18.8 27.15 19.4 ;
      RECT 20.95 21.6 34.75 21.8 ;
      RECT 20.95 21.2 21.15 21.8 ;
      RECT 16.95 21.2 21.15 21.4 ;
      RECT 16.95 20.8 17.15 21.4 ;
      RECT 29.35 18.4 34.35 18.6 ;
      RECT 34.15 18 34.35 18.6 ;
      RECT 29.35 18 29.55 18.6 ;
      RECT 22.15 18 29.55 18.2 ;
      RECT 28.15 17.6 28.35 18.2 ;
      RECT 22.15 17.6 22.35 18.2 ;
      RECT 28.15 12.8 30.35 13 ;
      RECT 30.15 12.4 30.35 13 ;
      RECT 29.75 17.2 29.95 17.8 ;
      RECT 29.55 17.2 30.15 17.4 ;
      RECT 28.95 7.6 29.15 8.2 ;
      RECT 24.95 7.6 25.15 8.2 ;
      RECT 24.95 7.6 29.15 7.8 ;
      RECT 20.15 8.4 20.35 9 ;
      RECT 20.15 8.4 25.95 8.6 ;
      RECT 25.75 8 25.95 8.6 ;
      RECT 20.15 22.8 23.55 23 ;
      RECT 23.35 22.4 23.55 23 ;
      RECT 20.15 22.4 20.35 23 ;
      RECT 23.35 22.4 24.75 22.6 ;
      RECT 24.55 22 24.75 22.6 ;
      RECT 12.55 22.4 20.35 22.6 ;
      RECT 12.55 22 12.75 22.6 ;
      RECT 23.75 15.6 23.95 16.2 ;
      RECT 22.15 15.6 23.95 15.8 ;
      RECT 22.15 15.2 22.35 15.8 ;
      RECT 20.15 19.6 20.35 20.2 ;
      RECT 20.15 19.6 23.55 19.8 ;
      RECT 22.55 7.6 22.75 8.2 ;
      RECT 22.15 7.6 22.75 7.8 ;
      RECT 15.35 5.2 21.95 5.4 ;
      RECT 21.75 4.8 21.95 5.4 ;
      RECT 19.75 4.8 19.95 5.4 ;
      RECT 15.35 4.8 15.55 5.4 ;
      RECT 18.15 15.2 20.75 15.4 ;
      RECT 20.55 14.8 20.75 15.4 ;
      RECT 13.35 16.8 13.55 17.4 ;
      RECT 12.95 16.8 13.55 17 ;
      RECT 10.55 12.8 10.75 13.4 ;
      RECT 10.55 12.8 13.15 13 ;
      RECT 2.95 21.6 4.75 21.8 ;
      RECT 2.95 21.2 3.15 21.8 ;
      RECT -1.55 21.2 3.15 21.4 ;
      RECT 3.35 21.2 3.95 21.4 ;
      RECT 3.75 20.8 3.95 21.4 ;
      RECT 3.35 7.2 3.55 7.8 ;
      RECT 2.95 7.2 3.55 7.4 ;
      RECT 2.15 13.2 3.15 13.4 ;
      RECT 2.95 12.8 3.15 13.4 ;
      RECT 2.55 7.2 2.75 7.8 ;
      RECT 2.15 7.2 2.75 7.4 ;
      RECT 35.01 56.7 50.3 56.9 ;
      RECT 29.94 58.2 50.3 58.4 ;
      RECT 41.75 22 46.45 22.2 ;
      RECT 41.55 2.62 44.53 3.62 ;
      RECT 42.05 5.42 44.53 5.82 ;
      RECT 42.85 6.22 44.53 7.22 ;
      RECT 42.85 7.62 44.53 8.62 ;
      RECT 42.85 9.02 44.53 10.02 ;
      RECT 42.85 10.42 44.53 11.42 ;
      RECT 42.85 11.82 44.53 12.82 ;
      RECT 42.85 13.22 44.53 14.22 ;
      RECT 42.85 14.62 44.53 15.62 ;
      RECT 42.85 16.02 44.53 17.02 ;
      RECT 42.85 17.42 44.53 18.42 ;
      RECT 42.85 18.82 44.53 19.82 ;
      RECT 41.25 24.5 44.53 25.5 ;
      RECT 41.25 25.9 44.53 26.9 ;
      RECT 41.25 27.3 44.53 28.3 ;
      RECT 41.25 28.7 44.53 29.7 ;
      RECT 43.25 31.5 44.53 32.5 ;
      RECT 43.25 32.9 44.53 33.9 ;
      RECT 43.25 34.3 44.53 35.3 ;
      RECT 43.25 35.7 44.53 36.7 ;
      RECT 40.15 4.02 44.15 5.02 ;
      RECT 39.85 34.5 42.85 35.5 ;
      RECT 41.65 35.9 42.85 36.7 ;
      RECT 41.25 8.3 42.45 9.3 ;
      RECT 41.25 9.7 42.45 10.7 ;
      RECT 41.25 11.1 42.45 12.1 ;
      RECT 41.25 12.5 42.45 13.5 ;
      RECT 41.25 13.9 42.45 14.9 ;
      RECT 41.25 15.3 42.45 16.3 ;
      RECT 41.25 16.7 42.45 17.7 ;
      RECT 41.25 18.1 42.45 19.1 ;
      RECT 3.35 32 42.35 32.2 ;
      RECT 27.35 43.02 42.31 43.22 ;
      RECT 27.35 47.02 42.31 47.22 ;
      RECT 2.55 20.4 41.55 20.6 ;
      RECT 37.25 35.9 41.25 36.7 ;
      RECT 37.15 2.62 41.15 3.62 ;
      RECT 3.75 6 41.15 6.2 ;
      RECT 37.91 54.33 41.1 54.53 ;
      RECT 39.65 7.9 40.85 8.9 ;
      RECT 39.65 9.3 40.85 10.3 ;
      RECT 39.65 10.7 40.85 11.7 ;
      RECT 39.65 12.1 40.85 13.1 ;
      RECT 39.65 13.5 40.85 14.5 ;
      RECT 39.65 14.9 40.85 15.9 ;
      RECT 39.65 16.3 40.85 17.3 ;
      RECT 39.65 17.7 40.85 18.7 ;
      RECT 39.85 22.9 40.85 23.9 ;
      RECT 39.85 24.3 40.85 25.3 ;
      RECT 39.85 25.7 40.85 26.7 ;
      RECT 36.71 53.93 40.11 54.13 ;
      RECT 35.75 4.02 39.75 5.02 ;
      RECT 36.54 51.41 39.54 51.61 ;
      RECT 35.65 22.9 39.45 23.9 ;
      RECT 35.65 24.3 39.45 25.3 ;
      RECT 35.45 34.5 39.45 35.5 ;
      RECT 38.05 10.1 39.25 11.1 ;
      RECT 38.05 11.5 39.25 12.5 ;
      RECT 38.05 12.9 39.25 13.3 ;
      RECT 36.35 15.2 39.25 15.8 ;
      RECT 37.75 17.6 39.25 18.6 ;
      RECT 2.55 28.4 39.15 28.6 ;
      RECT 30.95 31.2 38.75 31.4 ;
      RECT 23.35 27.6 38.35 27.8 ;
      RECT 35.25 9.5 37.65 10.5 ;
      RECT 35.35 12.1 37.55 13.1 ;
      RECT 33.45 10.9 37.45 11.7 ;
      RECT 6.73 67.84 36.93 68.04 ;
      RECT 32.85 35.9 36.85 36.7 ;
      RECT 32.75 2.62 36.75 3.62 ;
      RECT 31.95 15.2 35.95 15.8 ;
      RECT 31.35 4.02 35.35 5.02 ;
      RECT 29.91 51.41 35.34 51.61 ;
      RECT 0.7 64.62 35.31 64.82 ;
      RECT 34.15 22.7 35.25 23.7 ;
      RECT 32.35 24.1 35.25 25.1 ;
      RECT 31.05 34.5 35.05 35.5 ;
      RECT 30.95 12.1 34.95 13.1 ;
      RECT 30.85 9.5 34.85 10.5 ;
      RECT 31.11 54.33 34.51 54.53 ;
      RECT 29.75 22.7 33.75 23.7 ;
      RECT 29.91 53.93 33.31 54.13 ;
      RECT 30.85 10.9 33.05 11.7 ;
      RECT 28.45 35.9 32.45 36.7 ;
      RECT 28.35 2.62 32.35 3.62 ;
      RECT 27.95 24.1 31.95 25.1 ;
      RECT 27.55 15.2 31.55 15.8 ;
      RECT 26.95 4.02 30.95 5.02 ;
      RECT 26.65 34.5 30.65 35.5 ;
      RECT 28.95 11.1 30.45 11.7 ;
      RECT 13.35 31.6 30.35 31.8 ;
      RECT 26.15 10 29.95 10.2 ;
      RECT 25.35 22.7 29.35 23.7 ;
      RECT 24.55 11.1 28.55 11.7 ;
      RECT 24.05 35.9 28.05 36.7 ;
      RECT 23.95 2.62 27.95 3.62 ;
      RECT 25.35 24.1 27.55 25.1 ;
      RECT 24.55 15.2 27.15 16.2 ;
      RECT 22.55 4.02 26.55 5.02 ;
      RECT 22.25 34.5 26.25 35.5 ;
      RECT 20.44 52.24 26.09 52.44 ;
      RECT 23.55 16.8 25.95 17.2 ;
      RECT 24.25 9.6 25.25 10.6 ;
      RECT 20.43 51.5 24.85 51.7 ;
      RECT 20.15 11.1 24.15 11.7 ;
      RECT 22.95 6.4 23.95 6.6 ;
      RECT 19.95 9.6 23.85 10.6 ;
      RECT 19.65 35.9 23.65 36.7 ;
      RECT 19.55 2.62 23.55 3.62 ;
      RECT 19.95 23.7 23.55 24.7 ;
      RECT 19.95 25.1 23.55 26.1 ;
      RECT 21.85 16.4 23.15 17 ;
      RECT 3.75 14 22.75 14.2 ;
      RECT 17.85 34.5 21.85 35.5 ;
      RECT 18.15 6.4 20.35 6.6 ;
      RECT 14.15 17.6 20.35 17.8 ;
      RECT 18.53 47.34 19.93 47.54 ;
      RECT 18.53 56.54 19.93 56.74 ;
      RECT 17.65 8.3 19.55 8.9 ;
      RECT 16.95 9.3 19.55 10.3 ;
      RECT 17.35 11.2 19.55 11.4 ;
      RECT 16.75 23.2 19.55 24.2 ;
      RECT 18.55 24.6 19.55 25.6 ;
      RECT 14.53 45.74 19.53 45.94 ;
      RECT 14.53 58.14 19.53 58.34 ;
      RECT 15.25 35.9 19.25 36.7 ;
      RECT 15.15 2.62 19.15 3.62 ;
      RECT 16.15 4.02 19.15 4.42 ;
      RECT 14.93 44.94 19.13 45.14 ;
      RECT 14.93 58.94 19.13 59.14 ;
      RECT 17.33 46.54 18.73 46.74 ;
      RECT 17.33 57.34 18.73 57.54 ;
      RECT -5.57 61.8 18.43 62 ;
      RECT -1.56 39.3 18.33 40.88 ;
      RECT 14.95 24.6 18.15 25.6 ;
      RECT 16.13 42.55 17.93 42.75 ;
      RECT -0.27 51.74 17.93 51.94 ;
      RECT 16.13 61.33 17.93 61.53 ;
      RECT 15.75 13.2 17.55 13.4 ;
      RECT 13.45 34.5 17.45 35.5 ;
      RECT 13.25 8.3 17.25 8.9 ;
      RECT 16.05 15.1 17.05 15.9 ;
      RECT 13.15 10.5 16.55 11.5 ;
      RECT 13.35 9.6 16.35 9.8 ;
      RECT 12.35 23.2 16.35 24.2 ;
      RECT 14.53 44.54 15.93 44.74 ;
      RECT 14.53 59.34 15.93 59.54 ;
      RECT 10.85 35.9 14.85 36.7 ;
      RECT 11.65 2.62 14.75 3.62 ;
      RECT 13.25 4.02 14.75 5.02 ;
      RECT 12.35 24.6 14.55 25.6 ;
      RECT 11.35 13.6 13.55 13.8 ;
      RECT 9.05 34.5 13.05 35.5 ;
      RECT 10.35 8.7 12.75 9.7 ;
      RECT 10.35 10.1 12.75 11.1 ;
      RECT 10.35 11.5 12.75 12.1 ;
      RECT 12.15 5.2 12.35 5.8 ;
      RECT 10.25 16.5 12.05 17.5 ;
      RECT 9.75 21.5 11.95 22.5 ;
      RECT 9.75 22.9 11.95 23.9 ;
      RECT 9.75 24.3 11.95 25.3 ;
      RECT 9.75 25.7 11.95 26.7 ;
      RECT 9.17 2.62 11.25 3.62 ;
      RECT 7.37 4.02 11.25 5.02 ;
      RECT 6.45 35.9 10.45 36.7 ;
      RECT 8.85 7.9 9.95 8.9 ;
      RECT 8.85 9.3 9.95 10.3 ;
      RECT 8.85 10.7 9.95 11.7 ;
      RECT 8.85 12.1 9.95 13.1 ;
      RECT 5.85 16.5 9.85 17.5 ;
      RECT 5.35 21.5 9.35 22.5 ;
      RECT 5.35 22.9 9.35 23.9 ;
      RECT 5.35 24.3 9.35 25.3 ;
      RECT 5.35 25.7 9.35 26.7 ;
      RECT 4.77 2.62 8.77 3.62 ;
      RECT 4.65 34.5 8.65 35.5 ;
      RECT 4.45 9.3 8.45 10.3 ;
      RECT 4.45 10.7 8.45 11.7 ;
      RECT 4.45 12.1 8.45 13.1 ;
      RECT 2.97 4.02 6.97 5.02 ;
      RECT 2.05 35.9 6.05 36.7 ;
      RECT 3.25 16.5 5.45 17.5 ;
      RECT 2.75 25.2 4.95 26.2 ;
      RECT 0.37 2.62 4.37 3.62 ;
      RECT 2.05 34.5 4.25 35.5 ;
      RECT 2.05 10.1 4.05 11.1 ;
      RECT 0.37 15.7 2.85 16.7 ;
      RECT 0.37 17.1 2.85 18.1 ;
      RECT 0.37 4.02 2.57 5.02 ;
      RECT 0.37 23.4 2.35 24.4 ;
      RECT 0.37 24.8 2.35 25.8 ;
      RECT 0.37 5.42 2.05 6.22 ;
      RECT 0.37 9.7 1.65 10.7 ;
      RECT 0.37 19.9 1.65 20.5 ;
      RECT 0.37 29 1.65 30 ;
      RECT 0.37 30.4 1.65 31.4 ;
      RECT 0.37 31.8 1.65 32.8 ;
      RECT 0.37 33.2 1.65 34.2 ;
      RECT 0.37 34.6 1.65 35.6 ;
      RECT 0.37 36 1.65 36.6 ;
    LAYER M4 ;
      RECT 41.75 22 42.35 22.2 ;
      RECT 41.75 6.8 41.95 22.2 ;
      RECT 41.35 20.4 41.55 31.4 ;
      RECT 40.95 20.4 41.55 20.6 ;
      RECT 38.15 31.2 38.75 31.4 ;
      RECT 38.55 7.2 38.75 31.4 ;
      RECT 29.75 21.6 30.35 21.8 ;
      RECT 29.75 7.2 29.95 21.8 ;
      RECT 29.35 10 29.95 10.2 ;
      RECT 29.75 7.2 30.35 7.4 ;
      RECT 23.35 27.6 23.95 27.8 ;
      RECT 23.35 6.4 23.55 27.8 ;
      RECT 23.35 6.4 23.95 6.6 ;
      RECT 22.15 14 22.75 14.2 ;
      RECT 22.55 7.6 22.75 14.2 ;
      RECT 19.75 17.6 20.35 17.8 ;
      RECT 20.15 6.4 20.35 17.8 ;
      RECT 19.75 6.4 20.35 6.6 ;
      RECT 16.95 13.2 17.55 13.4 ;
      RECT 17.35 7.2 17.55 13.4 ;
      RECT 17.35 7.2 17.95 7.4 ;
      RECT 13.35 31.6 13.95 31.8 ;
      RECT 13.35 16.8 13.55 31.8 ;
      RECT 3.75 6 3.95 21.4 ;
      RECT 3.75 6 4.35 6.2 ;
      RECT 3.35 32 3.95 32.2 ;
      RECT 3.35 7.2 3.55 32.2 ;
      RECT 2.55 28.4 3.15 28.6 ;
      RECT 2.55 7.2 2.75 28.6 ;
      RECT 43.85 25.7 44.45 29.7 ;
      RECT 43.85 30.1 44.45 32.7 ;
      RECT 43.77 2.62 44.37 4.3 ;
      RECT 43.37 33.1 44.37 36.78 ;
      RECT 42.37 2.62 43.37 4.3 ;
      RECT 41.97 33.1 42.97 36.78 ;
      RECT 40.97 2.62 41.97 4.3 ;
      RECT 40.57 33.1 41.57 36.78 ;
      RECT 40.45 6.7 40.85 10.7 ;
      RECT 40.45 11.1 40.85 15.1 ;
      RECT 39.57 2.62 40.57 4.3 ;
      RECT 39.17 33.1 40.17 36.78 ;
      RECT 38.17 2.62 39.17 4.3 ;
      RECT 37.77 33.1 38.77 36.78 ;
      RECT 36.77 2.62 37.77 4.3 ;
      RECT 36.37 33.1 37.37 36.78 ;
      RECT 35.45 6.7 36.45 7.9 ;
      RECT 35.45 21.1 36.45 22.3 ;
      RECT 35.45 28.7 36.45 30.7 ;
      RECT 35.37 2.62 36.37 4.3 ;
      RECT 35.05 8.3 36.05 10.5 ;
      RECT 35.05 10.9 36.05 14.9 ;
      RECT 35.05 15.3 36.05 19.3 ;
      RECT 35.05 19.7 36.05 20.7 ;
      RECT 34.97 33.1 35.97 36.78 ;
      RECT 34.45 22.7 35.45 26.7 ;
      RECT 34.45 27.1 35.45 28.3 ;
      RECT 34.45 31.1 35.45 32.7 ;
      RECT 34.05 6.7 35.05 7.9 ;
      RECT 34.05 21.1 35.05 22.3 ;
      RECT 34.05 28.7 35.05 30.7 ;
      RECT 33.97 2.62 34.97 4.3 ;
      RECT 33.65 8.3 34.65 12.3 ;
      RECT 33.65 12.7 34.65 16.7 ;
      RECT 33.65 17.1 34.65 20.7 ;
      RECT 33.57 33.1 34.57 36.78 ;
      RECT 33.05 22.7 34.05 26.7 ;
      RECT 33.05 27.1 34.05 28.3 ;
      RECT 33.05 31.1 34.05 32.7 ;
      RECT 32.65 6.7 33.65 7.9 ;
      RECT 32.65 21.1 33.65 22.3 ;
      RECT 32.65 28.7 33.65 30.7 ;
      RECT 32.57 2.62 33.57 4.3 ;
      RECT 32.25 8.3 33.25 10.5 ;
      RECT 32.25 10.9 33.25 14.9 ;
      RECT 32.25 15.3 33.25 19.3 ;
      RECT 32.25 19.7 33.25 20.7 ;
      RECT 32.17 33.1 33.17 36.78 ;
      RECT 31.65 22.7 32.65 26.7 ;
      RECT 31.65 27.1 32.65 28.3 ;
      RECT 31.65 31.1 32.65 32.7 ;
      RECT 31.25 28.7 32.25 30.7 ;
      RECT 31.17 2.62 32.17 4.3 ;
      RECT 30.85 8.3 31.85 12.3 ;
      RECT 30.85 12.7 31.85 16.7 ;
      RECT 30.85 17.1 31.85 20.7 ;
      RECT 30.77 33.1 31.77 36.78 ;
      RECT 30.25 22.7 31.25 26.7 ;
      RECT 30.25 27.1 31.25 28.3 ;
      RECT 30.25 31.1 31.25 32.7 ;
      RECT 29.85 28.7 30.85 30.7 ;
      RECT 29.77 2.62 30.77 4.3 ;
      RECT 29.37 33.1 30.37 36.78 ;
      RECT 28.85 22.7 29.85 26.7 ;
      RECT 28.85 27.1 29.85 28.3 ;
      RECT 28.85 31.1 29.85 32.7 ;
      RECT 28.45 28.7 29.45 30.7 ;
      RECT 28.37 2.62 29.37 4.3 ;
      RECT 27.97 33.1 28.97 36.78 ;
      RECT 27.45 31.1 28.45 32.7 ;
      RECT 27.05 28.7 28.05 30.7 ;
      RECT 26.97 2.62 27.97 4.3 ;
      RECT 26.57 33.1 27.57 36.78 ;
      RECT 26.25 4.7 27.25 6.9 ;
      RECT 26.25 7.3 27.25 11.3 ;
      RECT 26.25 11.7 27.25 15.7 ;
      RECT 26.25 16.1 27.25 20.1 ;
      RECT 26.25 20.5 27.25 24.5 ;
      RECT 26.25 24.9 27.25 28.3 ;
      RECT 26.05 31.1 27.05 32.7 ;
      RECT 25.57 2.62 26.57 4.3 ;
      RECT 25.17 33.1 26.17 36.78 ;
      RECT 24.65 31.1 25.65 32.7 ;
      RECT 24.17 2.62 25.17 4.3 ;
      RECT 23.77 33.1 24.77 36.78 ;
      RECT 23.25 31.1 24.25 32.7 ;
      RECT 22.77 2.62 23.77 4.3 ;
      RECT 22.37 33.1 23.37 36.78 ;
      RECT 21.85 31.1 22.85 32.7 ;
      RECT 21.37 2.62 22.37 4.3 ;
      RECT 20.97 33.1 21.97 36.78 ;
      RECT 20.45 31.1 21.45 32.7 ;
      RECT 20.05 21.3 21.05 25.3 ;
      RECT 20.05 25.7 21.05 29.3 ;
      RECT 20.05 29.7 21.05 30.7 ;
      RECT 19.97 2.62 20.97 4.3 ;
      RECT 19.57 33.1 20.57 36.78 ;
      RECT 19.05 31.1 20.05 32.7 ;
      RECT 18.65 23.1 19.65 27.1 ;
      RECT 18.65 27.5 19.65 30.7 ;
      RECT 18.57 2.62 19.57 4.3 ;
      RECT 18.17 33.1 19.17 36.78 ;
      RECT 17.65 31.1 18.65 32.7 ;
      RECT 17.25 20.7 18.25 24.7 ;
      RECT 17.25 25.1 18.25 29.1 ;
      RECT 17.25 29.5 18.25 30.7 ;
      RECT 17.17 2.62 18.17 4.3 ;
      RECT 16.77 33.1 17.77 36.78 ;
      RECT 16.25 31.1 17.25 32.7 ;
      RECT 15.85 18.9 16.85 22.9 ;
      RECT 15.85 23.3 16.85 27.3 ;
      RECT 15.77 2.62 16.77 4.3 ;
      RECT 15.37 33.1 16.37 36.78 ;
      RECT 14.65 4.7 15.65 8.3 ;
      RECT 13.97 33.1 14.97 36.78 ;
      RECT 13.05 11.3 14.05 14.5 ;
      RECT 12.57 33.1 13.57 36.78 ;
      RECT 12.15 5.2 12.35 7.8 ;
      RECT 11.17 33.1 12.17 36.78 ;
      RECT 10.45 11.5 11.25 15.5 ;
      RECT 10.45 15.9 11.25 19.9 ;
      RECT 10.45 20.3 11.25 21.9 ;
      RECT 10.05 22.3 11.05 26.3 ;
      RECT 10.05 26.7 11.05 30.7 ;
      RECT 10.05 31.5 11.05 32.7 ;
      RECT 9.77 33.1 10.77 36.78 ;
      RECT 9.05 7.1 10.05 9.3 ;
      RECT 9.05 9.7 10.05 13.7 ;
      RECT 9.05 14.1 10.05 18.1 ;
      RECT 9.05 18.5 10.05 21.9 ;
      RECT 8.77 2.62 9.77 5.1 ;
      RECT 8.65 22.3 9.65 24.5 ;
      RECT 8.65 24.9 9.65 28.9 ;
      RECT 8.65 29.3 9.65 31.1 ;
      RECT 8.65 31.5 9.65 32.7 ;
      RECT 8.37 33.1 9.37 36.78 ;
      RECT 8.05 5.5 9.05 6.7 ;
      RECT 7.65 7.1 8.65 11.1 ;
      RECT 7.65 11.5 8.65 15.5 ;
      RECT 7.65 15.9 8.65 19.9 ;
      RECT 7.65 20.3 8.65 21.9 ;
      RECT 7.37 2.62 8.37 5.1 ;
      RECT 7.25 22.3 8.25 26.3 ;
      RECT 7.25 26.7 8.25 30.7 ;
      RECT 7.25 31.5 8.25 32.7 ;
      RECT 6.97 33.1 7.97 36.78 ;
      RECT 6.65 5.5 7.65 6.7 ;
      RECT 6.25 7.1 7.25 9.3 ;
      RECT 6.25 9.7 7.25 13.7 ;
      RECT 6.25 14.1 7.25 18.1 ;
      RECT 6.25 18.5 7.25 21.9 ;
      RECT 5.97 2.62 6.97 5.1 ;
      RECT 5.85 22.3 6.85 24.5 ;
      RECT 5.85 24.9 6.85 28.9 ;
      RECT 5.85 29.3 6.85 31.1 ;
      RECT 4.57 2.62 5.57 5.1 ;
      RECT 3.17 2.62 4.17 5.1 ;
      RECT 2.95 6.4 3.15 13.4 ;
      RECT 1.77 33.9 2.37 36.78 ;
      RECT 0.37 2.62 1.37 5.5 ;
      RECT 0.37 32.3 1.37 35.38 ;
      RECT 0.37 35.78 1.37 36.78 ;
    LAYER M5 ;
      RECT 43.53 2.62 44.53 3.62 ;
      RECT 42.57 4.02 44.53 5.02 ;
      RECT 42.57 6.82 44.53 7.82 ;
      RECT 42.57 9.62 44.53 10.62 ;
      RECT 42.57 12.42 44.53 13.42 ;
      RECT 42.57 15.22 44.53 16.22 ;
      RECT 42.57 18.02 44.53 19.02 ;
      RECT 42.57 20.82 44.53 21.82 ;
      RECT 42.57 23.62 44.53 24.62 ;
      RECT 42.57 26.42 44.53 27.42 ;
      RECT 42.57 29.22 44.53 30.22 ;
      RECT 43.53 33.42 44.53 34.42 ;
      RECT 43.53 36.22 44.53 36.62 ;
      RECT 39.97 2.62 43.13 3.62 ;
      RECT 39.97 33.42 43.13 34.42 ;
      RECT 39.97 36.22 43.13 36.62 ;
      RECT 38.17 4.02 42.17 5.02 ;
      RECT 38.17 6.82 42.17 7.82 ;
      RECT 38.17 9.62 42.17 10.62 ;
      RECT 38.17 12.42 42.17 13.42 ;
      RECT 38.17 15.22 42.17 16.22 ;
      RECT 38.17 18.02 42.17 19.02 ;
      RECT 38.17 20.82 42.17 21.82 ;
      RECT 38.17 23.62 42.17 24.62 ;
      RECT 38.17 26.42 42.17 27.42 ;
      RECT 38.17 29.22 42.17 30.22 ;
      RECT 35.57 2.62 39.57 3.62 ;
      RECT 35.57 33.42 39.57 34.42 ;
      RECT 35.57 36.22 39.57 36.62 ;
      RECT 33.77 4.02 37.77 5.02 ;
      RECT 33.77 6.82 37.77 7.82 ;
      RECT 33.77 9.62 37.77 10.62 ;
      RECT 33.77 12.42 37.77 13.42 ;
      RECT 33.77 15.22 37.77 16.22 ;
      RECT 33.77 18.02 37.77 19.02 ;
      RECT 33.77 20.82 37.77 21.82 ;
      RECT 33.77 23.62 37.77 24.62 ;
      RECT 33.77 26.42 37.77 27.42 ;
      RECT 33.77 29.22 37.77 30.22 ;
      RECT 31.17 2.62 35.17 3.62 ;
      RECT 31.17 33.42 35.17 34.42 ;
      RECT 31.17 36.22 35.17 36.62 ;
      RECT 29.37 6.82 33.37 7.82 ;
      RECT 29.37 9.62 33.37 10.62 ;
      RECT 29.37 12.42 33.37 13.42 ;
      RECT 29.37 15.22 33.37 16.22 ;
      RECT 29.37 18.02 33.37 19.02 ;
      RECT 29.37 20.82 33.37 21.82 ;
      RECT 29.37 23.62 33.37 24.62 ;
      RECT 29.37 26.42 33.37 27.42 ;
      RECT 29.37 29.22 33.37 30.22 ;
      RECT 26.77 2.62 30.77 3.62 ;
      RECT 26.77 33.42 30.77 34.42 ;
      RECT 26.77 36.22 30.77 36.62 ;
      RECT 24.97 6.82 28.97 7.82 ;
      RECT 24.97 9.62 28.97 10.62 ;
      RECT 24.97 12.42 28.97 13.42 ;
      RECT 24.97 15.22 28.97 16.22 ;
      RECT 24.97 18.02 28.97 19.02 ;
      RECT 24.97 20.82 28.97 21.82 ;
      RECT 24.97 23.62 28.97 24.62 ;
      RECT 24.97 26.42 28.97 27.42 ;
      RECT 24.97 29.22 28.97 30.22 ;
      RECT 22.37 2.62 26.37 3.62 ;
      RECT 22.37 33.42 26.37 34.42 ;
      RECT 22.37 36.22 26.37 36.62 ;
      RECT 20.57 6.82 24.57 7.82 ;
      RECT 20.57 9.62 24.57 10.62 ;
      RECT 20.57 12.42 24.57 13.42 ;
      RECT 20.57 15.22 24.57 16.22 ;
      RECT 20.57 18.02 24.57 19.02 ;
      RECT 20.57 20.82 24.57 21.82 ;
      RECT 20.57 23.62 24.57 24.62 ;
      RECT 20.57 26.42 24.57 27.42 ;
      RECT 20.57 29.22 24.57 30.22 ;
      RECT 17.97 2.62 21.97 3.62 ;
      RECT 17.97 33.42 21.97 34.42 ;
      RECT 17.97 36.22 21.97 36.62 ;
      RECT 16.17 6.82 20.17 7.82 ;
      RECT 16.17 9.62 20.17 10.62 ;
      RECT 16.17 12.42 20.17 13.42 ;
      RECT 16.17 15.22 20.17 16.22 ;
      RECT 16.17 18.02 20.17 19.02 ;
      RECT 16.17 20.82 20.17 21.82 ;
      RECT 16.17 23.62 20.17 24.62 ;
      RECT 16.17 26.42 20.17 27.42 ;
      RECT 16.17 29.22 20.17 30.22 ;
      RECT 13.57 2.62 17.57 3.62 ;
      RECT 13.57 33.42 17.57 34.42 ;
      RECT 13.57 36.22 17.57 36.62 ;
      RECT 11.77 6.82 15.77 7.82 ;
      RECT 11.77 9.62 15.77 10.62 ;
      RECT 11.77 12.42 15.77 13.42 ;
      RECT 11.77 15.22 15.77 16.22 ;
      RECT 11.77 18.02 15.77 19.02 ;
      RECT 11.77 20.82 15.77 21.82 ;
      RECT 11.77 23.62 15.77 24.62 ;
      RECT 11.77 26.42 15.77 27.42 ;
      RECT 11.77 29.22 15.77 30.22 ;
      RECT 9.17 2.62 13.17 3.62 ;
      RECT 9.17 33.42 13.17 34.42 ;
      RECT 9.17 36.22 13.17 36.62 ;
      RECT 7.37 6.82 11.37 7.82 ;
      RECT 7.37 9.62 11.37 10.62 ;
      RECT 7.37 12.42 11.37 13.42 ;
      RECT 7.37 15.22 11.37 16.22 ;
      RECT 7.37 18.02 11.37 19.02 ;
      RECT 7.37 20.82 11.37 21.82 ;
      RECT 7.37 23.62 11.37 24.62 ;
      RECT 7.37 26.42 11.37 27.42 ;
      RECT 7.37 29.22 11.37 30.22 ;
      RECT 4.77 2.62 8.77 3.62 ;
      RECT 4.77 33.42 8.77 34.42 ;
      RECT 4.77 36.22 8.77 36.62 ;
      RECT 2.97 6.82 6.97 7.82 ;
      RECT 2.97 9.62 6.97 10.62 ;
      RECT 2.97 12.42 6.97 13.42 ;
      RECT 2.97 15.22 6.97 16.22 ;
      RECT 2.97 18.02 6.97 19.02 ;
      RECT 2.97 20.82 6.97 21.82 ;
      RECT 2.97 23.62 6.97 24.62 ;
      RECT 2.97 26.42 6.97 27.42 ;
      RECT 2.97 29.22 6.97 30.22 ;
      RECT 0.37 2.62 4.37 3.62 ;
      RECT 0.37 33.42 4.37 34.42 ;
      RECT 0.37 36.22 4.37 36.62 ;
      RECT 0.37 6.82 2.57 7.82 ;
      RECT 0.37 9.62 2.57 10.62 ;
      RECT 0.37 12.42 2.57 13.42 ;
      RECT 0.37 15.22 2.57 16.22 ;
      RECT 0.37 18.02 2.57 19.02 ;
      RECT 0.37 20.82 2.57 21.82 ;
      RECT 0.37 23.62 2.57 24.62 ;
      RECT 0.37 26.42 2.57 27.42 ;
      RECT 0.37 29.22 2.57 30.22 ;
  END
END PLL_integerN_top_lef

END LIBRARY
