

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO PE_top 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0142 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8352 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.64655 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0272749 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.191571 LAYER V3 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 4.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0454 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9552 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.4025 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.569324 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER V3 ;
  END reset
  PIN pe_in_pk_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0598 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.8462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.358333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER V3 ;
  END pe_in_pk_PE_state__2_
  PIN pe_in_pk_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.0513 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.883974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__1_
  PIN pe_in_pk_PE_state__0_ 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 106.282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.07628 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__0_
  PIN pe_in_pk_A__3__7_ 
    ANTENNAPARTIALMETALAREA 8.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0854 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 169.423 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.70128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__7_
  PIN pe_in_pk_A__3__6_ 
    ANTENNAPARTIALMETALAREA 7.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0758 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 127.115 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.27821 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__6_
  PIN pe_in_pk_A__3__5_ 
    ANTENNAPARTIALMETALAREA 6.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0654 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 121.987 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.22692 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__5_
  PIN pe_in_pk_A__3__4_ 
    ANTENNAPARTIALMETALAREA 6.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0614 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 113.013 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.13718 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__4_
  PIN pe_in_pk_A__3__3_ 
    ANTENNAPARTIALMETALAREA 6.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0614 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 106.603 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.07308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__3_
  PIN pe_in_pk_A__3__2_ 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0622 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 107.885 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.0859 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__2_
  PIN pe_in_pk_A__3__1_ 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0638 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 109.167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.09872 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__1_
  PIN pe_in_pk_A__3__0_ 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0638 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 106.603 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.07308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__0_
  PIN pe_in_pk_A__2__7_ 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0646 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.295 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.15 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__7_
  PIN pe_in_pk_A__2__6_ 
    ANTENNAPARTIALMETALAREA 6.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0662 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.577 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.16282 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__6_
  PIN pe_in_pk_A__2__5_ 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0646 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 113.013 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.13718 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__5_
  PIN pe_in_pk_A__2__4_ 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0646 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 107.885 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.0859 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__4_
  PIN pe_in_pk_A__2__3_ 
    ANTENNAPARTIALMETALAREA 6.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0654 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 110.449 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.11154 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__3_
  PIN pe_in_pk_A__2__2_ 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 91.2179 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.919231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__2_
  PIN pe_in_pk_A__2__1_ 
    ANTENNAPARTIALMETALAREA 4.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0406 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 74.5513 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.752564 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__1_
  PIN pe_in_pk_A__2__0_ 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0334 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.859 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.675641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__0_
  PIN pe_in_pk_A__1__7_ 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.9103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.496154 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__7_
  PIN pe_in_pk_A__1__6_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9615 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__6_
  PIN pe_in_pk_A__1__5_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.355128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__5_
  PIN pe_in_pk_A__1__4_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.5256 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.342308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__4_
  PIN pe_in_pk_A__1__3_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9615 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__3_
  PIN pe_in_pk_A__1__2_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.0641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.457692 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__2_
  PIN pe_in_pk_A__1__1_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.40641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__1_
  PIN pe_in_pk_A__1__0_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.508974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__0_
  PIN pe_in_pk_A__0__7_ 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0334 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.4487 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.611538 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__7_
  PIN pe_in_pk_A__0__6_ 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0334 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.859 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.675641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__6_
  PIN pe_in_pk_A__0__5_ 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.688462 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__5_
  PIN pe_in_pk_A__0__4_ 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.039 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 70.7051 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.714103 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__4_
  PIN pe_in_pk_A__0__3_ 
    ANTENNAPARTIALMETALAREA 4.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.043 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 74.5513 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.752564 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__3_
  PIN pe_in_pk_A__0__2_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 59.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.598718 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__2_
  PIN pe_in_pk_A__0__1_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 55.641 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.576282 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__0__1_
  PIN pe_in_pk_A__0__0_ 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0478 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 133.526 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.34231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__0_
  PIN pe_in_pk_wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 11.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.076 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 19.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1928 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 111.191 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.136 LAYER M4 ;
    ANTENNAMAXCUTCAR 5.76923 LAYER V4 ;
  END pe_in_pk_wrb_data__7_
  PIN pe_in_pk_wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 8.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0886 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 78.3648 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.789937 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.88679 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 24.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2448 LAYER M4 ;
    ANTENNAGATEAREA 0.444 LAYER M4 ; 
    ANTENNAMAXAREACAR 133.41 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.34129 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_wrb_data__6_
  PIN pe_in_pk_wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 8.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0854 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 151.795 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.53782 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 4.48718 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2608 LAYER M4 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 220.36 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 2.22558 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.48718 LAYER V4 ;
  END pe_in_pk_wrb_data__5_
  PIN pe_in_pk_wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 17.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1718 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 53.8365 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.544654 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.88679 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 16.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1632 LAYER M4 ;
    ANTENNAGATEAREA 0.444 LAYER M4 ; 
    ANTENNAMAXAREACAR 90.4131 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.912222 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.48718 LAYER V4 ;
  END pe_in_pk_wrb_data__4_
  PIN pe_in_pk_wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 16.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1678 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 78.0769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.794231 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 18.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1816 LAYER M4 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 125.862 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.27313 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_wrb_data__3_
  PIN pe_in_pk_wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0312 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 22.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.228 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 129.98 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.31857 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.48718 LAYER V4 ;
  END pe_in_pk_wrb_data__2_
  PIN pe_in_pk_wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 28.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2856 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 102.055 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.02738 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.48718 LAYER V4 ;
  END pe_in_pk_wrb_data__1_
  PIN pe_in_pk_wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 6.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.067 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 26.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2632 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 LAYER M4 ; 
    ANTENNAMAXAREACAR 111.483 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.12935 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_wrb_data__0_
  PIN pe_in_pk_wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.047 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.264 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.50152 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0554545 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.909091 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 27.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2736 LAYER M4 ;
    ANTENNAGATEAREA 1.056 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.6758 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.417576 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.909091 LAYER V4 ;
  END pe_in_pk_wrb_addr__3_
  PIN pe_in_pk_wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0478 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.044 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8136 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.1259 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.142056 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.38038 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 25.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26 LAYER M4 ;
    ANTENNAGATEAREA 1.7808 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.6812 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.288058 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END pe_in_pk_wrb_addr__2_
  PIN pe_in_pk_wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 4.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0478 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M2 ; 
    ANTENNAMAXAREACAR 30.2736 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.306219 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.746269 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M3 ;
    ANTENNAGATEAREA 0.3384 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.5195 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.32986 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.746269 LAYER V3 ;
  END pe_in_pk_wrb_addr__1_
  PIN pe_in_pk_wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 4.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0414 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1776 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.0011 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.113739 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M4 ;
    ANTENNAGATEAREA 0.7512 LAYER M4 ; 
    ANTENNAMAXAREACAR 14.2696 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.148447 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER V4 ;
  END pe_in_pk_wrb_addr__0_
  PIN pe_in_pk_wrb__3_ 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.039 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4608 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.5236 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.141073 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V3 ;
  END pe_in_pk_wrb__3_
  PIN pe_in_pk_wrb__2_ 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 14.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.148 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4608 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.6838 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.3904 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.980063 LAYER V4 ;
  END pe_in_pk_wrb__2_
  PIN pe_in_pk_wrb__1_ 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.027 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0872 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 30.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3048 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4608 LAYER M4 ; 
    ANTENNAMAXAREACAR 71.7149 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.724362 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.34409 LAYER V4 ;
  END pe_in_pk_wrb__1_
  PIN pe_in_pk_wrb__0_ 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1856 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 34.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.344 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4608 LAYER M4 ; 
    ANTENNAMAXAREACAR 82.1232 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.826624 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.980063 LAYER V4 ;
  END pe_in_pk_wrb__0_
  PIN pe_in_pk_rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.027 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0944 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 33.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3328 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1304 LAYER M4 ; 
    ANTENNAMAXAREACAR 73.3277 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.737551 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.72792 LAYER V4 ;
  END pe_in_pk_rdb_addr__3_
  PIN pe_in_pk_rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 44.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4472 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.472 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.0791 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.657821 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.6983 LAYER V4 ;
  END pe_in_pk_rdb_addr__2_
  PIN pe_in_pk_rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 6.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0606 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7992 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0901 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.1 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.15015 LAYER V3 ;
  END pe_in_pk_rdb_addr__1_
  PIN pe_in_pk_rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 11.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.3588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.193207 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.606061 LAYER V3 ;
  END pe_in_pk_rdb_addr__0_
  PIN pe_out_pk_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0592 LAYER M3 ;
  END pe_out_pk_PE_state__2_
  PIN pe_out_pk_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 3.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0192 LAYER M3 ;
  END pe_out_pk_PE_state__1_
  PIN pe_out_pk_PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
  END pe_out_pk_PE_state__0_
  PIN pe_out_pk_data__7_ 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M3 ;
  END pe_out_pk_data__7_
  PIN pe_out_pk_data__6_ 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0408 LAYER M3 ;
  END pe_out_pk_data__6_
  PIN pe_out_pk_data__5_ 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER M3 ;
  END pe_out_pk_data__5_
  PIN pe_out_pk_data__4_ 
    ANTENNAPARTIALMETALAREA 5.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0456 LAYER M3 ;
  END pe_out_pk_data__4_
  PIN pe_out_pk_data__3_ 
    ANTENNAPARTIALMETALAREA 4.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0454 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0856 LAYER M3 ;
  END pe_out_pk_data__3_
  PIN pe_out_pk_data__2_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 12.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1296 LAYER M3 ;
  END pe_out_pk_data__2_
  PIN pe_out_pk_data__1_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 16.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1672 LAYER M3 ;
  END pe_out_pk_data__1_
  PIN pe_out_pk_data__0_ 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0142 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 20.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.208 LAYER M3 ;
  END pe_out_pk_data__0_
END PE_top

END LIBRARY
