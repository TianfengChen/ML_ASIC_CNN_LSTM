

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO PE_POOL_top 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8352 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.93391 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0301485 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.191571 LAYER V3 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 1.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.73764 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0287389 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.190114 LAYER V3 ;
  END reset
  PIN pe_in_pk_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.256 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.16603 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__2_
  PIN pe_in_pk_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 134.487 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.35833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__1_
  PIN pe_in_pk_PE_state__0_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.37115 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__0_
  PIN pe_in_pk_A__3__7_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 123.269 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.23974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__7_
  PIN pe_in_pk_A__3__6_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0897 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.367949 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__6_
  PIN pe_in_pk_A__3__5_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9615 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__5_
  PIN pe_in_pk_A__3__4_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.40641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__4_
  PIN pe_in_pk_A__3__3_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.432051 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__3_
  PIN pe_in_pk_A__3__2_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.508974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__2_
  PIN pe_in_pk_A__3__1_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.7564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.534615 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__1_
  PIN pe_in_pk_A__3__0_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0208 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 46.6667 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.486538 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__3__0_
  PIN pe_in_pk_A__2__7_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.7564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.534615 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__7_
  PIN pe_in_pk_A__2__6_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 22.3077 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.242949 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__2__6_
  PIN pe_in_pk_A__2__5_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.7821 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.444872 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__5_
  PIN pe_in_pk_A__2__4_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.355128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__4_
  PIN pe_in_pk_A__2__3_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__3_
  PIN pe_in_pk_A__2__2_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.9615 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__2_
  PIN pe_in_pk_A__2__1_ 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0142 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.5256 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.342308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__1_
  PIN pe_in_pk_A__2__0_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__0_
  PIN pe_in_pk_A__1__7_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.355128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__7_
  PIN pe_in_pk_A__1__6_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__6_
  PIN pe_in_pk_A__1__5_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__5_
  PIN pe_in_pk_A__1__4_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6795 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.303846 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__4_
  PIN pe_in_pk_A__1__3_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.432051 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__3_
  PIN pe_in_pk_A__1__2_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.6923 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.396795 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__1__2_
  PIN pe_in_pk_A__1__1_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.6026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.573077 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__1_
  PIN pe_in_pk_A__1__0_ 
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0198 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0176 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 35.1282 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.371154 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__1__0_
  PIN pe_in_pk_A__0__7_ 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.023 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0296 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.3333 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.653205 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__0__7_
  PIN pe_in_pk_A__0__6_ 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0262 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.9872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.483333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__6_
  PIN pe_in_pk_A__0__5_ 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.432051 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__5_
  PIN pe_in_pk_A__0__4_ 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 55.3205 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.560256 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__4_
  PIN pe_in_pk_A__0__3_ 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.5128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.512179 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__3_
  PIN pe_in_pk_A__0__2_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.3462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.470513 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__2_
  PIN pe_in_pk_A__0__1_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.3462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.470513 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__1_
  PIN pe_in_pk_A__0__0_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__0_
  PIN pe_in_pk_wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 84.4872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.858333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_wrb_data__7_
  PIN pe_in_pk_wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.4214 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.280503 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER V3 ;
  END pe_in_pk_wrb_data__6_
  PIN pe_in_pk_wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.409615 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_wrb_data__5_
  PIN pe_in_pk_wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 31.6026 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.316667 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END pe_in_pk_wrb_data__4_
  PIN pe_in_pk_wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.3846 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.217308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_wrb_data__3_
  PIN pe_in_pk_wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.327 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.12956 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER V3 ;
  END pe_in_pk_wrb_data__2_
  PIN pe_in_pk_wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.6981 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.12327 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER V3 ;
  END pe_in_pk_wrb_data__1_
  PIN pe_in_pk_wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 1.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.3846 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.217308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_wrb_data__0_
  PIN pe_in_pk_wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 1.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0126 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7248 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.29077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0687978 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.854701 LAYER V3 ;
  END pe_in_pk_wrb_addr__3_
  PIN pe_in_pk_wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0288 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.3846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.245513 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAGATEAREA 0.1248 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.3462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.258333 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.961538 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M4 ;
    ANTENNAGATEAREA 1.1808 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.4762 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.340312 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.961538 LAYER V4 ;
  END pe_in_pk_wrb_addr__2_
  PIN pe_in_pk_wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.264103 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 9.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0928 LAYER M4 ;
    ANTENNAGATEAREA 0.8784 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.1146 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.369749 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V4 ;
  END pe_in_pk_wrb_addr__1_
  PIN pe_in_pk_wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.7644 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.415385 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAMAXCUTCAR 0.961538 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0968 LAYER M4 ;
    ANTENNAGATEAREA 0.828 LAYER M4 ; 
    ANTENNAMAXAREACAR 52.3586 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.532293 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.961538 LAYER V4 ;
  END pe_in_pk_wrb_addr__0_
  PIN pe_in_pk_wrb__3_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M2 ; 
    ANTENNAMAXAREACAR 6.28455 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.0635501 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.135501 LAYER V2 ;
  END pe_in_pk_wrb__3_
  PIN pe_in_pk_wrb__2_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.4173 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.107588 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.406504 LAYER V3 ;
  END pe_in_pk_wrb__2_
  PIN pe_in_pk_wrb__1_ 
    ANTENNAPARTIALMETALAREA 0.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0078 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.1734 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.205149 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.406504 LAYER V3 ;
  END pe_in_pk_wrb__1_
  PIN pe_in_pk_wrb__0_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.0894 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.194309 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.406504 LAYER V3 ;
  END pe_in_pk_wrb__0_
  PIN pe_in_pk_rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.156 LAYER M3 ; 
    ANTENNAMAXAREACAR 61.1359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.616923 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAMAXCUTCAR 2.05128 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0296 LAYER M4 ;
    ANTENNAGATEAREA 0.3192 LAYER M4 ; 
    ANTENNAMAXAREACAR 70.2838 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.709655 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.05128 LAYER V4 ;
  END pe_in_pk_rdb_addr__3_
  PIN pe_in_pk_rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.108 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.264 LAYER M3 ; 
    ANTENNAMAXAREACAR 49.4409 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.494848 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.606061 LAYER V3 ;
  END pe_in_pk_rdb_addr__2_
  PIN pe_in_pk_rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1632 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8592 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6672 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.41238 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_rdb_addr__1_
  PIN pe_in_pk_rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.264 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.5318 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.585758 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.454545 LAYER V3 ;
  END pe_in_pk_rdb_addr__0_
  PIN pk_out_PE_state__2_ 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0958 LAYER M3 ;
  END pk_out_PE_state__2_
  PIN pk_out_PE_state__1_ 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1 LAYER M3 ;
  END pk_out_PE_state__1_
  PIN pk_out_PE_state__0_ 
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1006 LAYER M3 ;
  END pk_out_PE_state__0_
  PIN pk_out_data__7_ 
  END pk_out_data__7_
  PIN pk_out_data__6_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0646 LAYER M3 ;
  END pk_out_data__6_
  PIN pk_out_data__5_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0696 LAYER M3 ;
  END pk_out_data__5_
  PIN pk_out_data__4_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0694 LAYER M3 ;
  END pk_out_data__4_
  PIN pk_out_data__3_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0694 LAYER M3 ;
  END pk_out_data__3_
  PIN pk_out_data__2_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0678 LAYER M3 ;
  END pk_out_data__2_
  PIN pk_out_data__1_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER M3 ;
  END pk_out_data__1_
  PIN pk_out_data__0_ 
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0694 LAYER M3 ;
  END pk_out_data__0_
END PE_POOL_top

END LIBRARY
