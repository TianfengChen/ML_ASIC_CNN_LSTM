VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LDO_Top_lef
  CLASS BLOCK ;
  ORIGIN 0.34 96.4 ;
  FOREIGN LDO_Top_lef -0.34 -96.4 ;
  SIZE 125.45 BY 46 ;
  SYMMETRY X Y R90 ;
  PIN SW[2]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 22.94 -50.6 23.14 -50.4 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.68 -62.45 23.4 -61.73 ;
      LAYER M2 ;
        RECT 22.74 -62.39 23.34 -61.79 ;
      LAYER V1 ;
        RECT 22.74 -61.99 22.94 -61.79 ;
        RECT 22.74 -62.39 22.94 -62.19 ;
        RECT 23.14 -61.99 23.34 -61.79 ;
        RECT 23.14 -62.39 23.34 -62.19 ;
      LAYER V2 ;
        RECT 22.74 -61.99 22.94 -61.79 ;
        RECT 22.74 -62.39 22.94 -62.19 ;
        RECT 23.14 -61.99 23.34 -61.79 ;
        RECT 23.14 -62.39 23.34 -62.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -62 24.6 -61.84 ;
    END
  END SW[2]
  PIN SW[1]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 22.19 -50.6 22.39 -50.4 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.93 -58.78 22.65 -58.06 ;
      LAYER M2 ;
        RECT 21.99 -58.72 22.59 -58.12 ;
      LAYER V1 ;
        RECT 21.99 -58.32 22.19 -58.12 ;
        RECT 21.99 -58.72 22.19 -58.52 ;
        RECT 22.39 -58.32 22.59 -58.12 ;
        RECT 22.39 -58.72 22.59 -58.52 ;
      LAYER V2 ;
        RECT 21.99 -58.32 22.19 -58.12 ;
        RECT 21.99 -58.72 22.19 -58.52 ;
        RECT 22.39 -58.32 22.59 -58.12 ;
        RECT 22.39 -58.72 22.59 -58.52 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -58.64 24.6 -58.48 ;
    END
  END SW[1]
  PIN SW[0]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 21.42 -50.6 21.62 -50.4 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.16 -55.07 21.88 -54.35 ;
      LAYER M2 ;
        RECT 21.22 -55.01 21.82 -54.41 ;
      LAYER V1 ;
        RECT 21.22 -54.61 21.42 -54.41 ;
        RECT 21.22 -55.01 21.42 -54.81 ;
        RECT 21.62 -54.61 21.82 -54.41 ;
        RECT 21.62 -55.01 21.82 -54.81 ;
      LAYER V2 ;
        RECT 21.22 -54.61 21.42 -54.41 ;
        RECT 21.22 -55.01 21.42 -54.81 ;
        RECT 21.62 -54.61 21.82 -54.41 ;
        RECT 21.62 -55.01 21.82 -54.81 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.44 -54.8 24.6 -54.64 ;
    END
  END SW[0]
  PIN VB
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 47.82 -96.4 48.22 -96 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.8 -68.77 47.04 -68.53 ;
    END
  END VB
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 34.05 -53 35.05 -52.02 ;
        RECT 35.02 -53.02 35.05 -52.02 ;
        RECT 34.05 -53.02 34.12 -52.02 ;
      LAYER V2 ;
        RECT 34.05 -52.22 34.25 -52.02 ;
        RECT 34.05 -52.62 34.25 -52.42 ;
        RECT 34.05 -53.02 34.25 -52.82 ;
        RECT 34.45 -52.22 34.65 -52.02 ;
        RECT 34.45 -52.62 34.65 -52.42 ;
        RECT 34.45 -53.02 34.65 -52.82 ;
        RECT 34.85 -52.22 35.05 -52.02 ;
        RECT 34.85 -52.62 35.05 -52.42 ;
        RECT 34.85 -53.02 35.05 -52.82 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.48 -54.26 28.76 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.44 -54.26 29.72 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.4 -54.26 30.68 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.36 -54.26 31.64 -54 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4 -53.95 34.74 -53.78 ;
      LAYER V1 ;
        RECT 34.47 -54.02 34.67 -53.82 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.12 -90.61 65.38 -90.37 ;
      LAYER V1 ;
        RECT 65.15 -90.55 65.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.08 -90.61 66.34 -90.37 ;
      LAYER V1 ;
        RECT 66.11 -90.55 66.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.04 -90.61 67.3 -90.37 ;
      LAYER V1 ;
        RECT 67.07 -90.55 67.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68 -90.61 68.26 -90.37 ;
      LAYER V1 ;
        RECT 68.03 -90.55 68.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.96 -90.61 69.22 -90.37 ;
      LAYER V1 ;
        RECT 68.99 -90.55 69.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.92 -90.61 70.18 -90.37 ;
      LAYER V1 ;
        RECT 69.95 -90.55 70.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.88 -90.61 71.14 -90.37 ;
      LAYER V1 ;
        RECT 70.91 -90.55 71.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.84 -90.61 72.1 -90.37 ;
      LAYER V1 ;
        RECT 71.87 -90.55 72.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.8 -90.61 73.06 -90.37 ;
      LAYER V1 ;
        RECT 72.83 -90.55 73.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.76 -90.61 74.02 -90.37 ;
      LAYER V1 ;
        RECT 73.79 -90.55 73.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.72 -90.61 74.98 -90.37 ;
      LAYER V1 ;
        RECT 74.75 -90.55 74.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.68 -90.61 75.94 -90.37 ;
      LAYER V1 ;
        RECT 75.71 -90.55 75.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.64 -90.61 76.9 -90.37 ;
      LAYER V1 ;
        RECT 76.67 -90.55 76.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.6 -90.61 77.86 -90.37 ;
      LAYER V1 ;
        RECT 77.63 -90.55 77.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.56 -90.61 78.82 -90.37 ;
      LAYER V1 ;
        RECT 78.59 -90.55 78.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.52 -90.61 79.78 -90.37 ;
      LAYER V1 ;
        RECT 79.55 -90.55 79.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.48 -90.61 80.74 -90.37 ;
      LAYER V1 ;
        RECT 80.51 -90.55 80.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.44 -90.61 81.7 -90.37 ;
      LAYER V1 ;
        RECT 81.47 -90.55 81.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.4 -90.61 82.66 -90.37 ;
      LAYER V1 ;
        RECT 82.43 -90.55 82.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.36 -90.61 83.62 -90.37 ;
      LAYER V1 ;
        RECT 83.39 -90.55 83.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.32 -90.61 84.58 -90.37 ;
      LAYER V1 ;
        RECT 84.35 -90.55 84.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.28 -90.61 85.54 -90.37 ;
      LAYER V1 ;
        RECT 85.31 -90.55 85.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.24 -90.61 86.5 -90.37 ;
      LAYER V1 ;
        RECT 86.27 -90.55 86.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.2 -90.61 87.46 -90.37 ;
      LAYER V1 ;
        RECT 87.23 -90.55 87.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.16 -90.61 88.42 -90.37 ;
      LAYER V1 ;
        RECT 88.19 -90.55 88.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.12 -90.61 89.38 -90.37 ;
      LAYER V1 ;
        RECT 89.15 -90.55 89.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.08 -90.61 90.34 -90.37 ;
      LAYER V1 ;
        RECT 90.11 -90.55 90.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.04 -90.61 91.3 -90.37 ;
      LAYER V1 ;
        RECT 91.07 -90.55 91.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92 -90.61 92.26 -90.37 ;
      LAYER V1 ;
        RECT 92.03 -90.55 92.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.96 -90.61 93.22 -90.37 ;
      LAYER V1 ;
        RECT 92.99 -90.55 93.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.92 -90.61 94.18 -90.37 ;
      LAYER V1 ;
        RECT 93.95 -90.55 94.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.88 -90.61 95.14 -90.37 ;
      LAYER V1 ;
        RECT 94.91 -90.55 95.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.84 -90.61 96.1 -90.37 ;
      LAYER V1 ;
        RECT 95.87 -90.55 96.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.8 -90.61 97.06 -90.37 ;
      LAYER V1 ;
        RECT 96.83 -90.55 97.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.76 -90.61 98.02 -90.37 ;
      LAYER V1 ;
        RECT 97.79 -90.55 97.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.72 -90.61 98.98 -90.37 ;
      LAYER V1 ;
        RECT 98.75 -90.55 98.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.68 -90.61 99.94 -90.37 ;
      LAYER V1 ;
        RECT 99.71 -90.55 99.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.64 -90.61 100.9 -90.37 ;
      LAYER V1 ;
        RECT 100.67 -90.55 100.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.6 -90.61 101.86 -90.37 ;
      LAYER V1 ;
        RECT 101.63 -90.55 101.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.56 -90.61 102.82 -90.37 ;
      LAYER V1 ;
        RECT 102.59 -90.55 102.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.52 -90.61 103.78 -90.37 ;
      LAYER V1 ;
        RECT 103.55 -90.55 103.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.48 -90.61 104.74 -90.37 ;
      LAYER V1 ;
        RECT 104.51 -90.55 104.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.44 -90.61 105.7 -90.37 ;
      LAYER V1 ;
        RECT 105.47 -90.55 105.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.4 -90.61 106.66 -90.37 ;
      LAYER V1 ;
        RECT 106.43 -90.55 106.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.36 -90.61 107.62 -90.37 ;
      LAYER V1 ;
        RECT 107.39 -90.55 107.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.32 -90.61 108.58 -90.37 ;
      LAYER V1 ;
        RECT 108.35 -90.55 108.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.28 -90.61 109.54 -90.37 ;
      LAYER V1 ;
        RECT 109.31 -90.55 109.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.24 -90.61 110.5 -90.37 ;
      LAYER V1 ;
        RECT 110.27 -90.55 110.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.2 -90.61 111.46 -90.37 ;
      LAYER V1 ;
        RECT 111.23 -90.55 111.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.16 -90.61 112.42 -90.37 ;
      LAYER V1 ;
        RECT 112.19 -90.55 112.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.12 -90.61 113.38 -90.37 ;
      LAYER V1 ;
        RECT 113.15 -90.55 113.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.08 -90.61 114.34 -90.37 ;
      LAYER V1 ;
        RECT 114.11 -90.55 114.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.04 -90.61 115.3 -90.37 ;
      LAYER V1 ;
        RECT 115.07 -90.55 115.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116 -90.61 116.26 -90.37 ;
      LAYER V1 ;
        RECT 116.03 -90.55 116.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.96 -90.61 117.22 -90.37 ;
      LAYER V1 ;
        RECT 116.99 -90.55 117.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.92 -90.61 118.18 -90.37 ;
      LAYER V1 ;
        RECT 117.95 -90.55 118.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.88 -90.61 119.14 -90.37 ;
      LAYER V1 ;
        RECT 118.91 -90.55 119.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.84 -90.61 120.1 -90.37 ;
      LAYER V1 ;
        RECT 119.87 -90.55 120.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.8 -90.61 121.06 -90.37 ;
      LAYER V1 ;
        RECT 120.83 -90.55 121.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.76 -90.61 122.02 -90.37 ;
      LAYER V1 ;
        RECT 121.79 -90.55 121.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.72 -90.61 122.98 -90.37 ;
      LAYER V1 ;
        RECT 122.75 -90.55 122.95 -90.35 ;
    END
  END DVDD
  PIN AVDD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M2 ;
        RECT 7.38 -61.17 9.38 -59.17 ;
      LAYER V1 ;
        RECT 7.38 -59.45 7.58 -59.25 ;
        RECT 7.38 -59.85 7.58 -59.65 ;
        RECT 7.38 -60.25 7.58 -60.05 ;
        RECT 7.38 -60.65 7.58 -60.45 ;
        RECT 7.38 -61.05 7.58 -60.85 ;
        RECT 7.78 -59.45 7.98 -59.25 ;
        RECT 7.78 -59.85 7.98 -59.65 ;
        RECT 7.78 -60.25 7.98 -60.05 ;
        RECT 7.78 -60.65 7.98 -60.45 ;
        RECT 7.78 -61.05 7.98 -60.85 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.13 -68.33 36.43 -68.03 ;
      LAYER V1 ;
        RECT 36.2 -68.29 36.4 -68.09 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.55 -65.95 101.55 -50.95 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.9 -69.65 124.78 -68.77 ;
      LAYER V1 ;
        RECT 123.94 -69.09 124.14 -68.89 ;
        RECT 123.94 -69.53 124.14 -69.33 ;
        RECT 124.34 -69.09 124.54 -68.89 ;
        RECT 124.34 -69.53 124.54 -69.33 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.01 -60.63 4.17 -60.47 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.32 -61.91 8.04 -61.19 ;
      LAYER M2 ;
        RECT 7.38 -61.85 7.98 -61.25 ;
      LAYER V1 ;
        RECT 7.38 -61.45 7.58 -61.25 ;
        RECT 7.38 -61.85 7.58 -61.65 ;
        RECT 7.78 -61.45 7.98 -61.25 ;
        RECT 7.78 -61.85 7.98 -61.65 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -55.47 24.44 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -62.67 24.44 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.98 -56.88 24.46 -56.4 ;
      LAYER M2 ;
        RECT 24.08 -57.14 24.68 -56.54 ;
      LAYER V1 ;
        RECT 24.08 -56.74 24.28 -56.54 ;
        RECT 24.48 -56.74 24.68 -56.54 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.98 -64.08 24.46 -63.6 ;
      LAYER V1 ;
        RECT 24.08 -63.94 24.28 -63.74 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -55.47 25.4 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -62.67 25.4 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.67 -69.21 25.93 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -55.47 26.36 -55.19 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -62.67 26.36 -62.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -55.58 26.84 -55.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -62.78 26.84 -62.5 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -55.58 27.8 -55.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -62.78 27.8 -62.5 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.33 -69.42 28.8 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.05 -68.33 31.35 -68.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.05 -69.21 32.31 -68.95 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.55 -68.35 36.87 -68.03 ;
      LAYER V1 ;
        RECT 36.6 -68.29 36.8 -68.09 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.64 -69.59 47.8 -69.43 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.31 -69.16 51.63 -68.84 ;
        RECT 51.19 -69.3 51.45 -69.04 ;
      LAYER V1 ;
        RECT 51.37 -69.1 51.57 -68.9 ;
        RECT 51.37 -69.5 51.57 -69.3 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.8 -69.38 54.14 -69.04 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.44 -69.3 56.7 -69.04 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.32 -69.65 64.2 -68.77 ;
      LAYER V1 ;
        RECT 63.54 -69.09 63.74 -68.89 ;
        RECT 63.54 -69.53 63.74 -69.33 ;
        RECT 63.94 -69.09 64.14 -68.89 ;
        RECT 63.94 -69.53 64.14 -69.33 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.32 -92.61 64.2 -91.73 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6 -90.61 65.86 -90.35 ;
      LAYER M2 ;
        RECT 65.6 -90.61 65.86 -90.35 ;
      LAYER V1 ;
        RECT 65.63 -90.55 65.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.56 -90.61 66.82 -90.35 ;
      LAYER M2 ;
        RECT 66.56 -90.61 66.82 -90.35 ;
      LAYER V1 ;
        RECT 66.59 -90.55 66.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.52 -90.61 67.78 -90.35 ;
      LAYER M2 ;
        RECT 67.52 -90.61 67.78 -90.35 ;
      LAYER V1 ;
        RECT 67.55 -90.55 67.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.48 -90.61 68.74 -90.35 ;
      LAYER M2 ;
        RECT 68.48 -90.61 68.74 -90.35 ;
      LAYER V1 ;
        RECT 68.51 -90.55 68.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.44 -90.61 69.7 -90.35 ;
      LAYER M2 ;
        RECT 69.44 -90.61 69.7 -90.35 ;
      LAYER V1 ;
        RECT 69.47 -90.55 69.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4 -90.61 70.66 -90.35 ;
      LAYER M2 ;
        RECT 70.4 -90.61 70.66 -90.35 ;
      LAYER V1 ;
        RECT 70.43 -90.55 70.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.36 -90.61 71.62 -90.35 ;
      LAYER M2 ;
        RECT 71.36 -90.61 71.62 -90.35 ;
      LAYER V1 ;
        RECT 71.39 -90.55 71.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.32 -90.61 72.58 -90.35 ;
      LAYER M2 ;
        RECT 72.32 -90.61 72.58 -90.35 ;
      LAYER V1 ;
        RECT 72.35 -90.55 72.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.28 -90.61 73.54 -90.35 ;
      LAYER M2 ;
        RECT 73.28 -90.61 73.54 -90.35 ;
      LAYER V1 ;
        RECT 73.31 -90.55 73.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.24 -90.61 74.5 -90.35 ;
      LAYER M2 ;
        RECT 74.24 -90.61 74.5 -90.35 ;
      LAYER V1 ;
        RECT 74.27 -90.55 74.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2 -90.61 75.46 -90.35 ;
      LAYER M2 ;
        RECT 75.2 -90.61 75.46 -90.35 ;
      LAYER V1 ;
        RECT 75.23 -90.55 75.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.16 -90.61 76.42 -90.35 ;
      LAYER M2 ;
        RECT 76.16 -90.61 76.42 -90.35 ;
      LAYER V1 ;
        RECT 76.19 -90.55 76.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.12 -90.61 77.38 -90.35 ;
      LAYER M2 ;
        RECT 77.12 -90.61 77.38 -90.35 ;
      LAYER V1 ;
        RECT 77.15 -90.55 77.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.08 -90.61 78.34 -90.35 ;
      LAYER M2 ;
        RECT 78.08 -90.61 78.34 -90.35 ;
      LAYER V1 ;
        RECT 78.11 -90.55 78.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.04 -90.61 79.3 -90.35 ;
      LAYER M2 ;
        RECT 79.04 -90.61 79.3 -90.35 ;
      LAYER V1 ;
        RECT 79.07 -90.55 79.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80 -90.61 80.26 -90.35 ;
      LAYER M2 ;
        RECT 80 -90.61 80.26 -90.35 ;
      LAYER V1 ;
        RECT 80.03 -90.55 80.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.96 -90.61 81.22 -90.35 ;
      LAYER M2 ;
        RECT 80.96 -90.61 81.22 -90.35 ;
      LAYER V1 ;
        RECT 80.99 -90.55 81.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.92 -90.61 82.18 -90.35 ;
      LAYER M2 ;
        RECT 81.92 -90.61 82.18 -90.35 ;
      LAYER V1 ;
        RECT 81.95 -90.55 82.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.88 -90.61 83.14 -90.35 ;
      LAYER M2 ;
        RECT 82.88 -90.61 83.14 -90.35 ;
      LAYER V1 ;
        RECT 82.91 -90.55 83.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.84 -90.61 84.1 -90.35 ;
      LAYER M2 ;
        RECT 83.84 -90.61 84.1 -90.35 ;
      LAYER V1 ;
        RECT 83.87 -90.55 84.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8 -90.61 85.06 -90.35 ;
      LAYER M2 ;
        RECT 84.8 -90.61 85.06 -90.35 ;
      LAYER V1 ;
        RECT 84.83 -90.55 85.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.76 -90.61 86.02 -90.35 ;
      LAYER M2 ;
        RECT 85.76 -90.61 86.02 -90.35 ;
      LAYER V1 ;
        RECT 85.79 -90.55 85.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.72 -90.61 86.98 -90.35 ;
      LAYER M2 ;
        RECT 86.72 -90.61 86.98 -90.35 ;
      LAYER V1 ;
        RECT 86.75 -90.55 86.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.68 -90.61 87.94 -90.35 ;
      LAYER M2 ;
        RECT 87.68 -90.61 87.94 -90.35 ;
      LAYER V1 ;
        RECT 87.71 -90.55 87.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.64 -90.61 88.9 -90.35 ;
      LAYER M2 ;
        RECT 88.64 -90.61 88.9 -90.35 ;
      LAYER V1 ;
        RECT 88.67 -90.55 88.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.6 -90.61 89.86 -90.35 ;
      LAYER M2 ;
        RECT 89.6 -90.61 89.86 -90.35 ;
      LAYER V1 ;
        RECT 89.63 -90.55 89.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.56 -90.61 90.82 -90.35 ;
      LAYER M2 ;
        RECT 90.56 -90.61 90.82 -90.35 ;
      LAYER V1 ;
        RECT 90.59 -90.55 90.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.52 -90.61 91.78 -90.35 ;
      LAYER M2 ;
        RECT 91.52 -90.61 91.78 -90.35 ;
      LAYER V1 ;
        RECT 91.55 -90.55 91.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.48 -90.61 92.74 -90.35 ;
      LAYER M2 ;
        RECT 92.48 -90.61 92.74 -90.35 ;
      LAYER V1 ;
        RECT 92.51 -90.55 92.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.44 -90.61 93.7 -90.35 ;
      LAYER M2 ;
        RECT 93.44 -90.61 93.7 -90.35 ;
      LAYER V1 ;
        RECT 93.47 -90.55 93.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4 -90.61 94.66 -90.35 ;
      LAYER M2 ;
        RECT 94.4 -90.61 94.66 -90.35 ;
      LAYER V1 ;
        RECT 94.43 -90.55 94.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.36 -90.61 95.62 -90.35 ;
      LAYER M2 ;
        RECT 95.36 -90.61 95.62 -90.35 ;
      LAYER V1 ;
        RECT 95.39 -90.55 95.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.32 -90.61 96.58 -90.35 ;
      LAYER M2 ;
        RECT 96.32 -90.61 96.58 -90.35 ;
      LAYER V1 ;
        RECT 96.35 -90.55 96.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.28 -90.61 97.54 -90.35 ;
      LAYER M2 ;
        RECT 97.28 -90.61 97.54 -90.35 ;
      LAYER V1 ;
        RECT 97.31 -90.55 97.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.24 -90.61 98.5 -90.35 ;
      LAYER M2 ;
        RECT 98.24 -90.61 98.5 -90.35 ;
      LAYER V1 ;
        RECT 98.27 -90.55 98.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.2 -90.61 99.46 -90.35 ;
      LAYER M2 ;
        RECT 99.2 -90.61 99.46 -90.35 ;
      LAYER V1 ;
        RECT 99.23 -90.55 99.43 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.16 -90.61 100.42 -90.35 ;
      LAYER M2 ;
        RECT 100.16 -90.61 100.42 -90.35 ;
      LAYER V1 ;
        RECT 100.19 -90.55 100.39 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.12 -90.61 101.38 -90.35 ;
      LAYER M2 ;
        RECT 101.12 -90.61 101.38 -90.35 ;
      LAYER V1 ;
        RECT 101.15 -90.55 101.35 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.08 -90.61 102.34 -90.35 ;
      LAYER M2 ;
        RECT 102.08 -90.61 102.34 -90.35 ;
      LAYER V1 ;
        RECT 102.11 -90.55 102.31 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.04 -90.61 103.3 -90.35 ;
      LAYER M2 ;
        RECT 103.04 -90.61 103.3 -90.35 ;
      LAYER V1 ;
        RECT 103.07 -90.55 103.27 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104 -90.61 104.26 -90.35 ;
      LAYER M2 ;
        RECT 104 -90.61 104.26 -90.35 ;
      LAYER V1 ;
        RECT 104.03 -90.55 104.23 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.96 -90.61 105.22 -90.35 ;
      LAYER M2 ;
        RECT 104.96 -90.61 105.22 -90.35 ;
      LAYER V1 ;
        RECT 104.99 -90.55 105.19 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.92 -90.61 106.18 -90.35 ;
      LAYER M2 ;
        RECT 105.92 -90.61 106.18 -90.35 ;
      LAYER V1 ;
        RECT 105.95 -90.55 106.15 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.88 -90.61 107.14 -90.35 ;
      LAYER M2 ;
        RECT 106.88 -90.61 107.14 -90.35 ;
      LAYER V1 ;
        RECT 106.91 -90.55 107.11 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.84 -90.61 108.1 -90.35 ;
      LAYER M2 ;
        RECT 107.84 -90.61 108.1 -90.35 ;
      LAYER V1 ;
        RECT 107.87 -90.55 108.07 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.8 -90.61 109.06 -90.35 ;
      LAYER M2 ;
        RECT 108.8 -90.61 109.06 -90.35 ;
      LAYER V1 ;
        RECT 108.83 -90.55 109.03 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.76 -90.61 110.02 -90.35 ;
      LAYER M2 ;
        RECT 109.76 -90.61 110.02 -90.35 ;
      LAYER V1 ;
        RECT 109.79 -90.55 109.99 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.72 -90.61 110.98 -90.35 ;
      LAYER M2 ;
        RECT 110.72 -90.61 110.98 -90.35 ;
      LAYER V1 ;
        RECT 110.75 -90.55 110.95 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.68 -90.61 111.94 -90.35 ;
      LAYER M2 ;
        RECT 111.68 -90.61 111.94 -90.35 ;
      LAYER V1 ;
        RECT 111.71 -90.55 111.91 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.64 -90.61 112.9 -90.35 ;
      LAYER M2 ;
        RECT 112.64 -90.61 112.9 -90.35 ;
      LAYER V1 ;
        RECT 112.67 -90.55 112.87 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.6 -90.61 113.86 -90.35 ;
      LAYER M2 ;
        RECT 113.6 -90.61 113.86 -90.35 ;
      LAYER V1 ;
        RECT 113.63 -90.55 113.83 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.56 -90.61 114.82 -90.35 ;
      LAYER M2 ;
        RECT 114.56 -90.61 114.82 -90.35 ;
      LAYER V1 ;
        RECT 114.59 -90.55 114.79 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.52 -90.61 115.78 -90.35 ;
      LAYER M2 ;
        RECT 115.52 -90.61 115.78 -90.35 ;
      LAYER V1 ;
        RECT 115.55 -90.55 115.75 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.48 -90.61 116.74 -90.35 ;
      LAYER M2 ;
        RECT 116.48 -90.61 116.74 -90.35 ;
      LAYER V1 ;
        RECT 116.51 -90.55 116.71 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.44 -90.61 117.7 -90.35 ;
      LAYER M2 ;
        RECT 117.44 -90.61 117.7 -90.35 ;
      LAYER V1 ;
        RECT 117.47 -90.55 117.67 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.4 -90.61 118.66 -90.35 ;
      LAYER M2 ;
        RECT 118.4 -90.61 118.66 -90.35 ;
      LAYER V1 ;
        RECT 118.43 -90.55 118.63 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.36 -90.61 119.62 -90.35 ;
      LAYER M2 ;
        RECT 119.36 -90.61 119.62 -90.35 ;
      LAYER V1 ;
        RECT 119.39 -90.55 119.59 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.32 -90.61 120.58 -90.35 ;
      LAYER M2 ;
        RECT 120.32 -90.61 120.58 -90.35 ;
      LAYER V1 ;
        RECT 120.35 -90.55 120.55 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.28 -90.61 121.54 -90.35 ;
      LAYER M2 ;
        RECT 121.28 -90.61 121.54 -90.35 ;
      LAYER V1 ;
        RECT 121.31 -90.55 121.51 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.24 -90.61 122.5 -90.35 ;
      LAYER M2 ;
        RECT 122.24 -90.61 122.5 -90.35 ;
      LAYER V1 ;
        RECT 122.27 -90.55 122.47 -90.35 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.34 -92.61 124.78 -92.17 ;
    END
  END AVDD
  PIN VOUT
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M1 ;
        RECT 42.85 -82.58 43.15 -82.28 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.35 -85.91 43.51 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.05 -85.91 46.21 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.75 -85.91 48.91 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.45 -85.91 51.61 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.15 -85.91 54.31 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.85 -85.91 57.01 -85.75 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.47 -82.73 59.92 -82.28 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.32 -91.33 64.88 -90.77 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.32 -70.61 64.9 -70.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.38 -91.33 124 -90.71 ;
    END
  END VOUT
  PIN AVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER M3 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER M4 ;
        RECT 11.21 -78.61 21.57 -68.27 ;
      LAYER V3 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
      LAYER V1 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
      LAYER V2 ;
        RECT 11.25 -71.62 11.45 -71.42 ;
        RECT 11.25 -72.22 11.45 -72.02 ;
        RECT 11.25 -72.82 11.45 -72.62 ;
        RECT 11.25 -73.42 11.45 -73.22 ;
        RECT 11.25 -74.02 11.45 -73.82 ;
        RECT 11.25 -74.62 11.45 -74.42 ;
        RECT 11.25 -75.22 11.45 -75.02 ;
        RECT 11.25 -75.82 11.45 -75.62 ;
        RECT 11.25 -76.42 11.45 -76.22 ;
        RECT 11.25 -77.02 11.45 -76.82 ;
        RECT 11.25 -77.62 11.45 -77.42 ;
        RECT 11.25 -78.22 11.45 -78.02 ;
        RECT 11.73 -71.92 11.93 -71.72 ;
        RECT 11.73 -72.52 11.93 -72.32 ;
        RECT 11.73 -73.12 11.93 -72.92 ;
        RECT 11.73 -73.72 11.93 -73.52 ;
        RECT 11.73 -74.32 11.93 -74.12 ;
        RECT 11.73 -74.92 11.93 -74.72 ;
        RECT 11.73 -75.52 11.93 -75.32 ;
        RECT 11.73 -76.12 11.93 -75.92 ;
        RECT 11.73 -76.72 11.93 -76.52 ;
        RECT 11.73 -77.32 11.93 -77.12 ;
        RECT 11.73 -77.92 11.93 -77.72 ;
        RECT 11.73 -78.52 11.93 -78.32 ;
        RECT 11.79 -68.87 11.99 -68.67 ;
        RECT 11.79 -69.47 11.99 -69.27 ;
        RECT 11.79 -70.07 11.99 -69.87 ;
        RECT 11.79 -70.67 11.99 -70.47 ;
        RECT 12.21 -71.62 12.41 -71.42 ;
        RECT 12.21 -72.22 12.41 -72.02 ;
        RECT 12.21 -72.82 12.41 -72.62 ;
        RECT 12.21 -73.42 12.41 -73.22 ;
        RECT 12.21 -74.02 12.41 -73.82 ;
        RECT 12.21 -74.62 12.41 -74.42 ;
        RECT 12.21 -75.22 12.41 -75.02 ;
        RECT 12.21 -75.82 12.41 -75.62 ;
        RECT 12.21 -76.42 12.41 -76.22 ;
        RECT 12.21 -77.02 12.41 -76.82 ;
        RECT 12.21 -77.62 12.41 -77.42 ;
        RECT 12.21 -78.22 12.41 -78.02 ;
        RECT 12.39 -68.87 12.59 -68.67 ;
        RECT 12.39 -69.47 12.59 -69.27 ;
        RECT 12.39 -70.07 12.59 -69.87 ;
        RECT 12.39 -70.67 12.59 -70.47 ;
        RECT 12.69 -71.92 12.89 -71.72 ;
        RECT 12.69 -72.52 12.89 -72.32 ;
        RECT 12.69 -73.12 12.89 -72.92 ;
        RECT 12.69 -73.72 12.89 -73.52 ;
        RECT 12.69 -74.32 12.89 -74.12 ;
        RECT 12.69 -74.92 12.89 -74.72 ;
        RECT 12.69 -75.52 12.89 -75.32 ;
        RECT 12.69 -76.12 12.89 -75.92 ;
        RECT 12.69 -76.72 12.89 -76.52 ;
        RECT 12.69 -77.32 12.89 -77.12 ;
        RECT 12.69 -77.92 12.89 -77.72 ;
        RECT 12.69 -78.52 12.89 -78.32 ;
        RECT 12.99 -68.87 13.19 -68.67 ;
        RECT 12.99 -69.47 13.19 -69.27 ;
        RECT 12.99 -70.07 13.19 -69.87 ;
        RECT 12.99 -70.67 13.19 -70.47 ;
        RECT 13.17 -71.62 13.37 -71.42 ;
        RECT 13.17 -72.22 13.37 -72.02 ;
        RECT 13.17 -72.82 13.37 -72.62 ;
        RECT 13.17 -73.42 13.37 -73.22 ;
        RECT 13.17 -74.02 13.37 -73.82 ;
        RECT 13.17 -74.62 13.37 -74.42 ;
        RECT 13.17 -75.22 13.37 -75.02 ;
        RECT 13.17 -75.82 13.37 -75.62 ;
        RECT 13.17 -76.42 13.37 -76.22 ;
        RECT 13.17 -77.02 13.37 -76.82 ;
        RECT 13.17 -77.62 13.37 -77.42 ;
        RECT 13.17 -78.22 13.37 -78.02 ;
        RECT 13.59 -68.87 13.79 -68.67 ;
        RECT 13.59 -69.47 13.79 -69.27 ;
        RECT 13.59 -70.07 13.79 -69.87 ;
        RECT 13.59 -70.67 13.79 -70.47 ;
        RECT 13.65 -71.92 13.85 -71.72 ;
        RECT 13.65 -72.52 13.85 -72.32 ;
        RECT 13.65 -73.12 13.85 -72.92 ;
        RECT 13.65 -73.72 13.85 -73.52 ;
        RECT 13.65 -74.32 13.85 -74.12 ;
        RECT 13.65 -74.92 13.85 -74.72 ;
        RECT 13.65 -75.52 13.85 -75.32 ;
        RECT 13.65 -76.12 13.85 -75.92 ;
        RECT 13.65 -76.72 13.85 -76.52 ;
        RECT 13.65 -77.32 13.85 -77.12 ;
        RECT 13.65 -77.92 13.85 -77.72 ;
        RECT 13.65 -78.52 13.85 -78.32 ;
        RECT 14.13 -71.62 14.33 -71.42 ;
        RECT 14.13 -72.22 14.33 -72.02 ;
        RECT 14.13 -72.82 14.33 -72.62 ;
        RECT 14.13 -73.42 14.33 -73.22 ;
        RECT 14.13 -74.02 14.33 -73.82 ;
        RECT 14.13 -74.62 14.33 -74.42 ;
        RECT 14.13 -75.22 14.33 -75.02 ;
        RECT 14.13 -75.82 14.33 -75.62 ;
        RECT 14.13 -76.42 14.33 -76.22 ;
        RECT 14.13 -77.02 14.33 -76.82 ;
        RECT 14.13 -77.62 14.33 -77.42 ;
        RECT 14.13 -78.22 14.33 -78.02 ;
        RECT 14.19 -68.87 14.39 -68.67 ;
        RECT 14.19 -69.47 14.39 -69.27 ;
        RECT 14.19 -70.07 14.39 -69.87 ;
        RECT 14.19 -70.67 14.39 -70.47 ;
        RECT 14.61 -71.92 14.81 -71.72 ;
        RECT 14.61 -72.52 14.81 -72.32 ;
        RECT 14.61 -73.12 14.81 -72.92 ;
        RECT 14.61 -73.72 14.81 -73.52 ;
        RECT 14.61 -74.32 14.81 -74.12 ;
        RECT 14.61 -74.92 14.81 -74.72 ;
        RECT 14.61 -75.52 14.81 -75.32 ;
        RECT 14.61 -76.12 14.81 -75.92 ;
        RECT 14.61 -76.72 14.81 -76.52 ;
        RECT 14.61 -77.32 14.81 -77.12 ;
        RECT 14.61 -77.92 14.81 -77.72 ;
        RECT 14.61 -78.52 14.81 -78.32 ;
        RECT 14.79 -68.87 14.99 -68.67 ;
        RECT 14.79 -69.47 14.99 -69.27 ;
        RECT 14.79 -70.07 14.99 -69.87 ;
        RECT 14.79 -70.67 14.99 -70.47 ;
        RECT 15.09 -71.62 15.29 -71.42 ;
        RECT 15.09 -72.22 15.29 -72.02 ;
        RECT 15.09 -72.82 15.29 -72.62 ;
        RECT 15.09 -73.42 15.29 -73.22 ;
        RECT 15.09 -74.02 15.29 -73.82 ;
        RECT 15.09 -74.62 15.29 -74.42 ;
        RECT 15.09 -75.22 15.29 -75.02 ;
        RECT 15.09 -75.82 15.29 -75.62 ;
        RECT 15.09 -76.42 15.29 -76.22 ;
        RECT 15.09 -77.02 15.29 -76.82 ;
        RECT 15.09 -77.62 15.29 -77.42 ;
        RECT 15.09 -78.22 15.29 -78.02 ;
        RECT 15.39 -68.87 15.59 -68.67 ;
        RECT 15.39 -69.47 15.59 -69.27 ;
        RECT 15.39 -70.07 15.59 -69.87 ;
        RECT 15.39 -70.67 15.59 -70.47 ;
        RECT 15.57 -71.92 15.77 -71.72 ;
        RECT 15.57 -72.52 15.77 -72.32 ;
        RECT 15.57 -73.12 15.77 -72.92 ;
        RECT 15.57 -73.72 15.77 -73.52 ;
        RECT 15.57 -74.32 15.77 -74.12 ;
        RECT 15.57 -74.92 15.77 -74.72 ;
        RECT 15.57 -75.52 15.77 -75.32 ;
        RECT 15.57 -76.12 15.77 -75.92 ;
        RECT 15.57 -76.72 15.77 -76.52 ;
        RECT 15.57 -77.32 15.77 -77.12 ;
        RECT 15.57 -77.92 15.77 -77.72 ;
        RECT 15.57 -78.52 15.77 -78.32 ;
        RECT 15.99 -68.87 16.19 -68.67 ;
        RECT 15.99 -69.47 16.19 -69.27 ;
        RECT 15.99 -70.07 16.19 -69.87 ;
        RECT 15.99 -70.67 16.19 -70.47 ;
        RECT 16.05 -71.62 16.25 -71.42 ;
        RECT 16.05 -72.22 16.25 -72.02 ;
        RECT 16.05 -72.82 16.25 -72.62 ;
        RECT 16.05 -73.42 16.25 -73.22 ;
        RECT 16.05 -74.02 16.25 -73.82 ;
        RECT 16.05 -74.62 16.25 -74.42 ;
        RECT 16.05 -75.22 16.25 -75.02 ;
        RECT 16.05 -75.82 16.25 -75.62 ;
        RECT 16.05 -76.42 16.25 -76.22 ;
        RECT 16.05 -77.02 16.25 -76.82 ;
        RECT 16.05 -77.62 16.25 -77.42 ;
        RECT 16.05 -78.22 16.25 -78.02 ;
        RECT 16.53 -71.92 16.73 -71.72 ;
        RECT 16.53 -72.52 16.73 -72.32 ;
        RECT 16.53 -73.12 16.73 -72.92 ;
        RECT 16.53 -73.72 16.73 -73.52 ;
        RECT 16.53 -74.32 16.73 -74.12 ;
        RECT 16.53 -74.92 16.73 -74.72 ;
        RECT 16.53 -75.52 16.73 -75.32 ;
        RECT 16.53 -76.12 16.73 -75.92 ;
        RECT 16.53 -76.72 16.73 -76.52 ;
        RECT 16.53 -77.32 16.73 -77.12 ;
        RECT 16.53 -77.92 16.73 -77.72 ;
        RECT 16.53 -78.52 16.73 -78.32 ;
        RECT 16.59 -68.87 16.79 -68.67 ;
        RECT 16.59 -69.47 16.79 -69.27 ;
        RECT 16.59 -70.07 16.79 -69.87 ;
        RECT 16.59 -70.67 16.79 -70.47 ;
        RECT 17.01 -71.62 17.21 -71.42 ;
        RECT 17.01 -72.22 17.21 -72.02 ;
        RECT 17.01 -72.82 17.21 -72.62 ;
        RECT 17.01 -73.42 17.21 -73.22 ;
        RECT 17.01 -74.02 17.21 -73.82 ;
        RECT 17.01 -74.62 17.21 -74.42 ;
        RECT 17.01 -75.22 17.21 -75.02 ;
        RECT 17.01 -75.82 17.21 -75.62 ;
        RECT 17.01 -76.42 17.21 -76.22 ;
        RECT 17.01 -77.02 17.21 -76.82 ;
        RECT 17.01 -77.62 17.21 -77.42 ;
        RECT 17.01 -78.22 17.21 -78.02 ;
        RECT 17.19 -68.87 17.39 -68.67 ;
        RECT 17.19 -69.47 17.39 -69.27 ;
        RECT 17.19 -70.07 17.39 -69.87 ;
        RECT 17.19 -70.67 17.39 -70.47 ;
        RECT 17.49 -71.92 17.69 -71.72 ;
        RECT 17.49 -72.52 17.69 -72.32 ;
        RECT 17.49 -73.12 17.69 -72.92 ;
        RECT 17.49 -73.72 17.69 -73.52 ;
        RECT 17.49 -74.32 17.69 -74.12 ;
        RECT 17.49 -74.92 17.69 -74.72 ;
        RECT 17.49 -75.52 17.69 -75.32 ;
        RECT 17.49 -76.12 17.69 -75.92 ;
        RECT 17.49 -76.72 17.69 -76.52 ;
        RECT 17.49 -77.32 17.69 -77.12 ;
        RECT 17.49 -77.92 17.69 -77.72 ;
        RECT 17.49 -78.52 17.69 -78.32 ;
        RECT 17.79 -68.87 17.99 -68.67 ;
        RECT 17.79 -69.47 17.99 -69.27 ;
        RECT 17.79 -70.07 17.99 -69.87 ;
        RECT 17.79 -70.67 17.99 -70.47 ;
        RECT 17.97 -71.62 18.17 -71.42 ;
        RECT 17.97 -72.22 18.17 -72.02 ;
        RECT 17.97 -72.82 18.17 -72.62 ;
        RECT 17.97 -73.42 18.17 -73.22 ;
        RECT 17.97 -74.02 18.17 -73.82 ;
        RECT 17.97 -74.62 18.17 -74.42 ;
        RECT 17.97 -75.22 18.17 -75.02 ;
        RECT 17.97 -75.82 18.17 -75.62 ;
        RECT 17.97 -76.42 18.17 -76.22 ;
        RECT 17.97 -77.02 18.17 -76.82 ;
        RECT 17.97 -77.62 18.17 -77.42 ;
        RECT 17.97 -78.22 18.17 -78.02 ;
        RECT 18.39 -68.87 18.59 -68.67 ;
        RECT 18.39 -69.47 18.59 -69.27 ;
        RECT 18.39 -70.07 18.59 -69.87 ;
        RECT 18.39 -70.67 18.59 -70.47 ;
        RECT 18.45 -71.92 18.65 -71.72 ;
        RECT 18.45 -72.52 18.65 -72.32 ;
        RECT 18.45 -73.12 18.65 -72.92 ;
        RECT 18.45 -73.72 18.65 -73.52 ;
        RECT 18.45 -74.32 18.65 -74.12 ;
        RECT 18.45 -74.92 18.65 -74.72 ;
        RECT 18.45 -75.52 18.65 -75.32 ;
        RECT 18.45 -76.12 18.65 -75.92 ;
        RECT 18.45 -76.72 18.65 -76.52 ;
        RECT 18.45 -77.32 18.65 -77.12 ;
        RECT 18.45 -77.92 18.65 -77.72 ;
        RECT 18.45 -78.52 18.65 -78.32 ;
        RECT 18.93 -71.62 19.13 -71.42 ;
        RECT 18.93 -72.22 19.13 -72.02 ;
        RECT 18.93 -72.82 19.13 -72.62 ;
        RECT 18.93 -73.42 19.13 -73.22 ;
        RECT 18.93 -74.02 19.13 -73.82 ;
        RECT 18.93 -74.62 19.13 -74.42 ;
        RECT 18.93 -75.22 19.13 -75.02 ;
        RECT 18.93 -75.82 19.13 -75.62 ;
        RECT 18.93 -76.42 19.13 -76.22 ;
        RECT 18.93 -77.02 19.13 -76.82 ;
        RECT 18.93 -77.62 19.13 -77.42 ;
        RECT 18.93 -78.22 19.13 -78.02 ;
        RECT 18.99 -68.87 19.19 -68.67 ;
        RECT 18.99 -69.47 19.19 -69.27 ;
        RECT 18.99 -70.07 19.19 -69.87 ;
        RECT 18.99 -70.67 19.19 -70.47 ;
        RECT 19.41 -71.92 19.61 -71.72 ;
        RECT 19.41 -72.52 19.61 -72.32 ;
        RECT 19.41 -73.12 19.61 -72.92 ;
        RECT 19.41 -73.72 19.61 -73.52 ;
        RECT 19.41 -74.32 19.61 -74.12 ;
        RECT 19.41 -74.92 19.61 -74.72 ;
        RECT 19.41 -75.52 19.61 -75.32 ;
        RECT 19.41 -76.12 19.61 -75.92 ;
        RECT 19.41 -76.72 19.61 -76.52 ;
        RECT 19.41 -77.32 19.61 -77.12 ;
        RECT 19.41 -77.92 19.61 -77.72 ;
        RECT 19.41 -78.52 19.61 -78.32 ;
        RECT 19.59 -68.87 19.79 -68.67 ;
        RECT 19.59 -69.47 19.79 -69.27 ;
        RECT 19.59 -70.07 19.79 -69.87 ;
        RECT 19.59 -70.67 19.79 -70.47 ;
        RECT 19.89 -71.62 20.09 -71.42 ;
        RECT 19.89 -72.22 20.09 -72.02 ;
        RECT 19.89 -72.82 20.09 -72.62 ;
        RECT 19.89 -73.42 20.09 -73.22 ;
        RECT 19.89 -74.02 20.09 -73.82 ;
        RECT 19.89 -74.62 20.09 -74.42 ;
        RECT 19.89 -75.22 20.09 -75.02 ;
        RECT 19.89 -75.82 20.09 -75.62 ;
        RECT 19.89 -76.42 20.09 -76.22 ;
        RECT 19.89 -77.02 20.09 -76.82 ;
        RECT 19.89 -77.62 20.09 -77.42 ;
        RECT 19.89 -78.22 20.09 -78.02 ;
        RECT 20.19 -68.87 20.39 -68.67 ;
        RECT 20.19 -69.47 20.39 -69.27 ;
        RECT 20.19 -70.07 20.39 -69.87 ;
        RECT 20.19 -70.67 20.39 -70.47 ;
        RECT 20.37 -71.92 20.57 -71.72 ;
        RECT 20.37 -72.52 20.57 -72.32 ;
        RECT 20.37 -73.12 20.57 -72.92 ;
        RECT 20.37 -73.72 20.57 -73.52 ;
        RECT 20.37 -74.32 20.57 -74.12 ;
        RECT 20.37 -74.92 20.57 -74.72 ;
        RECT 20.37 -75.52 20.57 -75.32 ;
        RECT 20.37 -76.12 20.57 -75.92 ;
        RECT 20.37 -76.72 20.57 -76.52 ;
        RECT 20.37 -77.32 20.57 -77.12 ;
        RECT 20.37 -77.92 20.57 -77.72 ;
        RECT 20.37 -78.52 20.57 -78.32 ;
        RECT 20.79 -68.87 20.99 -68.67 ;
        RECT 20.79 -69.47 20.99 -69.27 ;
        RECT 20.79 -70.07 20.99 -69.87 ;
        RECT 20.79 -70.67 20.99 -70.47 ;
        RECT 20.85 -71.62 21.05 -71.42 ;
        RECT 20.85 -72.22 21.05 -72.02 ;
        RECT 20.85 -72.82 21.05 -72.62 ;
        RECT 20.85 -73.42 21.05 -73.22 ;
        RECT 20.85 -74.02 21.05 -73.82 ;
        RECT 20.85 -74.62 21.05 -74.42 ;
        RECT 20.85 -75.22 21.05 -75.02 ;
        RECT 20.85 -75.82 21.05 -75.62 ;
        RECT 20.85 -76.42 21.05 -76.22 ;
        RECT 20.85 -77.02 21.05 -76.82 ;
        RECT 20.85 -77.62 21.05 -77.42 ;
        RECT 20.85 -78.22 21.05 -78.02 ;
        RECT 21.33 -71.92 21.53 -71.72 ;
        RECT 21.33 -72.52 21.53 -72.32 ;
        RECT 21.33 -73.12 21.53 -72.92 ;
        RECT 21.33 -73.72 21.53 -73.52 ;
        RECT 21.33 -74.32 21.53 -74.12 ;
        RECT 21.33 -74.92 21.53 -74.72 ;
        RECT 21.33 -75.52 21.53 -75.32 ;
        RECT 21.33 -76.12 21.53 -75.92 ;
        RECT 21.33 -76.72 21.53 -76.52 ;
        RECT 21.33 -77.32 21.53 -77.12 ;
        RECT 21.33 -77.92 21.53 -77.72 ;
        RECT 21.33 -78.52 21.53 -78.32 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER M3 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER M4 ;
        RECT 11.21 -93.67 21.57 -83.33 ;
      LAYER V3 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
      LAYER V1 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
      LAYER V2 ;
        RECT 11.25 -83.62 11.45 -83.42 ;
        RECT 11.25 -84.22 11.45 -84.02 ;
        RECT 11.25 -84.82 11.45 -84.62 ;
        RECT 11.25 -85.42 11.45 -85.22 ;
        RECT 11.25 -86.02 11.45 -85.82 ;
        RECT 11.25 -86.62 11.45 -86.42 ;
        RECT 11.25 -87.22 11.45 -87.02 ;
        RECT 11.25 -87.82 11.45 -87.62 ;
        RECT 11.25 -88.42 11.45 -88.22 ;
        RECT 11.25 -89.02 11.45 -88.82 ;
        RECT 11.25 -89.62 11.45 -89.42 ;
        RECT 11.25 -90.22 11.45 -90.02 ;
        RECT 11.73 -83.92 11.93 -83.72 ;
        RECT 11.73 -84.52 11.93 -84.32 ;
        RECT 11.73 -85.12 11.93 -84.92 ;
        RECT 11.73 -85.72 11.93 -85.52 ;
        RECT 11.73 -86.32 11.93 -86.12 ;
        RECT 11.73 -86.92 11.93 -86.72 ;
        RECT 11.73 -87.52 11.93 -87.32 ;
        RECT 11.73 -88.12 11.93 -87.92 ;
        RECT 11.73 -88.72 11.93 -88.52 ;
        RECT 11.73 -89.32 11.93 -89.12 ;
        RECT 11.73 -89.92 11.93 -89.72 ;
        RECT 11.73 -90.52 11.93 -90.32 ;
        RECT 11.79 -91.47 11.99 -91.27 ;
        RECT 11.79 -92.07 11.99 -91.87 ;
        RECT 11.79 -92.67 11.99 -92.47 ;
        RECT 11.79 -93.27 11.99 -93.07 ;
        RECT 12.21 -83.62 12.41 -83.42 ;
        RECT 12.21 -84.22 12.41 -84.02 ;
        RECT 12.21 -84.82 12.41 -84.62 ;
        RECT 12.21 -85.42 12.41 -85.22 ;
        RECT 12.21 -86.02 12.41 -85.82 ;
        RECT 12.21 -86.62 12.41 -86.42 ;
        RECT 12.21 -87.22 12.41 -87.02 ;
        RECT 12.21 -87.82 12.41 -87.62 ;
        RECT 12.21 -88.42 12.41 -88.22 ;
        RECT 12.21 -89.02 12.41 -88.82 ;
        RECT 12.21 -89.62 12.41 -89.42 ;
        RECT 12.21 -90.22 12.41 -90.02 ;
        RECT 12.39 -91.47 12.59 -91.27 ;
        RECT 12.39 -92.07 12.59 -91.87 ;
        RECT 12.39 -92.67 12.59 -92.47 ;
        RECT 12.39 -93.27 12.59 -93.07 ;
        RECT 12.69 -83.92 12.89 -83.72 ;
        RECT 12.69 -84.52 12.89 -84.32 ;
        RECT 12.69 -85.12 12.89 -84.92 ;
        RECT 12.69 -85.72 12.89 -85.52 ;
        RECT 12.69 -86.32 12.89 -86.12 ;
        RECT 12.69 -86.92 12.89 -86.72 ;
        RECT 12.69 -87.52 12.89 -87.32 ;
        RECT 12.69 -88.12 12.89 -87.92 ;
        RECT 12.69 -88.72 12.89 -88.52 ;
        RECT 12.69 -89.32 12.89 -89.12 ;
        RECT 12.69 -89.92 12.89 -89.72 ;
        RECT 12.69 -90.52 12.89 -90.32 ;
        RECT 12.99 -91.47 13.19 -91.27 ;
        RECT 12.99 -92.07 13.19 -91.87 ;
        RECT 12.99 -92.67 13.19 -92.47 ;
        RECT 12.99 -93.27 13.19 -93.07 ;
        RECT 13.17 -83.62 13.37 -83.42 ;
        RECT 13.17 -84.22 13.37 -84.02 ;
        RECT 13.17 -84.82 13.37 -84.62 ;
        RECT 13.17 -85.42 13.37 -85.22 ;
        RECT 13.17 -86.02 13.37 -85.82 ;
        RECT 13.17 -86.62 13.37 -86.42 ;
        RECT 13.17 -87.22 13.37 -87.02 ;
        RECT 13.17 -87.82 13.37 -87.62 ;
        RECT 13.17 -88.42 13.37 -88.22 ;
        RECT 13.17 -89.02 13.37 -88.82 ;
        RECT 13.17 -89.62 13.37 -89.42 ;
        RECT 13.17 -90.22 13.37 -90.02 ;
        RECT 13.59 -91.47 13.79 -91.27 ;
        RECT 13.59 -92.07 13.79 -91.87 ;
        RECT 13.59 -92.67 13.79 -92.47 ;
        RECT 13.59 -93.27 13.79 -93.07 ;
        RECT 13.65 -83.92 13.85 -83.72 ;
        RECT 13.65 -84.52 13.85 -84.32 ;
        RECT 13.65 -85.12 13.85 -84.92 ;
        RECT 13.65 -85.72 13.85 -85.52 ;
        RECT 13.65 -86.32 13.85 -86.12 ;
        RECT 13.65 -86.92 13.85 -86.72 ;
        RECT 13.65 -87.52 13.85 -87.32 ;
        RECT 13.65 -88.12 13.85 -87.92 ;
        RECT 13.65 -88.72 13.85 -88.52 ;
        RECT 13.65 -89.32 13.85 -89.12 ;
        RECT 13.65 -89.92 13.85 -89.72 ;
        RECT 13.65 -90.52 13.85 -90.32 ;
        RECT 14.13 -83.62 14.33 -83.42 ;
        RECT 14.13 -84.22 14.33 -84.02 ;
        RECT 14.13 -84.82 14.33 -84.62 ;
        RECT 14.13 -85.42 14.33 -85.22 ;
        RECT 14.13 -86.02 14.33 -85.82 ;
        RECT 14.13 -86.62 14.33 -86.42 ;
        RECT 14.13 -87.22 14.33 -87.02 ;
        RECT 14.13 -87.82 14.33 -87.62 ;
        RECT 14.13 -88.42 14.33 -88.22 ;
        RECT 14.13 -89.02 14.33 -88.82 ;
        RECT 14.13 -89.62 14.33 -89.42 ;
        RECT 14.13 -90.22 14.33 -90.02 ;
        RECT 14.19 -91.47 14.39 -91.27 ;
        RECT 14.19 -92.07 14.39 -91.87 ;
        RECT 14.19 -92.67 14.39 -92.47 ;
        RECT 14.19 -93.27 14.39 -93.07 ;
        RECT 14.61 -83.92 14.81 -83.72 ;
        RECT 14.61 -84.52 14.81 -84.32 ;
        RECT 14.61 -85.12 14.81 -84.92 ;
        RECT 14.61 -85.72 14.81 -85.52 ;
        RECT 14.61 -86.32 14.81 -86.12 ;
        RECT 14.61 -86.92 14.81 -86.72 ;
        RECT 14.61 -87.52 14.81 -87.32 ;
        RECT 14.61 -88.12 14.81 -87.92 ;
        RECT 14.61 -88.72 14.81 -88.52 ;
        RECT 14.61 -89.32 14.81 -89.12 ;
        RECT 14.61 -89.92 14.81 -89.72 ;
        RECT 14.61 -90.52 14.81 -90.32 ;
        RECT 14.79 -91.47 14.99 -91.27 ;
        RECT 14.79 -92.07 14.99 -91.87 ;
        RECT 14.79 -92.67 14.99 -92.47 ;
        RECT 14.79 -93.27 14.99 -93.07 ;
        RECT 15.09 -83.62 15.29 -83.42 ;
        RECT 15.09 -84.22 15.29 -84.02 ;
        RECT 15.09 -84.82 15.29 -84.62 ;
        RECT 15.09 -85.42 15.29 -85.22 ;
        RECT 15.09 -86.02 15.29 -85.82 ;
        RECT 15.09 -86.62 15.29 -86.42 ;
        RECT 15.09 -87.22 15.29 -87.02 ;
        RECT 15.09 -87.82 15.29 -87.62 ;
        RECT 15.09 -88.42 15.29 -88.22 ;
        RECT 15.09 -89.02 15.29 -88.82 ;
        RECT 15.09 -89.62 15.29 -89.42 ;
        RECT 15.09 -90.22 15.29 -90.02 ;
        RECT 15.39 -91.47 15.59 -91.27 ;
        RECT 15.39 -92.07 15.59 -91.87 ;
        RECT 15.39 -92.67 15.59 -92.47 ;
        RECT 15.39 -93.27 15.59 -93.07 ;
        RECT 15.57 -83.92 15.77 -83.72 ;
        RECT 15.57 -84.52 15.77 -84.32 ;
        RECT 15.57 -85.12 15.77 -84.92 ;
        RECT 15.57 -85.72 15.77 -85.52 ;
        RECT 15.57 -86.32 15.77 -86.12 ;
        RECT 15.57 -86.92 15.77 -86.72 ;
        RECT 15.57 -87.52 15.77 -87.32 ;
        RECT 15.57 -88.12 15.77 -87.92 ;
        RECT 15.57 -88.72 15.77 -88.52 ;
        RECT 15.57 -89.32 15.77 -89.12 ;
        RECT 15.57 -89.92 15.77 -89.72 ;
        RECT 15.57 -90.52 15.77 -90.32 ;
        RECT 15.99 -91.47 16.19 -91.27 ;
        RECT 15.99 -92.07 16.19 -91.87 ;
        RECT 15.99 -92.67 16.19 -92.47 ;
        RECT 15.99 -93.27 16.19 -93.07 ;
        RECT 16.05 -83.62 16.25 -83.42 ;
        RECT 16.05 -84.22 16.25 -84.02 ;
        RECT 16.05 -84.82 16.25 -84.62 ;
        RECT 16.05 -85.42 16.25 -85.22 ;
        RECT 16.05 -86.02 16.25 -85.82 ;
        RECT 16.05 -86.62 16.25 -86.42 ;
        RECT 16.05 -87.22 16.25 -87.02 ;
        RECT 16.05 -87.82 16.25 -87.62 ;
        RECT 16.05 -88.42 16.25 -88.22 ;
        RECT 16.05 -89.02 16.25 -88.82 ;
        RECT 16.05 -89.62 16.25 -89.42 ;
        RECT 16.05 -90.22 16.25 -90.02 ;
        RECT 16.53 -83.92 16.73 -83.72 ;
        RECT 16.53 -84.52 16.73 -84.32 ;
        RECT 16.53 -85.12 16.73 -84.92 ;
        RECT 16.53 -85.72 16.73 -85.52 ;
        RECT 16.53 -86.32 16.73 -86.12 ;
        RECT 16.53 -86.92 16.73 -86.72 ;
        RECT 16.53 -87.52 16.73 -87.32 ;
        RECT 16.53 -88.12 16.73 -87.92 ;
        RECT 16.53 -88.72 16.73 -88.52 ;
        RECT 16.53 -89.32 16.73 -89.12 ;
        RECT 16.53 -89.92 16.73 -89.72 ;
        RECT 16.53 -90.52 16.73 -90.32 ;
        RECT 16.59 -91.47 16.79 -91.27 ;
        RECT 16.59 -92.07 16.79 -91.87 ;
        RECT 16.59 -92.67 16.79 -92.47 ;
        RECT 16.59 -93.27 16.79 -93.07 ;
        RECT 17.01 -83.62 17.21 -83.42 ;
        RECT 17.01 -84.22 17.21 -84.02 ;
        RECT 17.01 -84.82 17.21 -84.62 ;
        RECT 17.01 -85.42 17.21 -85.22 ;
        RECT 17.01 -86.02 17.21 -85.82 ;
        RECT 17.01 -86.62 17.21 -86.42 ;
        RECT 17.01 -87.22 17.21 -87.02 ;
        RECT 17.01 -87.82 17.21 -87.62 ;
        RECT 17.01 -88.42 17.21 -88.22 ;
        RECT 17.01 -89.02 17.21 -88.82 ;
        RECT 17.01 -89.62 17.21 -89.42 ;
        RECT 17.01 -90.22 17.21 -90.02 ;
        RECT 17.19 -91.47 17.39 -91.27 ;
        RECT 17.19 -92.07 17.39 -91.87 ;
        RECT 17.19 -92.67 17.39 -92.47 ;
        RECT 17.19 -93.27 17.39 -93.07 ;
        RECT 17.49 -83.92 17.69 -83.72 ;
        RECT 17.49 -84.52 17.69 -84.32 ;
        RECT 17.49 -85.12 17.69 -84.92 ;
        RECT 17.49 -85.72 17.69 -85.52 ;
        RECT 17.49 -86.32 17.69 -86.12 ;
        RECT 17.49 -86.92 17.69 -86.72 ;
        RECT 17.49 -87.52 17.69 -87.32 ;
        RECT 17.49 -88.12 17.69 -87.92 ;
        RECT 17.49 -88.72 17.69 -88.52 ;
        RECT 17.49 -89.32 17.69 -89.12 ;
        RECT 17.49 -89.92 17.69 -89.72 ;
        RECT 17.49 -90.52 17.69 -90.32 ;
        RECT 17.79 -91.47 17.99 -91.27 ;
        RECT 17.79 -92.07 17.99 -91.87 ;
        RECT 17.79 -92.67 17.99 -92.47 ;
        RECT 17.79 -93.27 17.99 -93.07 ;
        RECT 17.97 -83.62 18.17 -83.42 ;
        RECT 17.97 -84.22 18.17 -84.02 ;
        RECT 17.97 -84.82 18.17 -84.62 ;
        RECT 17.97 -85.42 18.17 -85.22 ;
        RECT 17.97 -86.02 18.17 -85.82 ;
        RECT 17.97 -86.62 18.17 -86.42 ;
        RECT 17.97 -87.22 18.17 -87.02 ;
        RECT 17.97 -87.82 18.17 -87.62 ;
        RECT 17.97 -88.42 18.17 -88.22 ;
        RECT 17.97 -89.02 18.17 -88.82 ;
        RECT 17.97 -89.62 18.17 -89.42 ;
        RECT 17.97 -90.22 18.17 -90.02 ;
        RECT 18.39 -91.47 18.59 -91.27 ;
        RECT 18.39 -92.07 18.59 -91.87 ;
        RECT 18.39 -92.67 18.59 -92.47 ;
        RECT 18.39 -93.27 18.59 -93.07 ;
        RECT 18.45 -83.92 18.65 -83.72 ;
        RECT 18.45 -84.52 18.65 -84.32 ;
        RECT 18.45 -85.12 18.65 -84.92 ;
        RECT 18.45 -85.72 18.65 -85.52 ;
        RECT 18.45 -86.32 18.65 -86.12 ;
        RECT 18.45 -86.92 18.65 -86.72 ;
        RECT 18.45 -87.52 18.65 -87.32 ;
        RECT 18.45 -88.12 18.65 -87.92 ;
        RECT 18.45 -88.72 18.65 -88.52 ;
        RECT 18.45 -89.32 18.65 -89.12 ;
        RECT 18.45 -89.92 18.65 -89.72 ;
        RECT 18.45 -90.52 18.65 -90.32 ;
        RECT 18.93 -83.62 19.13 -83.42 ;
        RECT 18.93 -84.22 19.13 -84.02 ;
        RECT 18.93 -84.82 19.13 -84.62 ;
        RECT 18.93 -85.42 19.13 -85.22 ;
        RECT 18.93 -86.02 19.13 -85.82 ;
        RECT 18.93 -86.62 19.13 -86.42 ;
        RECT 18.93 -87.22 19.13 -87.02 ;
        RECT 18.93 -87.82 19.13 -87.62 ;
        RECT 18.93 -88.42 19.13 -88.22 ;
        RECT 18.93 -89.02 19.13 -88.82 ;
        RECT 18.93 -89.62 19.13 -89.42 ;
        RECT 18.93 -90.22 19.13 -90.02 ;
        RECT 18.99 -91.47 19.19 -91.27 ;
        RECT 18.99 -92.07 19.19 -91.87 ;
        RECT 18.99 -92.67 19.19 -92.47 ;
        RECT 18.99 -93.27 19.19 -93.07 ;
        RECT 19.41 -83.92 19.61 -83.72 ;
        RECT 19.41 -84.52 19.61 -84.32 ;
        RECT 19.41 -85.12 19.61 -84.92 ;
        RECT 19.41 -85.72 19.61 -85.52 ;
        RECT 19.41 -86.32 19.61 -86.12 ;
        RECT 19.41 -86.92 19.61 -86.72 ;
        RECT 19.41 -87.52 19.61 -87.32 ;
        RECT 19.41 -88.12 19.61 -87.92 ;
        RECT 19.41 -88.72 19.61 -88.52 ;
        RECT 19.41 -89.32 19.61 -89.12 ;
        RECT 19.41 -89.92 19.61 -89.72 ;
        RECT 19.41 -90.52 19.61 -90.32 ;
        RECT 19.59 -91.47 19.79 -91.27 ;
        RECT 19.59 -92.07 19.79 -91.87 ;
        RECT 19.59 -92.67 19.79 -92.47 ;
        RECT 19.59 -93.27 19.79 -93.07 ;
        RECT 19.89 -83.62 20.09 -83.42 ;
        RECT 19.89 -84.22 20.09 -84.02 ;
        RECT 19.89 -84.82 20.09 -84.62 ;
        RECT 19.89 -85.42 20.09 -85.22 ;
        RECT 19.89 -86.02 20.09 -85.82 ;
        RECT 19.89 -86.62 20.09 -86.42 ;
        RECT 19.89 -87.22 20.09 -87.02 ;
        RECT 19.89 -87.82 20.09 -87.62 ;
        RECT 19.89 -88.42 20.09 -88.22 ;
        RECT 19.89 -89.02 20.09 -88.82 ;
        RECT 19.89 -89.62 20.09 -89.42 ;
        RECT 19.89 -90.22 20.09 -90.02 ;
        RECT 20.19 -91.47 20.39 -91.27 ;
        RECT 20.19 -92.07 20.39 -91.87 ;
        RECT 20.19 -92.67 20.39 -92.47 ;
        RECT 20.19 -93.27 20.39 -93.07 ;
        RECT 20.37 -83.92 20.57 -83.72 ;
        RECT 20.37 -84.52 20.57 -84.32 ;
        RECT 20.37 -85.12 20.57 -84.92 ;
        RECT 20.37 -85.72 20.57 -85.52 ;
        RECT 20.37 -86.32 20.57 -86.12 ;
        RECT 20.37 -86.92 20.57 -86.72 ;
        RECT 20.37 -87.52 20.57 -87.32 ;
        RECT 20.37 -88.12 20.57 -87.92 ;
        RECT 20.37 -88.72 20.57 -88.52 ;
        RECT 20.37 -89.32 20.57 -89.12 ;
        RECT 20.37 -89.92 20.57 -89.72 ;
        RECT 20.37 -90.52 20.57 -90.32 ;
        RECT 20.79 -91.47 20.99 -91.27 ;
        RECT 20.79 -92.07 20.99 -91.87 ;
        RECT 20.79 -92.67 20.99 -92.47 ;
        RECT 20.79 -93.27 20.99 -93.07 ;
        RECT 20.85 -83.62 21.05 -83.42 ;
        RECT 20.85 -84.22 21.05 -84.02 ;
        RECT 20.85 -84.82 21.05 -84.62 ;
        RECT 20.85 -85.42 21.05 -85.22 ;
        RECT 20.85 -86.02 21.05 -85.82 ;
        RECT 20.85 -86.62 21.05 -86.42 ;
        RECT 20.85 -87.22 21.05 -87.02 ;
        RECT 20.85 -87.82 21.05 -87.62 ;
        RECT 20.85 -88.42 21.05 -88.22 ;
        RECT 20.85 -89.02 21.05 -88.82 ;
        RECT 20.85 -89.62 21.05 -89.42 ;
        RECT 20.85 -90.22 21.05 -90.02 ;
        RECT 21.33 -83.92 21.53 -83.72 ;
        RECT 21.33 -84.52 21.53 -84.32 ;
        RECT 21.33 -85.12 21.53 -84.92 ;
        RECT 21.33 -85.72 21.53 -85.52 ;
        RECT 21.33 -86.32 21.53 -86.12 ;
        RECT 21.33 -86.92 21.53 -86.72 ;
        RECT 21.33 -87.52 21.53 -87.32 ;
        RECT 21.33 -88.12 21.53 -87.92 ;
        RECT 21.33 -88.72 21.53 -88.52 ;
        RECT 21.33 -89.32 21.53 -89.12 ;
        RECT 21.33 -89.92 21.53 -89.72 ;
        RECT 21.33 -90.52 21.53 -90.32 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.93 -69.17 22.93 -68.17 ;
      LAYER M3 ;
        RECT 21.93 -69.17 22.93 -68.17 ;
      LAYER V3 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
      LAYER V1 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
      LAYER V2 ;
        RECT 21.93 -68.37 22.13 -68.17 ;
        RECT 21.93 -68.77 22.13 -68.57 ;
        RECT 21.93 -69.17 22.13 -68.97 ;
        RECT 22.33 -68.37 22.53 -68.17 ;
        RECT 22.33 -68.77 22.53 -68.57 ;
        RECT 22.33 -69.17 22.53 -68.97 ;
        RECT 22.73 -68.37 22.93 -68.17 ;
        RECT 22.73 -68.77 22.93 -68.57 ;
        RECT 22.73 -69.17 22.93 -68.97 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.28 -53.12 27.88 -52.54 ;
      LAYER V1 ;
        RECT 27.28 -52.74 27.48 -52.54 ;
        RECT 27.28 -53.14 27.48 -52.94 ;
        RECT 27.68 -52.74 27.88 -52.54 ;
        RECT 27.68 -53.14 27.88 -52.94 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.22 -90.74 38.82 -90.14 ;
      LAYER M3 ;
        RECT 38.22 -90.74 38.82 -90.52 ;
        RECT 38.52 -90.8 38.82 -90.52 ;
      LAYER V1 ;
        RECT 38.22 -90.34 38.42 -90.14 ;
        RECT 38.22 -90.74 38.42 -90.54 ;
        RECT 38.62 -90.34 38.82 -90.14 ;
        RECT 38.62 -90.74 38.82 -90.54 ;
      LAYER V2 ;
        RECT 38.22 -90.34 38.42 -90.14 ;
        RECT 38.22 -90.74 38.42 -90.54 ;
        RECT 38.62 -90.34 38.82 -90.14 ;
        RECT 38.62 -90.74 38.82 -90.54 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.16 -92.22 3.4 -91.98 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.01 -68.27 4.15 -68.11 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.72 -63.63 9.98 -63.39 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.16 -59.29 24.44 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.12 -59.29 25.4 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.08 -59.29 26.36 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.56 -59.29 26.84 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.52 -59.29 27.8 -59.03 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.82 -77.96 59.94 -76.84 ;
      LAYER M2 ;
        RECT 58.88 -77.9 59.88 -76.9 ;
      LAYER M3 ;
        RECT 58.88 -77.9 59.88 -76.9 ;
      LAYER M4 ;
        RECT 58.88 -77.9 59.88 -76.92 ;
      LAYER V3 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
      LAYER V1 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
      LAYER V2 ;
        RECT 58.88 -77.1 59.08 -76.9 ;
        RECT 58.88 -77.5 59.08 -77.3 ;
        RECT 58.88 -77.9 59.08 -77.7 ;
        RECT 59.28 -77.1 59.48 -76.9 ;
        RECT 59.28 -77.5 59.48 -77.3 ;
        RECT 59.28 -77.9 59.48 -77.7 ;
        RECT 59.68 -77.1 59.88 -76.9 ;
        RECT 59.68 -77.5 59.88 -77.3 ;
        RECT 59.68 -77.9 59.88 -77.7 ;
    END
  END AVSS
  OBS
    LAYER M1 ;
      RECT 66.12 -69.65 124.78 -68.77 ;
      RECT 124.34 -90.25 124.78 -68.77 ;
      RECT 66.82 -70.61 124 -70.03 ;
      RECT 123.38 -88.79 124 -70.03 ;
      RECT 64.32 -88.85 64.72 -72.53 ;
      RECT 59.93 -80.36 62.62 -78.73 ;
      RECT 61.84 -82.73 62.62 -78.73 ;
      RECT 61.84 -82.33 64.72 -79.13 ;
      RECT 57.35 -82.58 57.51 -78.63 ;
      RECT 54.45 -82.58 54.61 -78.63 ;
      RECT 51.55 -82.58 51.71 -78.63 ;
      RECT 48.65 -82.58 48.81 -78.63 ;
      RECT 45.75 -82.58 45.91 -78.63 ;
      RECT 45.07 -82.58 57.55 -82.28 ;
      RECT 56.85 -83.83 57.01 -82.28 ;
      RECT 54.15 -83.83 54.31 -82.28 ;
      RECT 51.45 -83.83 51.61 -82.28 ;
      RECT 48.75 -83.83 48.91 -82.28 ;
      RECT 46.05 -83.83 46.21 -82.28 ;
      RECT -0.34 -52.94 51.16 -50.94 ;
      RECT 23.98 -52.99 51.15 -50.94 ;
      RECT 50.75 -62.45 51.15 -50.94 ;
      RECT -0.34 -96.32 1.66 -50.94 ;
      RECT 23.98 -53.28 32.38 -50.94 ;
      RECT 27.63 -54.25 27.79 -50.94 ;
      RECT 26.57 -54.25 26.73 -50.94 ;
      RECT 26.2 -54.25 26.36 -50.94 ;
      RECT 25.13 -54.25 25.29 -50.94 ;
      RECT 24.16 -54.25 24.32 -50.94 ;
      RECT 27.52 -54.25 27.8 -53.96 ;
      RECT 26.56 -54.25 26.84 -53.96 ;
      RECT 26.08 -54.25 26.36 -53.96 ;
      RECT 25.12 -54.25 25.4 -53.96 ;
      RECT 24.16 -54.25 24.44 -53.96 ;
      RECT 50.03 -62.45 51.15 -62.05 ;
      RECT 9.72 -66.39 9.98 -65.55 ;
      RECT 9.82 -69.75 9.98 -65.55 ;
      RECT 9.72 -69.75 9.98 -67.87 ;
      RECT 6.07 -68.27 22.99 -68.11 ;
      RECT 21.87 -69.23 22.99 -68.11 ;
      RECT 11.21 -93.67 21.57 -68.11 ;
      RECT 45.6 -92.77 45.76 -86.99 ;
      RECT 43.15 -92.77 43.31 -86.99 ;
      RECT 38.61 -92.77 38.77 -87 ;
      RECT 36.16 -92.77 36.32 -87 ;
      RECT 45.54 -87.45 45.76 -87.05 ;
      RECT 45.54 -88.87 45.76 -88.47 ;
      RECT 45.54 -92.77 45.76 -89.91 ;
      RECT 38.16 -92.77 38.88 -90.08 ;
      RECT 45.53 -92.77 45.83 -90.12 ;
      RECT 43.08 -92.77 43.38 -90.21 ;
      RECT 36.09 -92.77 36.39 -90.21 ;
      RECT 36.09 -92.77 43.38 -90.52 ;
      RECT 36.09 -92.77 45.83 -90.58 ;
      RECT 33.94 -92.77 46.82 -90.77 ;
      RECT 33.94 -96.32 35.94 -90.77 ;
      RECT 14.61 -96.32 14.85 -68.11 ;
      RECT 11.22 -96.32 11.46 -68.11 ;
      RECT 5.32 -96.32 14.85 -94.13 ;
      RECT 3.16 -96.32 14.85 -94.14 ;
      RECT -0.34 -96.32 35.94 -94.32 ;
      RECT 66.12 -92.61 122.42 -91.73 ;
      RECT 66.8 -91.33 121.46 -90.77 ;
      RECT 42.85 -80.36 43.01 -78.63 ;
      RECT 5.32 -93.03 9.21 -92.87 ;
    LAYER M1 SPACING 0.16 ;
      RECT -0.34 -53.46 125.11 -50.4 ;
      RECT 124.32 -91.85 125.11 -50.4 ;
      RECT 35.06 -67.71 125.11 -50.4 ;
      RECT 123.3 -90.39 125.11 -50.4 ;
      RECT -0.34 -53.72 34.08 -50.4 ;
      RECT 31.96 -68.63 34.08 -50.4 ;
      RECT 31 -54.29 31.16 -50.4 ;
      RECT 30.04 -54.29 30.2 -50.4 ;
      RECT 29.08 -54.29 29.24 -50.4 ;
      RECT -0.34 -54.03 28.28 -50.4 ;
      RECT 22.2 -54.29 28.28 -50.4 ;
      RECT 31.84 -54.29 34.08 -54 ;
      RECT 30.88 -54.29 31.16 -54 ;
      RECT 29.92 -54.29 30.2 -54 ;
      RECT 28.96 -54.29 29.24 -54 ;
      RECT -0.34 -60.15 20.84 -50.4 ;
      RECT 32.63 -96.4 36.23 -54.27 ;
      RECT 22.2 -54.32 28.16 -50.4 ;
      RECT 24.76 -54.87 28.16 -50.4 ;
      RECT 27.16 -55.12 28.16 -50.4 ;
      RECT 22.2 -54.87 24.12 -50.4 ;
      RECT 31.67 -68.63 36.23 -54.58 ;
      RECT 26.68 -54.98 125.11 -54.58 ;
      RECT 28.12 -67.71 125.11 -54.58 ;
      RECT 25.72 -59.32 25.89 -50.4 ;
      RECT 24.76 -56.08 24.92 -50.4 ;
      RECT 22.2 -56.08 23.84 -50.4 ;
      RECT 27.16 -55.48 27.33 -50.4 ;
      RECT 25.6 -58.71 25.89 -55.19 ;
      RECT 24.64 -56.08 24.92 -55.19 ;
      RECT 27.04 -55.59 27.32 -55.3 ;
      RECT -0.34 -57.74 23.66 -55.39 ;
      RECT 28 -58.71 125.11 -55.49 ;
      RECT -0.34 -56.08 26.36 -55.79 ;
      RECT 24.78 -58.71 125.11 -55.9 ;
      RECT 24.76 -59.32 24.92 -57.2 ;
      RECT 22.97 -58.16 125.11 -57.2 ;
      RECT -0.34 -60.15 21.61 -55.39 ;
      RECT 22.97 -58.71 24.12 -57.2 ;
      RECT 27.16 -59.32 27.33 -55.9 ;
      RECT 22.97 -61.41 23.84 -57.2 ;
      RECT 28 -59.28 125.11 -58.99 ;
      RECT 27.04 -59.32 27.33 -59.03 ;
      RECT 25.6 -59.32 25.89 -59.03 ;
      RECT 24.64 -59.32 24.92 -59.03 ;
      RECT 8.36 -61.41 23.84 -59.1 ;
      RECT 27.16 -62.32 125.11 -59.61 ;
      RECT 4.49 -60.87 125.11 -59.61 ;
      RECT 26.68 -62.18 125.11 -59.61 ;
      RECT -0.34 -91.66 3.69 -50.4 ;
      RECT 24.76 -62.07 125.11 -59.61 ;
      RECT 4.49 -96.4 7 -50.4 ;
      RECT -0.34 -67.79 7 -60.95 ;
      RECT 23.72 -61.52 125.11 -59.61 ;
      RECT 8.36 -63.07 22.36 -59.1 ;
      RECT -0.34 -61.67 7.01 -61.51 ;
      RECT 23.72 -62.07 24.12 -59.61 ;
      RECT 25.72 -68.63 25.89 -59.61 ;
      RECT 24.76 -63.28 24.92 -59.61 ;
      RECT 4.47 -96.4 9.4 -62.23 ;
      RECT 27.16 -62.68 27.33 -59.61 ;
      RECT 25.6 -68.63 25.89 -62.39 ;
      RECT 24.64 -63.28 24.92 -62.39 ;
      RECT 27.04 -62.79 27.32 -62.5 ;
      RECT 28 -68.63 30.73 -62.69 ;
      RECT -0.34 -63.07 23.84 -62.77 ;
      RECT 10.3 -63.28 26.36 -62.99 ;
      RECT 24.78 -68.63 26.36 -62.99 ;
      RECT 26.25 -96.4 28.01 -63.1 ;
      RECT 10.3 -96.4 23.66 -62.77 ;
      RECT -0.34 -67.79 23.66 -63.95 ;
      RECT 4.47 -96.4 25.35 -64.4 ;
      RECT 37.19 -68.21 125.11 -50.4 ;
      RECT 122.72 -90.05 125.11 -50.4 ;
      RECT 47.36 -68.45 125.11 -50.4 ;
      RECT 65.22 -90.03 125.11 -50.4 ;
      RECT 37.19 -81.96 46.48 -50.4 ;
      RECT 64.52 -69.71 125.11 -50.4 ;
      RECT 47.36 -68.52 63 -50.4 ;
      RECT 32.63 -96.4 36.38 -68.52 ;
      RECT 51.95 -68.72 63 -50.4 ;
      RECT 57.02 -76.52 63 -50.4 ;
      RECT 47.36 -68.72 50.99 -50.4 ;
      RECT 29.12 -96.4 30.73 -54.58 ;
      RECT -0.34 -91.66 25.35 -68.59 ;
      RECT 29.12 -96.4 31.73 -68.65 ;
      RECT 32.63 -81.96 46.48 -68.67 ;
      RECT 54.46 -85.43 56.12 -50.4 ;
      RECT 51.95 -96.4 53.48 -50.4 ;
      RECT 47.36 -69.11 50.87 -50.4 ;
      RECT 32.63 -81.96 47.32 -69.09 ;
      RECT 48.12 -85.43 50.87 -50.4 ;
      RECT 51.77 -85.43 53.48 -69.48 ;
      RECT 29.12 -81.96 47.32 -69.53 ;
      RECT -0.34 -91.66 28.01 -69.53 ;
      RECT 54.46 -76.52 63 -69.62 ;
      RECT 48.12 -85.43 53.48 -69.62 ;
      RECT 48.12 -85.43 58.5 -69.7 ;
      RECT 3.72 -96.4 42.53 -69.74 ;
      RECT 46.53 -96.4 48.43 -69.91 ;
      RECT 60.26 -91.41 64 -69.97 ;
      RECT 65.12 -90.03 125.11 -70.77 ;
      RECT 60.26 -90.05 65.38 -70.93 ;
      RECT -0.34 -81.96 125.11 -78.28 ;
      RECT 60.24 -96.4 63 -78.28 ;
      RECT 43.47 -85.43 59.15 -78.28 ;
      RECT -0.34 -85.43 59.15 -82.9 ;
      RECT 57.33 -96.4 63 -83.05 ;
      RECT 54.63 -96.4 56.53 -69.62 ;
      RECT 51.93 -96.4 53.83 -69.7 ;
      RECT 49.23 -96.4 51.13 -69.62 ;
      RECT 43.83 -96.4 45.73 -50.4 ;
      RECT -0.34 -91.66 43.03 -82.9 ;
      RECT 43.83 -90.03 125.11 -86.18 ;
      RECT 3.72 -96.4 63 -86.23 ;
      RECT 121.76 -90.05 122.02 -50.4 ;
      RECT 120.8 -90.05 121.06 -50.4 ;
      RECT 119.84 -90.05 120.1 -50.4 ;
      RECT 118.88 -90.05 119.14 -50.4 ;
      RECT 117.92 -90.05 118.18 -50.4 ;
      RECT 116.96 -90.05 117.22 -50.4 ;
      RECT 116 -90.05 116.26 -50.4 ;
      RECT 115.04 -90.05 115.3 -50.4 ;
      RECT 114.08 -90.05 114.34 -50.4 ;
      RECT 113.12 -90.05 113.38 -50.4 ;
      RECT 112.16 -90.05 112.42 -50.4 ;
      RECT 111.2 -90.05 111.46 -50.4 ;
      RECT 110.24 -90.05 110.5 -50.4 ;
      RECT 109.28 -90.05 109.54 -50.4 ;
      RECT 108.32 -90.05 108.58 -50.4 ;
      RECT 107.36 -90.05 107.62 -50.4 ;
      RECT 106.4 -90.05 106.66 -50.4 ;
      RECT 105.44 -90.05 105.7 -50.4 ;
      RECT 104.48 -90.05 104.74 -50.4 ;
      RECT 103.52 -90.05 103.78 -50.4 ;
      RECT 102.56 -90.05 102.82 -50.4 ;
      RECT 101.6 -90.05 101.86 -50.4 ;
      RECT 100.64 -90.05 100.9 -50.4 ;
      RECT 99.68 -90.05 99.94 -50.4 ;
      RECT 98.72 -90.05 98.98 -50.4 ;
      RECT 97.76 -90.05 98.02 -50.4 ;
      RECT 96.8 -90.05 97.06 -50.4 ;
      RECT 95.84 -90.05 96.1 -50.4 ;
      RECT 94.88 -90.05 95.14 -50.4 ;
      RECT 93.92 -90.05 94.18 -50.4 ;
      RECT 92.96 -90.05 93.22 -50.4 ;
      RECT 92 -90.05 92.26 -50.4 ;
      RECT 91.04 -90.05 91.3 -50.4 ;
      RECT 90.08 -90.05 90.34 -50.4 ;
      RECT 89.12 -90.05 89.38 -50.4 ;
      RECT 88.16 -90.05 88.42 -50.4 ;
      RECT 87.2 -90.05 87.46 -50.4 ;
      RECT 86.24 -90.05 86.5 -50.4 ;
      RECT 85.28 -90.05 85.54 -50.4 ;
      RECT 84.32 -90.05 84.58 -50.4 ;
      RECT 83.36 -90.05 83.62 -50.4 ;
      RECT 82.4 -90.05 82.66 -50.4 ;
      RECT 81.44 -90.05 81.7 -50.4 ;
      RECT 80.48 -90.05 80.74 -50.4 ;
      RECT 79.52 -90.05 79.78 -50.4 ;
      RECT 78.56 -90.05 78.82 -50.4 ;
      RECT 77.6 -90.05 77.86 -50.4 ;
      RECT 76.64 -90.05 76.9 -50.4 ;
      RECT 75.68 -90.05 75.94 -50.4 ;
      RECT 74.72 -90.05 74.98 -50.4 ;
      RECT 73.76 -90.05 74.02 -50.4 ;
      RECT 72.8 -90.05 73.06 -50.4 ;
      RECT 71.84 -90.05 72.1 -50.4 ;
      RECT 70.88 -90.05 71.14 -50.4 ;
      RECT 69.92 -90.05 70.18 -50.4 ;
      RECT 68.96 -90.05 69.22 -50.4 ;
      RECT 68 -90.05 68.26 -50.4 ;
      RECT 67.04 -90.05 67.3 -50.4 ;
      RECT 66.08 -90.05 66.34 -50.4 ;
      RECT -0.34 -90.45 64.8 -86.23 ;
      RECT 65.2 -96.4 123.06 -90.77 ;
      RECT 64.52 -91.85 125.11 -91.65 ;
      RECT -0.34 -96.4 2.84 -50.4 ;
      RECT 64.52 -96.4 124.02 -91.65 ;
      RECT -0.34 -96.4 63 -92.54 ;
      RECT -0.34 -96.4 125.11 -92.93 ;
    LAYER M2 ;
      RECT 122.72 -92.5 122.98 -70.77 ;
      RECT 121.76 -92.5 122.02 -70.77 ;
      RECT 120.8 -92.5 121.06 -70.77 ;
      RECT 119.84 -92.5 120.1 -70.77 ;
      RECT 118.88 -92.5 119.14 -70.77 ;
      RECT 117.92 -92.5 118.18 -70.77 ;
      RECT 116.96 -92.5 117.22 -70.77 ;
      RECT 116 -92.5 116.26 -70.77 ;
      RECT 115.04 -92.5 115.3 -70.77 ;
      RECT 114.08 -92.5 114.34 -70.77 ;
      RECT 113.12 -92.5 113.38 -70.77 ;
      RECT 112.16 -92.5 112.42 -70.77 ;
      RECT 111.2 -92.5 111.46 -70.77 ;
      RECT 110.24 -92.5 110.5 -70.77 ;
      RECT 109.28 -92.5 109.54 -70.77 ;
      RECT 108.32 -92.5 108.58 -70.77 ;
      RECT 107.36 -92.5 107.62 -70.77 ;
      RECT 106.4 -92.5 106.66 -70.77 ;
      RECT 105.44 -92.5 105.7 -70.77 ;
      RECT 104.48 -92.5 104.74 -70.77 ;
      RECT 103.52 -92.5 103.78 -70.77 ;
      RECT 102.56 -92.5 102.82 -70.77 ;
      RECT 101.6 -92.5 101.86 -70.77 ;
      RECT 100.64 -96.35 100.9 -70.77 ;
      RECT 99.68 -96.35 99.94 -70.77 ;
      RECT 98.72 -96.35 98.98 -70.77 ;
      RECT 97.76 -96.35 98.02 -70.77 ;
      RECT 96.8 -96.35 97.06 -70.77 ;
      RECT 95.84 -96.35 96.1 -70.77 ;
      RECT 94.88 -96.35 95.14 -70.77 ;
      RECT 93.92 -96.35 94.18 -70.77 ;
      RECT 92.96 -96.35 93.22 -70.77 ;
      RECT 92 -96.35 92.26 -70.77 ;
      RECT 91.04 -96.35 91.3 -70.77 ;
      RECT 90.08 -96.35 90.34 -70.77 ;
      RECT 89.12 -96.35 89.38 -70.77 ;
      RECT 88.16 -96.35 88.42 -70.77 ;
      RECT 87.2 -96.35 87.46 -70.77 ;
      RECT 86.24 -92.5 86.5 -70.77 ;
      RECT 85.28 -92.5 85.54 -70.77 ;
      RECT 84.32 -92.5 84.58 -70.77 ;
      RECT 83.36 -92.5 83.62 -70.77 ;
      RECT 82.4 -92.5 82.66 -70.77 ;
      RECT 81.44 -92.5 81.7 -70.77 ;
      RECT 80.48 -92.5 80.74 -70.77 ;
      RECT 79.52 -92.5 79.78 -70.77 ;
      RECT 78.56 -92.5 78.82 -70.77 ;
      RECT 77.6 -92.5 77.86 -70.77 ;
      RECT 76.64 -92.5 76.9 -70.77 ;
      RECT 75.68 -92.5 75.94 -70.77 ;
      RECT 74.72 -92.5 74.98 -70.77 ;
      RECT 73.76 -92.5 74.02 -70.77 ;
      RECT 72.8 -92.5 73.06 -70.77 ;
      RECT 71.84 -92.5 72.1 -70.77 ;
      RECT 70.88 -92.5 71.14 -70.77 ;
      RECT 69.92 -92.5 70.18 -70.77 ;
      RECT 68.96 -92.5 69.22 -70.77 ;
      RECT 68 -92.5 68.26 -70.77 ;
      RECT 67.04 -92.5 67.3 -70.77 ;
      RECT 66.08 -92.5 66.34 -70.77 ;
      RECT 65.12 -92.5 65.38 -70.77 ;
      RECT 65.12 -92.5 122.98 -92.22 ;
      RECT 86.55 -96.35 101.55 -92.22 ;
      RECT 86.55 -69.65 101.55 -67.87 ;
      RECT 63.32 -69.65 121.98 -68.77 ;
      RECT 121.28 -88.43 121.54 -68.77 ;
      RECT 120.32 -88.43 120.58 -68.77 ;
      RECT 119.36 -88.43 119.62 -68.77 ;
      RECT 118.4 -88.43 118.66 -68.77 ;
      RECT 117.44 -88.43 117.7 -68.77 ;
      RECT 116.48 -88.43 116.74 -68.77 ;
      RECT 115.52 -88.43 115.78 -68.77 ;
      RECT 114.56 -88.43 114.82 -68.77 ;
      RECT 113.6 -88.43 113.86 -68.77 ;
      RECT 112.64 -88.43 112.9 -68.77 ;
      RECT 111.68 -88.43 111.94 -68.77 ;
      RECT 110.72 -88.43 110.98 -68.77 ;
      RECT 109.76 -88.43 110.02 -68.77 ;
      RECT 108.8 -88.43 109.06 -68.77 ;
      RECT 107.84 -88.43 108.1 -68.77 ;
      RECT 106.88 -88.43 107.14 -68.77 ;
      RECT 105.92 -88.43 106.18 -68.77 ;
      RECT 104.96 -88.43 105.22 -68.77 ;
      RECT 104 -88.43 104.26 -68.77 ;
      RECT 103.04 -88.43 103.3 -68.77 ;
      RECT 102.08 -88.43 102.34 -68.77 ;
      RECT 101.12 -88.43 101.38 -67.87 ;
      RECT 100.16 -88.43 100.42 -67.87 ;
      RECT 99.2 -88.43 99.46 -67.87 ;
      RECT 98.24 -88.43 98.5 -67.87 ;
      RECT 97.28 -88.43 97.54 -67.87 ;
      RECT 96.32 -88.43 96.58 -67.87 ;
      RECT 95.36 -88.43 95.62 -67.87 ;
      RECT 94.4 -88.43 94.66 -67.87 ;
      RECT 93.44 -88.43 93.7 -67.87 ;
      RECT 92.48 -88.43 92.74 -67.87 ;
      RECT 91.52 -88.43 91.78 -67.87 ;
      RECT 90.56 -88.43 90.82 -67.87 ;
      RECT 89.6 -88.43 89.86 -67.87 ;
      RECT 88.64 -88.43 88.9 -67.87 ;
      RECT 87.68 -88.43 87.94 -67.87 ;
      RECT 86.72 -88.43 86.98 -67.87 ;
      RECT 85.76 -88.43 86.02 -68.77 ;
      RECT 84.8 -88.43 85.06 -68.77 ;
      RECT 83.84 -88.43 84.1 -68.77 ;
      RECT 82.88 -88.43 83.14 -68.77 ;
      RECT 81.92 -88.43 82.18 -68.77 ;
      RECT 80.96 -88.43 81.22 -68.77 ;
      RECT 80 -88.43 80.26 -68.77 ;
      RECT 79.04 -88.43 79.3 -68.77 ;
      RECT 78.08 -88.43 78.34 -68.77 ;
      RECT 77.12 -88.43 77.38 -68.77 ;
      RECT 76.16 -88.43 76.42 -68.77 ;
      RECT 75.2 -88.43 75.46 -68.77 ;
      RECT 74.24 -88.43 74.5 -68.77 ;
      RECT 73.28 -88.43 73.54 -68.77 ;
      RECT 72.32 -88.43 72.58 -68.77 ;
      RECT 71.36 -88.43 71.62 -68.77 ;
      RECT 70.4 -88.43 70.66 -68.77 ;
      RECT 69.44 -88.43 69.7 -68.77 ;
      RECT 68.48 -88.43 68.74 -68.77 ;
      RECT 67.52 -88.43 67.78 -68.77 ;
      RECT 66.56 -88.43 66.82 -68.77 ;
      RECT 65.6 -88.43 65.86 -68.77 ;
      RECT 24.08 -63.94 24.68 -59.06 ;
      RECT 11.3 -61.17 24.68 -59.17 ;
      RECT 20.1 -67.25 22.1 -59.17 ;
      RECT 20.1 -66.11 84.63 -65.25 ;
      RECT 38.35 -67.25 84.63 -65.25 ;
      RECT 20.1 -67.25 34.21 -65.25 ;
      RECT 38.35 -68.33 39.11 -65.25 ;
      RECT 38.35 -68.33 51.61 -68.03 ;
      RECT 51.31 -69.55 51.61 -68.03 ;
      RECT 50.1 -71.66 50.3 -71.06 ;
      RECT 32.99 -71.69 33.19 -71.09 ;
      RECT 32.92 -71.56 50.37 -71.16 ;
      RECT 47.82 -94.08 48.22 -71.16 ;
      RECT 122.24 -88.43 122.5 -71.57 ;
    LAYER M2 SPACING 0.2 ;
      RECT -0.34 -50.65 125.11 -50.4 ;
      RECT 101.85 -68.47 125.11 -50.4 ;
      RECT -0.34 -51.72 86.25 -50.4 ;
      RECT 35.35 -67.73 86.25 -50.4 ;
      RECT -0.34 -52.24 33.75 -50.4 ;
      RECT 28.18 -53.7 33.75 -50.4 ;
      RECT 31.94 -68.65 33.75 -50.4 ;
      RECT -0.34 -54.05 26.98 -50.4 ;
      RECT 35.04 -67.73 86.25 -53.32 ;
      RECT 32.61 -96.4 34.1 -53.32 ;
      RECT 27.14 -62.2 28.18 -53.42 ;
      RECT 22.18 -54.34 28.18 -53.42 ;
      RECT 26.66 -55 28.18 -53.42 ;
      RECT -0.34 -58.87 20.86 -50.4 ;
      RECT 31.94 -67.73 86.25 -54.25 ;
      RECT 24.9 -54.89 28.18 -53.42 ;
      RECT 22.18 -54.89 24.14 -50.4 ;
      RECT 31.65 -68.65 35.83 -54.56 ;
      RECT 28.1 -67.73 86.25 -54.56 ;
      RECT 22.18 -56.1 23.86 -50.4 ;
      RECT -0.34 -57.76 23.68 -55.37 ;
      RECT -0.34 -56.1 26.26 -55.77 ;
      RECT 24.98 -58.73 86.25 -55.88 ;
      RECT 24.76 -56.24 86.25 -55.88 ;
      RECT -0.34 -57.76 23.78 -57.18 ;
      RECT 24.9 -58.73 86.25 -57.44 ;
      RECT 22.95 -58.18 86.25 -57.44 ;
      RECT 10.28 -67.97 21.63 -55.37 ;
      RECT 22.95 -61.43 24.68 -57.44 ;
      RECT 9.68 -63.09 21.63 -55.37 ;
      RECT -0.34 -60.17 7.08 -50.4 ;
      RECT 4.47 -60.89 7.08 -50.4 ;
      RECT 22.95 -61.43 24.82 -58.94 ;
      RECT 9.68 -61.43 24.82 -59.08 ;
      RECT 26.66 -62.2 86.25 -59.59 ;
      RECT -0.34 -91.68 3.71 -50.4 ;
      RECT 4.47 -96.4 7.02 -50.4 ;
      RECT -0.34 -67.81 7.02 -60.93 ;
      RECT 23.7 -61.54 86.25 -59.59 ;
      RECT 24.9 -62.09 86.25 -59.59 ;
      RECT 9.68 -63.09 22.38 -59.08 ;
      RECT 8.34 -63.09 22.38 -61.47 ;
      RECT 23.7 -63.3 24.68 -57.44 ;
      RECT 4.45 -96.4 9.42 -62.21 ;
      RECT 23.7 -63.3 24.82 -62.3 ;
      RECT 10.28 -63.3 24.82 -62.75 ;
      RECT -0.34 -63.09 26.26 -62.97 ;
      RECT 24.76 -68.65 30.75 -63.08 ;
      RECT 24.08 -63.94 86.25 -63.08 ;
      RECT 10.28 -67.87 23.68 -62.75 ;
      RECT 4.45 -96.4 10.91 -63.93 ;
      RECT 23.23 -96.4 25.37 -64.38 ;
      RECT 101.6 -96.4 101.86 -66.25 ;
      RECT 37.11 -68.33 125.11 -66.25 ;
      RECT 65.2 -90.05 123.6 -66.25 ;
      RECT 36.73 -68.33 125.11 -68.03 ;
      RECT 47.34 -68.47 125.11 -66.25 ;
      RECT 64.5 -69.73 86.25 -50.4 ;
      RECT 37.17 -81.98 46.5 -50.4 ;
      RECT 47.34 -68.54 63.02 -50.4 ;
      RECT 51.93 -68.74 63.02 -50.4 ;
      RECT 57 -76.54 63.02 -50.4 ;
      RECT 51.31 -85.45 51.61 -50.4 ;
      RECT 47.34 -68.74 51.01 -50.4 ;
      RECT 3.7 -96.4 10.91 -68.57 ;
      RECT 23.23 -68.65 36.25 -68.63 ;
      RECT 32.61 -96.4 37.92 -68.65 ;
      RECT 29.1 -96.4 31.75 -68.63 ;
      RECT 26.23 -96.4 28.03 -63.08 ;
      RECT 54.44 -85.45 56.14 -50.4 ;
      RECT 51.93 -96.4 53.5 -50.4 ;
      RECT 47.34 -69.13 50.89 -50.4 ;
      RECT 63.32 -69.65 123.6 -68.77 ;
      RECT 48.1 -85.45 50.89 -50.4 ;
      RECT 32.61 -81.98 47.34 -69.07 ;
      RECT 51.31 -85.45 53.5 -69.46 ;
      RECT 21.87 -96.4 25.37 -69.47 ;
      RECT 29.1 -81.98 47.34 -69.51 ;
      RECT 21.87 -96.4 28.03 -69.51 ;
      RECT 54.44 -76.54 63.02 -69.6 ;
      RECT 48.1 -85.45 53.5 -69.6 ;
      RECT 48.1 -85.45 58.52 -69.68 ;
      RECT 21.87 -96.4 37.92 -69.72 ;
      RECT 46.51 -95.7 48.45 -69.89 ;
      RECT 124.3 -91.87 125.11 -69.95 ;
      RECT 60.24 -91.43 64.02 -69.95 ;
      RECT 65.12 -96.4 65.38 -70.77 ;
      RECT 60.24 -90.07 65.38 -70.91 ;
      RECT 21.87 -81.98 125.11 -78.26 ;
      RECT 60.22 -96.4 63.02 -78.26 ;
      RECT -0.34 -83.03 42.55 -78.91 ;
      RECT 43.45 -85.45 59.17 -78.26 ;
      RECT 21.87 -85.45 59.17 -82.88 ;
      RECT 57.31 -96.4 63.02 -83.03 ;
      RECT 54.61 -96.4 56.55 -69.6 ;
      RECT 51.91 -96.4 53.85 -69.68 ;
      RECT 49.21 -96.4 51.15 -69.6 ;
      RECT 43.81 -96.4 45.75 -50.4 ;
      RECT 21.87 -89.84 43.05 -82.88 ;
      RECT 39.12 -95.7 63.02 -86.21 ;
      RECT 122.72 -90.07 125.11 -69.95 ;
      RECT 123.28 -90.41 125.11 -69.95 ;
      RECT 121.76 -96.4 122.02 -50.4 ;
      RECT 120.8 -96.4 121.06 -50.4 ;
      RECT 119.84 -96.4 120.1 -50.4 ;
      RECT 118.88 -96.4 119.14 -50.4 ;
      RECT 117.92 -96.4 118.18 -50.4 ;
      RECT 116.96 -96.4 117.22 -50.4 ;
      RECT 116 -96.4 116.26 -50.4 ;
      RECT 115.04 -96.4 115.3 -50.4 ;
      RECT 114.08 -96.4 114.34 -50.4 ;
      RECT 113.12 -96.4 113.38 -50.4 ;
      RECT 112.16 -96.4 112.42 -50.4 ;
      RECT 111.2 -96.4 111.46 -50.4 ;
      RECT 110.24 -96.4 110.5 -50.4 ;
      RECT 109.28 -96.4 109.54 -50.4 ;
      RECT 108.32 -96.4 108.58 -50.4 ;
      RECT 107.36 -96.4 107.62 -50.4 ;
      RECT 106.4 -96.4 106.66 -50.4 ;
      RECT 105.44 -96.4 105.7 -50.4 ;
      RECT 104.48 -96.4 104.74 -50.4 ;
      RECT 103.52 -96.4 103.78 -50.4 ;
      RECT 102.56 -96.4 102.82 -50.4 ;
      RECT 100.64 -96.4 100.9 -66.25 ;
      RECT 99.68 -96.4 99.94 -66.25 ;
      RECT 98.72 -96.4 98.98 -66.25 ;
      RECT 97.76 -96.4 98.02 -66.25 ;
      RECT 96.8 -96.4 97.06 -66.25 ;
      RECT 95.84 -96.4 96.1 -66.25 ;
      RECT 94.88 -96.4 95.14 -66.25 ;
      RECT 93.92 -96.4 94.18 -66.25 ;
      RECT 92.96 -96.4 93.22 -66.25 ;
      RECT 92 -96.4 92.26 -66.25 ;
      RECT 91.04 -96.4 91.3 -66.25 ;
      RECT 90.08 -96.4 90.34 -66.25 ;
      RECT 89.12 -96.4 89.38 -66.25 ;
      RECT 88.16 -96.4 88.42 -66.25 ;
      RECT 87.2 -96.4 87.46 -66.25 ;
      RECT 86.24 -96.4 86.5 -66.25 ;
      RECT 85.28 -96.4 85.54 -50.4 ;
      RECT 84.32 -96.4 84.58 -50.4 ;
      RECT 83.36 -96.4 83.62 -50.4 ;
      RECT 82.4 -96.4 82.66 -50.4 ;
      RECT 81.44 -96.4 81.7 -50.4 ;
      RECT 80.48 -96.4 80.74 -50.4 ;
      RECT 79.52 -96.4 79.78 -50.4 ;
      RECT 78.56 -96.4 78.82 -50.4 ;
      RECT 77.6 -96.4 77.86 -50.4 ;
      RECT 76.64 -96.4 76.9 -50.4 ;
      RECT 75.68 -96.4 75.94 -50.4 ;
      RECT 74.72 -96.4 74.98 -50.4 ;
      RECT 73.76 -96.4 74.02 -50.4 ;
      RECT 72.8 -96.4 73.06 -50.4 ;
      RECT 71.84 -96.4 72.1 -50.4 ;
      RECT 70.88 -96.4 71.14 -50.4 ;
      RECT 69.92 -96.4 70.18 -50.4 ;
      RECT 68.96 -96.4 69.22 -50.4 ;
      RECT 68 -96.4 68.26 -50.4 ;
      RECT 67.04 -96.4 67.3 -50.4 ;
      RECT 66.08 -96.4 66.34 -50.4 ;
      RECT 122.72 -96.4 122.98 -50.4 ;
      RECT 39.12 -90.47 64.82 -86.21 ;
      RECT 65.12 -96.4 123.08 -90.91 ;
      RECT 21.87 -96.4 47.52 -91.04 ;
      RECT 64.5 -91.87 125.11 -91.63 ;
      RECT -0.34 -96.4 2.86 -50.4 ;
      RECT 64.5 -96.4 124.04 -91.63 ;
      RECT -0.34 -96.4 10.91 -92.52 ;
      RECT 48.52 -96.4 125.11 -92.91 ;
      RECT -0.34 -96.4 47.52 -93.97 ;
      RECT 34.42 -54.02 34.72 -53.3 ;
    LAYER M3 SPACING 0.2 ;
      RECT 11.21 -83.03 21.57 -82.11 ;
      RECT 11.21 -79.83 21.57 -78.91 ;
    LAYER M3 ;
      RECT 34.05 -53.02 56.55 -52.02 ;
      RECT 55.55 -96.34 56.55 -52.02 ;
      RECT 55.55 -96.34 95.61 -95.34 ;
      RECT 38.38 -69 38.98 -68.8 ;
      RECT 38.52 -90.22 38.82 -68.8 ;
      RECT 38.22 -90.22 38.82 -90.14 ;
      RECT 22.94 -62.39 23.14 -50.9 ;
      RECT 22.74 -62.39 23.34 -61.79 ;
      RECT 22.19 -58.72 22.39 -50.9 ;
      RECT 21.99 -58.72 22.59 -58.12 ;
      RECT 21.42 -55.01 21.62 -50.9 ;
      RECT 21.22 -55.01 21.82 -54.41 ;
      RECT 37.76 -53.87 49.99 -53.67 ;
      RECT 11.21 -82.11 21.57 -79.83 ;
    LAYER M4 SPACING 0.2 ;
      RECT 11.21 -83.03 21.57 -82.11 ;
      RECT 11.21 -79.83 21.57 -78.91 ;
    LAYER M4 ;
      RECT 21.93 -69.17 59.88 -68.17 ;
      RECT 58.88 -76.62 59.88 -68.17 ;
      RECT 11.21 -82.11 21.57 -79.83 ;
  END
END LDO_Top_lef

END LIBRARY
