

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO PE_POOL 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8352 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.83812 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0291906 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.143678 LAYER V3 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 1.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0134 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4848 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.5759 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.186427 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.330033 LAYER V3 ;
  END reset
  PIN pe_in_pk_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 84.1667 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.842308 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END pe_in_pk_PE_state__2_
  PIN pe_in_pk_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 3.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.319872 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__1_
  PIN pe_in_pk_PE_state__0_ 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0326 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.5641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.589103 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_PE_state__0_
  PIN pe_in_pk_A__3__7_ 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0358 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.688462 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__7_
  PIN pe_in_pk_A__3__6_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.9103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.496154 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__6_
  PIN pe_in_pk_A__3__5_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.40641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__5_
  PIN pe_in_pk_A__3__4_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.3718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.380769 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__4_
  PIN pe_in_pk_A__3__3_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.355128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__3_
  PIN pe_in_pk_A__3__2_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.2179 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.419231 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__2_
  PIN pe_in_pk_A__3__1_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__1_
  PIN pe_in_pk_A__3__0_ 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0206 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.3462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.470513 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__3__0_
  PIN pe_in_pk_A__2__7_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.432051 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__7_
  PIN pe_in_pk_A__2__6_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__6_
  PIN pe_in_pk_A__2__5_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__5_
  PIN pe_in_pk_A__2__4_ 
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0897 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.367949 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__4_
  PIN pe_in_pk_A__2__3_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.39359 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__3_
  PIN pe_in_pk_A__2__2_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__2_
  PIN pe_in_pk_A__2__1_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.8077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.355128 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__1_
  PIN pe_in_pk_A__2__0_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.3718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.380769 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__2__0_
  PIN pe_in_pk_A__1__7_ 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0142 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.40641 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__7_
  PIN pe_in_pk_A__1__6_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.4103 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.383974 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__1__6_
  PIN pe_in_pk_A__1__5_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.6282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.483333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__5_
  PIN pe_in_pk_A__1__4_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.0641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.457692 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__4_
  PIN pe_in_pk_A__1__3_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.5256 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.342308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__3_
  PIN pe_in_pk_A__1__2_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 56.6026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.573077 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__2_
  PIN pe_in_pk_A__1__1_ 
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0174 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.7564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.534615 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER V3 ;
  END pe_in_pk_A__1__1_
  PIN pe_in_pk_A__1__0_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__1__0_
  PIN pe_in_pk_A__0__7_ 
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.1923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.508974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER V3 ;
  END pe_in_pk_A__0__7_
  PIN pe_in_pk_A__0__6_ 
    ANTENNAPARTIALMETALAREA 1.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.8846 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.342308 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__6_
  PIN pe_in_pk_A__0__5_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0072 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 17.1795 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.191667 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_A__0__5_
  PIN pe_in_pk_A__0__4_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.0897 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.367949 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__4_
  PIN pe_in_pk_A__0__3_ 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0214 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.432051 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__3_
  PIN pe_in_pk_A__0__2_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.329487 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__2_
  PIN pe_in_pk_A__0__1_ 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.6795 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.303846 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__1_
  PIN pe_in_pk_A__0__0_ 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.3462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.470513 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_A__0__0_
  PIN pe_in_pk_wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.1447 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.437736 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER V3 ;
  END pe_in_pk_wrb_data__7_
  PIN pe_in_pk_wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0334 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.6923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.640385 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER V3 ;
  END pe_in_pk_wrb_data__6_
  PIN pe_in_pk_wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 7.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0742 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.6164 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.192453 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.25786 LAYER V3 ;
  END pe_in_pk_wrb_data__5_
  PIN pe_in_pk_wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 6.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0648 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 106.282 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 1.06346 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END pe_in_pk_wrb_data__4_
  PIN pe_in_pk_wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 3.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0342 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 57.2436 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 0.573077 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END pe_in_pk_wrb_data__3_
  PIN pe_in_pk_wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 7.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0776 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 130 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.31987 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_wrb_data__2_
  PIN pe_in_pk_wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 7.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0792 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M4 ; 
    ANTENNAMAXAREACAR 132.564 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.34551 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.20513 LAYER V4 ;
  END pe_in_pk_wrb_data__1_
  PIN pe_in_pk_wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.035 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0136 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 8.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M4 ; 
    ANTENNAMAXAREACAR 79.3082 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.802516 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.88679 LAYER V4 ;
  END pe_in_pk_wrb_data__0_
  PIN pe_in_pk_wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0416 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 14.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5592 LAYER M4 ; 
    ANTENNAMAXAREACAR 30.7524 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.309317 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.589153 LAYER V4 ;
  END pe_in_pk_wrb_addr__3_
  PIN pe_in_pk_wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 12.52 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1256 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7536 LAYER M4 ; 
    ANTENNAMAXAREACAR 22.6146 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.22642 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.33165 LAYER V4 ;
  END pe_in_pk_wrb_addr__2_
  PIN pe_in_pk_wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0254 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 11.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1192 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9936 LAYER M4 ; 
    ANTENNAMAXAREACAR 20.7069 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.210811 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.06091 LAYER V4 ;
  END pe_in_pk_wrb_addr__1_
  PIN pe_in_pk_wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 12.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1288 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7536 LAYER M4 ; 
    ANTENNAMAXAREACAR 26.4289 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.265337 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.33165 LAYER V4 ;
  END pe_in_pk_wrb_addr__0_
  PIN pe_in_pk_wrb__3_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 13 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1304 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M4 ; 
    ANTENNAMAXAREACAR 94.7399 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.954435 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.6129 LAYER V4 ;
  END pe_in_pk_wrb__3_
  PIN pe_in_pk_wrb__2_ 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 12.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1224 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.2412 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.457182 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.677507 LAYER V4 ;
  END pe_in_pk_wrb__2_
  PIN pe_in_pk_wrb__1_ 
    ANTENNAPARTIALMETALAREA 4.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0446 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 11.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M4 ; 
    ANTENNAMAXAREACAR 44.9702 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.454472 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.677507 LAYER V4 ;
  END pe_in_pk_wrb__1_
  PIN pe_in_pk_wrb__0_ 
    ANTENNAPARTIALMETALAREA 12.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1294 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0488 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0184 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER M4 ; 
    ANTENNAMAXAREACAR 11.0949 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.115718 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.677507 LAYER V4 ;
  END pe_in_pk_wrb__0_
  PIN pe_in_pk_rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.051 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0368 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 9.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0992 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3192 LAYER M4 ; 
    ANTENNAMAXAREACAR 36.5205 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.368147 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.01986 LAYER V4 ;
  END pe_in_pk_rdb_addr__3_
  PIN pe_in_pk_rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5304 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.0349 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.316064 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.903965 LAYER V3 ;
  END pe_in_pk_rdb_addr__2_
  PIN pe_in_pk_rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5304 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.6439 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.274941 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.35135 LAYER V3 ;
  END pe_in_pk_rdb_addr__1_
  PIN pe_in_pk_rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0262 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7368 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.4426 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.230003 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02041 LAYER V3 ;
  END pe_in_pk_rdb_addr__0_
  PIN pk_out_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0056 LAYER M3 ;
  END pk_out_PE_state__2_
  PIN pk_out_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 2.014 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M3 ;
  END pk_out_PE_state__1_
  PIN pk_out_PE_state__0_ 
    ANTENNADIFFAREA 2.014 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0566 LAYER M2 ;
  END pk_out_PE_state__0_
  PIN pk_out_data__7_ 
  END pk_out_data__7_
  PIN pk_out_data__6_ 
    ANTENNAPARTIALMETALAREA 2.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M3 ;
  END pk_out_data__6_
  PIN pk_out_data__5_ 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M3 ;
  END pk_out_data__5_
  PIN pk_out_data__4_ 
    ANTENNAPARTIALMETALAREA 1.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0392 LAYER M3 ;
  END pk_out_data__4_
  PIN pk_out_data__3_ 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0208 LAYER M3 ;
  END pk_out_data__3_
  PIN pk_out_data__2_ 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0246 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0592 LAYER M3 ;
  END pk_out_data__2_
  PIN pk_out_data__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0992 LAYER M3 ;
  END pk_out_data__1_
  PIN pk_out_data__0_ 
    ANTENNAPARTIALMETALAREA 3.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0382 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNADIFFAREA 1.76 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1304 LAYER M3 ;
  END pk_out_data__0_
END PE_POOL

END LIBRARY
