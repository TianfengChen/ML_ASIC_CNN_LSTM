

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO decoder 
  PIN clk 
    ANTENNAPARTIALMETALAREA 7.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0776 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2136 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.7463 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.384363 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.93633 LAYER V4 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0022 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 64.3829 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.66509 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END reset
  PIN CNTR_pk_in_PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0088 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 5.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0552 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 95.6892 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.973649 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_PE_state__2_
  PIN CNTR_pk_in_PE_state__1_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 68.2117 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.703378 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_PE_state__1_
  PIN CNTR_pk_in_PE_state__0_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 3.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0392 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 63.7072 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.658333 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_PE_state__0_
  PIN CNTR_pk_in_wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 4.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0408 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 57.8514 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.59527 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__7_
  PIN CNTR_pk_in_wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 49.7432 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.514189 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__6_
  PIN CNTR_pk_in_wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 1.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 3.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 61.455 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.631306 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__5_
  PIN CNTR_pk_in_wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.527 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.352027 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__4_
  PIN CNTR_pk_in_wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0168 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.2207 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.288964 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__3_
  PIN CNTR_pk_in_wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 1.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.5811 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.397072 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__2_
  PIN CNTR_pk_in_wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0696 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 87.5811 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.892568 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__1_
  PIN CNTR_pk_in_wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 31.2748 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.334009 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_data__0_
  PIN CNTR_pk_in_wrb_addr__7_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0168 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.4369 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.451126 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__7_
  PIN CNTR_pk_in_wrb_addr__6_ 
    ANTENNAPARTIALMETALAREA 0.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0096 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.482 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.406081 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__6_
  PIN CNTR_pk_in_wrb_addr__5_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 7.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.08 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 101.095 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.0277 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__5_
  PIN CNTR_pk_in_wrb_addr__4_ 
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0136 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 25.8694 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.279955 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__4_
  PIN CNTR_pk_in_wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.288964 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__3_
  PIN CNTR_pk_in_wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 1.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0472 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.509 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.676351 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__2_
  PIN CNTR_pk_in_wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0208 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.9775 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.361036 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__1_
  PIN CNTR_pk_in_wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 38.482 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.406081 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_addr__0_
  PIN CNTR_pk_in_wrb_ 
    ANTENNAPARTIALMETALAREA 1.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0168 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 27.6712 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.297973 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_wrb_
  PIN CNTR_pk_in_rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0048 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0632 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 80.3739 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.820495 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_rdb_addr__3_
  PIN CNTR_pk_in_rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 26.7703 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.288964 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_rdb_addr__2_
  PIN CNTR_pk_in_rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 5.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0544 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 82.1757 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.838514 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_rdb_addr__1_
  PIN CNTR_pk_in_rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0014 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M4 ; 
    ANTENNAMAXAREACAR 44.3378 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.460135 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.25225 LAYER V4 ;
  END CNTR_pk_in_rdb_addr__0_
  PIN CNN_pk_out_3__wrb__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M4 ;
  END CNN_pk_out_3__wrb__3_
  PIN CNN_pk_out_3__wrb__2_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02 LAYER M4 ;
  END CNN_pk_out_3__wrb__2_
  PIN CNN_pk_out_3__wrb__1_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0392 LAYER M4 ;
  END CNN_pk_out_3__wrb__1_
  PIN CNN_pk_out_3__wrb__0_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER M4 ;
  END CNN_pk_out_3__wrb__0_
  PIN CNN_pk_out_2__wrb__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0152 LAYER M4 ;
  END CNN_pk_out_2__wrb__3_
  PIN CNN_pk_out_2__wrb__2_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M4 ;
  END CNN_pk_out_2__wrb__2_
  PIN CNN_pk_out_2__wrb__1_ 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0264 LAYER M4 ;
  END CNN_pk_out_2__wrb__1_
  PIN CNN_pk_out_2__wrb__0_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M4 ;
  END CNN_pk_out_2__wrb__0_
  PIN CNN_pk_out_1__wrb__3_ 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0128 LAYER M4 ;
  END CNN_pk_out_1__wrb__3_
  PIN CNN_pk_out_1__wrb__2_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0144 LAYER M4 ;
  END CNN_pk_out_1__wrb__2_
  PIN CNN_pk_out_1__wrb__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02 LAYER M4 ;
  END CNN_pk_out_1__wrb__1_
  PIN CNN_pk_out_1__wrb__0_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0192 LAYER M4 ;
  END CNN_pk_out_1__wrb__0_
  PIN CNN_pk_out_0__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 30.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3048 LAYER M4 ;
  END CNN_pk_out_0__PE_state__2_
  PIN CNN_pk_out_1__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 30.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3048 LAYER M4 ;
  END CNN_pk_out_1__PE_state__2_
  PIN CNN_pk_out_2__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0014 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 30.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3048 LAYER M4 ;
  END CNN_pk_out_2__PE_state__2_
  PIN CNN_pk_out_3__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 30.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3048 LAYER M4 ;
  END CNN_pk_out_3__PE_state__2_
  PIN CNN_pk_out_0__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0904 LAYER M4 ;
  END CNN_pk_out_0__PE_state__1_
  PIN CNN_pk_out_1__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0904 LAYER M4 ;
  END CNN_pk_out_1__PE_state__1_
  PIN CNN_pk_out_2__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0904 LAYER M4 ;
  END CNN_pk_out_2__PE_state__1_
  PIN CNN_pk_out_3__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0904 LAYER M4 ;
  END CNN_pk_out_3__PE_state__1_
  PIN CNN_pk_out_0__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M4 ;
  END CNN_pk_out_0__PE_state__0_
  PIN CNN_pk_out_1__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M4 ;
  END CNN_pk_out_1__PE_state__0_
  PIN CNN_pk_out_2__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M4 ;
  END CNN_pk_out_2__PE_state__0_
  PIN CNN_pk_out_3__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0816 LAYER M4 ;
  END CNN_pk_out_3__PE_state__0_
  PIN CNN_pk_out_0__wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__7_
  PIN CNN_pk_out_1__wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__7_
  PIN CNN_pk_out_2__wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__7_
  PIN CNN_pk_out_3__wrb_data__7_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__7_
  PIN CNN_pk_out_0__wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0928 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__6_
  PIN CNN_pk_out_1__wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0928 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__6_
  PIN CNN_pk_out_2__wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0928 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__6_
  PIN CNN_pk_out_3__wrb_data__6_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0928 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__6_
  PIN CNN_pk_out_0__wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 26.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2632 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__5_
  PIN CNN_pk_out_1__wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 26.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2632 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__5_
  PIN CNN_pk_out_2__wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 0.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0006 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 26.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2632 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__5_
  PIN CNN_pk_out_3__wrb_data__5_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 26.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2632 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__5_
  PIN CNN_pk_out_0__wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__4_
  PIN CNN_pk_out_1__wrb_data__4_ 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__4_
  PIN CNN_pk_out_2__wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__4_
  PIN CNN_pk_out_3__wrb_data__4_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0432 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__4_
  PIN CNN_pk_out_0__wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2328 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__3_
  PIN CNN_pk_out_1__wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2328 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__3_
  PIN CNN_pk_out_2__wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2328 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__3_
  PIN CNN_pk_out_3__wrb_data__3_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.12 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2328 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__3_
  PIN CNN_pk_out_0__wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__2_
  PIN CNN_pk_out_1__wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__2_
  PIN CNN_pk_out_2__wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 1.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0168 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__2_
  PIN CNN_pk_out_3__wrb_data__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 15.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__2_
  PIN CNN_pk_out_0__wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__1_
  PIN CNN_pk_out_1__wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__1_
  PIN CNN_pk_out_2__wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__1_
  PIN CNN_pk_out_3__wrb_data__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 23.6 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2376 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__1_
  PIN CNN_pk_out_0__wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 20.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M4 ;
  END CNN_pk_out_0__wrb_data__0_
  PIN CNN_pk_out_1__wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 20.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M4 ;
  END CNN_pk_out_1__wrb_data__0_
  PIN CNN_pk_out_2__wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 20.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M4 ;
  END CNN_pk_out_2__wrb_data__0_
  PIN CNN_pk_out_3__wrb_data__0_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 20.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M4 ;
  END CNN_pk_out_3__wrb_data__0_
  PIN CNN_pk_out_0__wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 22.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2232 LAYER M4 ;
  END CNN_pk_out_0__wrb_addr__3_
  PIN CNN_pk_out_1__wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 22.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2232 LAYER M4 ;
  END CNN_pk_out_1__wrb_addr__3_
  PIN CNN_pk_out_2__wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 22.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2232 LAYER M4 ;
  END CNN_pk_out_2__wrb_addr__3_
  PIN CNN_pk_out_3__wrb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0046 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 22.16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2232 LAYER M4 ;
  END CNN_pk_out_3__wrb_addr__3_
  PIN CNN_pk_out_0__wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 27.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER M4 ;
  END CNN_pk_out_0__wrb_addr__2_
  PIN CNN_pk_out_1__wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0008 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 27.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER M4 ;
  END CNN_pk_out_1__wrb_addr__2_
  PIN CNN_pk_out_2__wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 27.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER M4 ;
  END CNN_pk_out_2__wrb_addr__2_
  PIN CNN_pk_out_3__wrb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 27.92 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER M4 ;
  END CNN_pk_out_3__wrb_addr__2_
  PIN CNN_pk_out_0__wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 24.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER M4 ;
  END CNN_pk_out_0__wrb_addr__1_
  PIN CNN_pk_out_1__wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 24.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER M4 ;
  END CNN_pk_out_1__wrb_addr__1_
  PIN CNN_pk_out_2__wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 24.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER M4 ;
  END CNN_pk_out_2__wrb_addr__1_
  PIN CNN_pk_out_3__wrb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 24.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER M4 ;
  END CNN_pk_out_3__wrb_addr__1_
  PIN CNN_pk_out_0__wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1216 LAYER M4 ;
  END CNN_pk_out_0__wrb_addr__0_
  PIN CNN_pk_out_1__wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1216 LAYER M4 ;
  END CNN_pk_out_1__wrb_addr__0_
  PIN CNN_pk_out_2__wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1216 LAYER M4 ;
  END CNN_pk_out_2__wrb_addr__0_
  PIN CNN_pk_out_3__wrb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1216 LAYER M4 ;
  END CNN_pk_out_3__wrb_addr__0_
  PIN CNN_pk_out_0__wrb__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M4 ;
  END CNN_pk_out_0__wrb__3_
  PIN CNN_pk_out_0__wrb__2_ 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNADIFFAREA 2.172 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0128 LAYER M4 ;
  END CNN_pk_out_0__wrb__2_
  PIN CNN_pk_out_0__wrb__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0176 LAYER M4 ;
  END CNN_pk_out_0__wrb__1_
  PIN CNN_pk_out_0__wrb__0_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.196 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.68 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M4 ;
  END CNN_pk_out_0__wrb__0_
  PIN CNN_pk_out_0__rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1624 LAYER M4 ;
  END CNN_pk_out_0__rdb_addr__3_
  PIN CNN_pk_out_1__rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1624 LAYER M4 ;
  END CNN_pk_out_1__rdb_addr__3_
  PIN CNN_pk_out_2__rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1624 LAYER M4 ;
  END CNN_pk_out_2__rdb_addr__3_
  PIN CNN_pk_out_3__rdb_addr__3_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1624 LAYER M4 ;
  END CNN_pk_out_3__rdb_addr__3_
  PIN CNN_pk_out_0__rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1016 LAYER M4 ;
  END CNN_pk_out_0__rdb_addr__2_
  PIN CNN_pk_out_1__rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1016 LAYER M4 ;
  END CNN_pk_out_1__rdb_addr__2_
  PIN CNN_pk_out_2__rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1016 LAYER M4 ;
  END CNN_pk_out_2__rdb_addr__2_
  PIN CNN_pk_out_3__rdb_addr__2_ 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1016 LAYER M4 ;
  END CNN_pk_out_3__rdb_addr__2_
  PIN CNN_pk_out_0__rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M4 ;
  END CNN_pk_out_0__rdb_addr__1_
  PIN CNN_pk_out_1__rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M4 ;
  END CNN_pk_out_1__rdb_addr__1_
  PIN CNN_pk_out_2__rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M4 ;
  END CNN_pk_out_2__rdb_addr__1_
  PIN CNN_pk_out_3__rdb_addr__1_ 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0014 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER M4 ;
  END CNN_pk_out_3__rdb_addr__1_
  PIN CNN_pk_out_0__rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1696 LAYER M4 ;
  END CNN_pk_out_0__rdb_addr__0_
  PIN CNN_pk_out_1__rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1696 LAYER M4 ;
  END CNN_pk_out_1__rdb_addr__0_
  PIN CNN_pk_out_2__rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0016 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1696 LAYER M4 ;
  END CNN_pk_out_2__rdb_addr__0_
  PIN CNN_pk_out_3__rdb_addr__0_ 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 16.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1696 LAYER M4 ;
  END CNN_pk_out_3__rdb_addr__0_
END decoder

END LIBRARY
