

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO wb_controller 
  PIN clk 
    ANTENNAPARTIALMETALAREA 12.7 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1286 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2696 LAYER M4 ; 
    ANTENNAMAXAREACAR 112.833 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.14215 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.71901 LAYER V4 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 1.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.672 LAYER M4 ; 
    ANTENNAMAXAREACAR 76.5483 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.768033 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.736532 LAYER V4 ;
  END reset
  PIN DRAM_wbegin_sft[15] 
    ANTENNAPARTIALMETALAREA 6.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 43.1343 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.440162 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END DRAM_wbegin_sft[15]
  PIN DRAM_wbegin_sft[14] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.027 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 29.5926 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.304745 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END DRAM_wbegin_sft[14]
  PIN DRAM_wbegin_sft[13] 
    ANTENNAPARTIALMETALAREA 6.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0612 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 39.1991 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.40081 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END DRAM_wbegin_sft[13]
  PIN DRAM_wbegin_sft[12] 
    ANTENNAPARTIALMETALAREA 7.7 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0778 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 65.2407 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.663542 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END DRAM_wbegin_sft[12]
  PIN DRAM_wbegin_sft[11] 
    ANTENNAPARTIALMETALAREA 5.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0552 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.5787 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.384606 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[11]
  PIN DRAM_wbegin_sft[10] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0238 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 41.1667 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.420486 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[10]
  PIN DRAM_wbegin_sft[9] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 111.421 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.12303 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END DRAM_wbegin_sft[9]
  PIN DRAM_wbegin_sft[8] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0026 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 22.1852 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.228356 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[8]
  PIN DRAM_wbegin_sft[7] 
    ANTENNAPARTIALMETALAREA 6.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 50.7731 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.514236 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END DRAM_wbegin_sft[7]
  PIN DRAM_wbegin_sft[6] 
    ANTENNAPARTIALMETALAREA 1.58 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0158 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.8981 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.295486 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[6]
  PIN DRAM_wbegin_sft[5] 
    ANTENNAPARTIALMETALAREA 5.84 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 81.0972 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.822106 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[5]
  PIN DRAM_wbegin_sft[4] 
    ANTENNAPARTIALMETALAREA 6.5 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0658 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 49.037 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.501505 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[4]
  PIN DRAM_wbegin_sft[3] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 37.1157 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.379977 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END DRAM_wbegin_sft[3]
  PIN DRAM_wbegin_sft[2] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0486 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 129.593 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.30475 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END DRAM_wbegin_sft[2]
  PIN DRAM_wbegin_sft[1] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0236 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 35.2639 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.359144 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V4 ;
  END DRAM_wbegin_sft[1]
  PIN DRAM_wbegin_sft[0] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0378 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 40.7778 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.418403 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.15741 LAYER V4 ;
  END DRAM_wbegin_sft[0]
  PIN pk_out_3__PE_state__2_ 
  END pk_out_3__PE_state__2_
  PIN pk_out_3__PE_state__1_ 
  END pk_out_3__PE_state__1_
  PIN pk_out_3__PE_state__0_ 
  END pk_out_3__PE_state__0_
  PIN pk_out_3__data__7_ 
  END pk_out_3__data__7_
  PIN pk_out_3__data__6_ 
  END pk_out_3__data__6_
  PIN pk_out_3__data__5_ 
  END pk_out_3__data__5_
  PIN pk_out_3__data__4_ 
  END pk_out_3__data__4_
  PIN pk_out_3__data__3_ 
  END pk_out_3__data__3_
  PIN pk_out_3__data__2_ 
  END pk_out_3__data__2_
  PIN pk_out_3__data__1_ 
  END pk_out_3__data__1_
  PIN pk_out_3__data__0_ 
  END pk_out_3__data__0_
  PIN pk_out_2__PE_state__2_ 
  END pk_out_2__PE_state__2_
  PIN pk_out_2__PE_state__1_ 
  END pk_out_2__PE_state__1_
  PIN pk_out_2__PE_state__0_ 
  END pk_out_2__PE_state__0_
  PIN pk_out_2__data__7_ 
  END pk_out_2__data__7_
  PIN pk_out_2__data__6_ 
  END pk_out_2__data__6_
  PIN pk_out_2__data__5_ 
  END pk_out_2__data__5_
  PIN pk_out_2__data__4_ 
  END pk_out_2__data__4_
  PIN pk_out_2__data__3_ 
  END pk_out_2__data__3_
  PIN pk_out_2__data__2_ 
  END pk_out_2__data__2_
  PIN pk_out_2__data__1_ 
  END pk_out_2__data__1_
  PIN pk_out_2__data__0_ 
  END pk_out_2__data__0_
  PIN pk_out_1__PE_state__2_ 
  END pk_out_1__PE_state__2_
  PIN pk_out_1__PE_state__1_ 
  END pk_out_1__PE_state__1_
  PIN pk_out_1__PE_state__0_ 
  END pk_out_1__PE_state__0_
  PIN pk_out_1__data__7_ 
  END pk_out_1__data__7_
  PIN pk_out_1__data__6_ 
  END pk_out_1__data__6_
  PIN pk_out_1__data__5_ 
  END pk_out_1__data__5_
  PIN pk_out_1__data__4_ 
  END pk_out_1__data__4_
  PIN pk_out_1__data__3_ 
  END pk_out_1__data__3_
  PIN pk_out_1__data__2_ 
  END pk_out_1__data__2_
  PIN pk_out_1__data__1_ 
  END pk_out_1__data__1_
  PIN pk_out_1__data__0_ 
  END pk_out_1__data__0_
  PIN pk_out_0__PE_state__2_ 
    ANTENNAPARTIALMETALAREA 2.6024 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02596 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.312 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.28462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.095 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.384615 LAYER V3 ;
  END pk_out_0__PE_state__2_
  PIN pk_out_0__PE_state__1_ 
    ANTENNAPARTIALMETALAREA 2.2824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02276 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.166 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.174462 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.806452 LAYER V3 ;
  END pk_out_0__PE_state__1_
  PIN pk_out_0__PE_state__0_ 
    ANTENNAPARTIALMETALAREA 2.3224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02356 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.412 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.188038 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.07527 LAYER V3 ;
  END pk_out_0__PE_state__0_
  PIN pk_out_0__data__7_ 
    ANTENNAPARTIALMETALAREA 4.2824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04276 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 109.194 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.09525 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END pk_out_0__data__7_
  PIN pk_out_0__data__6_ 
    ANTENNAPARTIALMETALAREA 2.9624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02996 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.0741 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.206366 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END pk_out_0__data__6_
  PIN pk_out_0__data__5_ 
    ANTENNAPARTIALMETALAREA 4.2824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04276 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 21.2176 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.222801 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.925926 LAYER V4 ;
  END pk_out_0__data__5_
  PIN pk_out_0__data__4_ 
    ANTENNAPARTIALMETALAREA 2.844 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02884 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.4815 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.25081 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END pk_out_0__data__4_
  PIN pk_out_0__data__3_ 
    ANTENNAPARTIALMETALAREA 3.1224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03156 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.6111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.201736 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END pk_out_0__data__3_
  PIN pk_out_0__data__2_ 
    ANTENNAPARTIALMETALAREA 4.5624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04596 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.13229 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V3 ;
  END pk_out_0__data__2_
  PIN pk_out_0__data__1_ 
    ANTENNAPARTIALMETALAREA 5.9624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0184 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M4 ; 
    ANTENNAMAXAREACAR 14.0417 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.148727 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V4 ;
  END pk_out_0__data__1_
  PIN pk_out_0__data__0_ 
    ANTENNAPARTIALMETALAREA 2.9624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02996 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.537 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.210995 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V3 ;
  END pk_out_0__data__0_
  PIN DRAM_in3_Data__7_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.58 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0458 LAYER M4 ;
  END DRAM_in3_Data__7_
  PIN DRAM_in3_Data__6_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.034 LAYER M4 ;
  END DRAM_in3_Data__6_
  PIN DRAM_in3_Data__5_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0326 LAYER M4 ;
  END DRAM_in3_Data__5_
  PIN DRAM_in3_Data__4_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.48 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0656 LAYER M4 ;
  END DRAM_in3_Data__4_
  PIN DRAM_in3_Data__3_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0322 LAYER M4 ;
  END DRAM_in3_Data__3_
  PIN DRAM_in3_Data__2_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 1.24 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0124 LAYER M4 ;
  END DRAM_in3_Data__2_
  PIN DRAM_in3_Data__1_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.14 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1118 LAYER M4 ;
  END DRAM_in3_Data__1_
  PIN DRAM_in3_Data__0_ 
    ANTENNADIFFAREA 2.112 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.96 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04 LAYER M4 ;
  END DRAM_in3_Data__0_
  PIN DRAM_in3_WEN_ 
    ANTENNADIFFAREA 3.52 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.76 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.028 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5592 LAYER M4 ; 
    ANTENNAMAXAREACAR 12.5473 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.130169 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.647249 LAYER V4 ;
  END DRAM_in3_WEN_
  PIN DRAM_in3_Addr__15_ 
    ANTENNADIFFAREA 1.728 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.58 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.077 LAYER M4 ;
  END DRAM_in3_Addr__15_
  PIN DRAM_in3_Addr__14_ 
    ANTENNADIFFAREA 0.996 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0244 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M4 ; 
    ANTENNAMAXAREACAR 92.0905 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.945977 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.72414 LAYER V4 ;
  END DRAM_in3_Addr__14_
  PIN DRAM_in3_Addr__13_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.74 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0582 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 82.035 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.841958 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.29885 LAYER V4 ;
  END DRAM_in3_Addr__13_
  PIN DRAM_in3_Addr__12_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0264 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 78.1321 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.797182 LAYER M4 ;
    ANTENNAMAXCUTCAR 5.17241 LAYER V4 ;
  END DRAM_in3_Addr__12_
  PIN DRAM_in3_Addr__11_ 
    ANTENNADIFFAREA 3.2 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.025 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2184 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.6683 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.470008 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.51573 LAYER V4 ;
  END DRAM_in3_Addr__11_
  PIN DRAM_in3_Addr__10_ 
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.08 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0212 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 116.241 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.17106 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.87356 LAYER V4 ;
  END DRAM_in3_Addr__10_
  PIN DRAM_in3_Addr__9_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.9 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0494 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 89.4079 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.920292 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER V4 ;
  END DRAM_in3_Addr__9_
  PIN DRAM_in3_Addr__8_ 
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0232 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER M4 ; 
    ANTENNAMAXAREACAR 103.554 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 1.06716 LAYER M4 ;
    ANTENNAMAXCUTCAR 6.32184 LAYER V4 ;
  END DRAM_in3_Addr__8_
  PIN DRAM_in3_Addr__7_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.065 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 95.0093 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.964813 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER V4 ;
  END DRAM_in3_Addr__7_
  PIN DRAM_in3_Addr__6_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0244 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER M4 ; 
    ANTENNAMAXAREACAR 34.2601 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.352835 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.22955 LAYER V4 ;
  END DRAM_in3_Addr__6_
  PIN DRAM_in3_Addr__5_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 90.4786 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.925252 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER V4 ;
  END DRAM_in3_Addr__5_
  PIN DRAM_in3_Addr__4_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.04 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0608 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 87.4889 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.895355 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER V4 ;
  END DRAM_in3_Addr__4_
  PIN DRAM_in3_Addr__3_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0506 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 62.5105 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.647855 LAYER M4 ;
    ANTENNAMAXCUTCAR 4.02299 LAYER V4 ;
  END DRAM_in3_Addr__3_
  PIN DRAM_in3_Addr__2_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.4 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0548 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 LAYER M4 ; 
    ANTENNAMAXAREACAR 53.6241 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.545266 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.51779 LAYER V4 ;
  END DRAM_in3_Addr__2_
  PIN DRAM_in3_Addr__1_ 
    ANTENNADIFFAREA 2.014 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0028 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3504 LAYER M4 ; 
    ANTENNAMAXAREACAR 15.6852 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.168107 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.95245 LAYER V4 ;
  END DRAM_in3_Addr__1_
  PIN DRAM_in3_Addr__0_ 
    ANTENNADIFFAREA 4.168 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 3.72 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0376 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER M4 ; 
    ANTENNAMAXAREACAR 30.9679 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.315925 LAYER M4 ;
    ANTENNAMAXCUTCAR 1.60437 LAYER V4 ;
  END DRAM_in3_Addr__0_
END wb_controller

END LIBRARY
