* SPICE NETLIST
***************************************

.SUBCKT esdscr A K PD SX
.ENDS
***************************************
.SUBCKT subc SUBCON SUB
.ENDS
***************************************
.SUBCKT nfettw G S D B PI sx
.ENDS
***************************************
.SUBCKT dgnfettw G S D B PI sx
.ENDS
***************************************
.SUBCKT nfet33tw G S D B PI sx
.ENDS
***************************************
.SUBCKT hvtnfet33tw G S D B PI sx
.ENDS
***************************************
.SUBCKT lvtnfettw G S D B PI sx
.ENDS
***************************************
.SUBCKT lpnfettw G S D B PI sx
.ENDS
***************************************
.SUBCKT nfettw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT dgnfettw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT hvtnfet33tw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT lvtnfettw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT nfet33tw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT lpnfettw_rf G S D B PI sx
.ENDS
***************************************
.SUBCKT sblkndres D S G
.ENDS
***************************************
.SUBCKT ncap G S B D
.ENDS
***************************************
.SUBCKT dgncap G S B D
.ENDS
***************************************
.SUBCKT diffhavar ANODE1 ANODE2 CATHODE BULK
.ENDS
***************************************
.SUBCKT diffncap GA GB NW SX
.ENDS
***************************************
.SUBCKT esdnsh_base d g s b
.ENDS
***************************************
.SUBCKT esdpsh_base d g s b
.ENDS
***************************************
.SUBCKT bondpad in gp sub
.ENDS
***************************************
.SUBCKT devicepad pad
.ENDS
***************************************
.SUBCKT efuse IN OUT
.ENDS
***************************************
.SUBCKT indp out in bulk
.ENDS
***************************************
.SUBCKT ind out in bulk
.ENDS
***************************************
.SUBCKT inds out in bulk
.ENDS
***************************************
.SUBCKT symindp outpr outse ct BULK
.ENDS
***************************************
.SUBCKT symind outpr outse ct BULK
.ENDS
***************************************
.SUBCKT rfline in out bulk
.ENDS
***************************************
.SUBCKT singlewire VA VB VSHIELD
.ENDS
***************************************
.SUBCKT coupledwires VA1 VA2 VB1 VB2 VSHIELD
.ENDS
***************************************
.SUBCKT singlecpw va vb vshield
.ENDS
***************************************
.SUBCKT coupledcpw va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT corrPoint cp
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=308 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=976 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=4088 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=4014 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=4887 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=4914 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PCORNER
** N=17 EP=0 IP=47 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD DVSS VDD
.ENDS
***************************************
.SUBCKT ICV_148
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT fillqbp_i
** N=102 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS
.ENDS
***************************************
.SUBCKT PFILLH
** N=5124 EP=0 IP=4 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVSS DVDD VDD
.ENDS
***************************************
.SUBCKT ICV_262
** N=4 EP=0 IP=16 FDC=0
.ENDS
***************************************
.SUBCKT ICV_145
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_261
** N=4 EP=0 IP=32 FDC=0
.ENDS
***************************************
.SUBCKT PFILLQ
** N=2664 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVSS DVDD VDD
.ENDS
***************************************
.SUBCKT PFILL1
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVSS DVDD VDD
.ENDS
***************************************
.SUBCKT ppoly_res_w2_l25 1 2 3
** N=13 EP=3 IP=0 FDC=1
R0 1 2 4371.76 L=2.5e-05 W=2e-06 sbar=1 m=1 par=1 bp=3 $SUB=3 $[opppcres] $X=0 $Y=590 $D=355
.ENDS
***************************************
.SUBCKT ICV_151 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 ppoly_res_w2_l25 $T=0 0 0 0 $X=-320 $Y=-300
X1 1 3 4 ppoly_res_w2_l25 $T=2800 0 0 0 $X=2480 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_152 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_151 $T=0 0 0 0 $X=-320 $Y=-300
X1 4 3 5 6 ICV_151 $T=5600 0 0 0 $X=5280 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_153 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=8
X0 1 2 3 4 5 10 ICV_152 $T=0 0 0 0 $X=-320 $Y=-300
X1 6 5 7 8 9 10 ICV_152 $T=11200 0 0 0 $X=10880 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_2 1 VSS 3
** N=2176 EP=3 IP=32 FDC=24
X0 14 8 9 15 3 VSS ICV_152 $T=33550 79300 0 90 $X=7070 $Y=78980
X1 20 25 26 21 1 VSS ICV_152 $T=36450 79300 1 90 $X=36150 $Y=78980
X2 10 4 5 11 6 12 7 13 8 VSS ICV_153 $T=33550 56900 0 90 $X=7070 $Y=56580
X3 16 4 22 17 23 18 24 19 25 VSS ICV_153 $T=36450 56900 1 90 $X=36150 $Y=56580
.ENDS
***************************************
.SUBCKT ICV_3 VSS DVDD 5
** N=27458 EP=3 IP=0 FDC=196
*.CALIBRE ISOLATED NETS: DVSS VDD
M0 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=5370 $D=106
M1 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=6050 $D=106
M2 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=6730 $D=106
M3 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=7410 $D=106
M4 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=8090 $D=106
M5 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=8770 $D=106
M6 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=9450 $D=106
M7 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=10130 $D=106
M8 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=10810 $D=106
M9 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=11490 $D=106
M10 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=12170 $D=106
M11 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=12850 $D=106
M12 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=13530 $D=106
M13 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=14210 $D=106
M14 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=14890 $D=106
M15 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=17910 $D=106
M16 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=18590 $D=106
M17 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=19270 $D=106
M18 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=19950 $D=106
M19 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=20630 $D=106
M20 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=21310 $D=106
M21 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=21990 $D=106
M22 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=22670 $D=106
M23 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=23350 $D=106
M24 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=24030 $D=106
M25 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=24710 $D=106
M26 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=25390 $D=106
M27 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=26070 $D=106
M28 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=26750 $D=106
M29 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=27430 $D=106
M30 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=30450 $D=106
M31 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=31130 $D=106
M32 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=31810 $D=106
M33 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=32490 $D=106
M34 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=33170 $D=106
M35 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=33850 $D=106
M36 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=34530 $D=106
M37 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=35210 $D=106
M38 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=35890 $D=106
M39 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=36570 $D=106
M40 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=37250 $D=106
M41 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=37930 $D=106
M42 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=38610 $D=106
M43 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=39290 $D=106
M44 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=39970 $D=106
M45 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=42990 $D=106
M46 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=43670 $D=106
M47 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=44350 $D=106
M48 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=45030 $D=106
M49 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=45710 $D=106
M50 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=46390 $D=106
M51 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=47070 $D=106
M52 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=47750 $D=106
M53 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=48430 $D=106
M54 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=49110 $D=106
M55 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=49790 $D=106
M56 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=50470 $D=106
M57 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=51150 $D=106
M58 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=51830 $D=106
M59 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=52510 $D=106
M60 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=55530 $D=106
M61 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=56210 $D=106
M62 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=56890 $D=106
M63 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=57570 $D=106
M64 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=58250 $D=106
M65 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=58930 $D=106
M66 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=59610 $D=106
M67 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=60290 $D=106
M68 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=60970 $D=106
M69 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=61650 $D=106
M70 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=62330 $D=106
M71 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=63010 $D=106
M72 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=63690 $D=106
M73 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=64370 $D=106
M74 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=65050 $D=106
M75 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=68810 $D=106
M76 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=69490 $D=106
M77 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=70170 $D=106
M78 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=70850 $D=106
M79 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=5370 $D=106
M80 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=6050 $D=106
M81 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=6730 $D=106
M82 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=7410 $D=106
M83 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=8090 $D=106
M84 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=8770 $D=106
M85 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=9450 $D=106
M86 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=10130 $D=106
M87 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=10810 $D=106
M88 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=11490 $D=106
M89 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=12170 $D=106
M90 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=12850 $D=106
M91 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=13530 $D=106
M92 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=14210 $D=106
M93 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=14890 $D=106
M94 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=17910 $D=106
M95 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=18590 $D=106
M96 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=19270 $D=106
M97 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=19950 $D=106
M98 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=20630 $D=106
M99 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=21310 $D=106
M100 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=21990 $D=106
M101 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=22670 $D=106
M102 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=23350 $D=106
M103 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=24030 $D=106
M104 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=24710 $D=106
M105 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=25390 $D=106
M106 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=26070 $D=106
M107 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=26750 $D=106
M108 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=27430 $D=106
M109 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=30450 $D=106
M110 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=31130 $D=106
M111 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=31810 $D=106
M112 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=32490 $D=106
M113 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=33170 $D=106
M114 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=33850 $D=106
M115 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=34530 $D=106
M116 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=35210 $D=106
M117 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=35890 $D=106
M118 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=36570 $D=106
M119 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=37250 $D=106
M120 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=37930 $D=106
M121 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=38610 $D=106
M122 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=39290 $D=106
M123 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=39970 $D=106
M124 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=42990 $D=106
M125 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=43670 $D=106
M126 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=44350 $D=106
M127 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=45030 $D=106
M128 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=45710 $D=106
M129 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=46390 $D=106
M130 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=47070 $D=106
M131 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=47750 $D=106
M132 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=48430 $D=106
M133 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=49110 $D=106
M134 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=49790 $D=106
M135 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=50470 $D=106
M136 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=51150 $D=106
M137 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=51830 $D=106
M138 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=52510 $D=106
M139 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=55530 $D=106
M140 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=56210 $D=106
M141 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=56890 $D=106
M142 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=57570 $D=106
M143 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=58250 $D=106
M144 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=58930 $D=106
M145 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=59610 $D=106
M146 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=60290 $D=106
M147 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=60970 $D=106
M148 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=61650 $D=106
M149 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=62330 $D=106
M150 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=63010 $D=106
M151 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=63690 $D=106
M152 VSS 6 DVDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=64370 $D=106
M153 DVDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=65050 $D=106
M154 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=68810 $D=106
M155 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=69490 $D=106
M156 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=70170 $D=106
M157 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=70850 $D=106
M158 6 5 DVDD DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=68810 $D=193
M159 DVDD 5 6 DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=69490 $D=193
M160 6 5 DVDD DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=70170 $D=193
M161 DVDD 5 6 DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=70850 $D=193
M162 6 5 DVDD DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=68810 $D=193
M163 DVDD 5 6 DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=69490 $D=193
M164 6 5 DVDD DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=70170 $D=193
M165 DVDD 5 6 DVDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=70850 $D=193
X166 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=76490 $D=397
X167 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=84470 $D=397
X168 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=92450 $D=397
X169 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=100430 $D=397
X170 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=108410 $D=397
X171 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=116390 $D=397
X172 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=76490 $D=397
X173 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=84470 $D=397
X174 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=92450 $D=397
X175 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=100430 $D=397
X176 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=108410 $D=397
X177 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=116390 $D=397
X178 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=76490 $D=397
X179 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=84470 $D=397
X180 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=92450 $D=397
X181 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=100430 $D=397
X182 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=108410 $D=397
X183 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=116390 $D=397
X184 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=76490 $D=397
X185 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=84470 $D=397
X186 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=92450 $D=397
X187 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=100430 $D=397
X188 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=108410 $D=397
X189 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=116390 $D=397
X190 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=76490 $D=397
X191 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=84470 $D=397
X192 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=92450 $D=397
X193 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=100430 $D=397
X194 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=108410 $D=397
X195 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=116390 $D=397
.ENDS
***************************************
.SUBCKT PDVDD VSS DVSS DVDD VDD
** N=5 EP=4 IP=8 FDC=220
X0 DVDD VSS 5 ICV_2 $T=0 0 0 0 $X=-140 $Y=0
X1 VSS DVDD 5 ICV_3 $T=0 117000 0 0 $X=-140 $Y=117000
.ENDS
***************************************
.SUBCKT ICV_176
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT dvssbp_i
** N=1785 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS
.ENDS
***************************************
.SUBCKT ICV_26
** N=1812 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=2067 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=1952 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1394 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=786 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=2112 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1309 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1590 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nc_grounds_l
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: pad vss_dvss_l1
.ENDS
***************************************
.SUBCKT nc_grounds_r
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_l1 pad
.ENDS
***************************************
.SUBCKT dvss_oly
** N=20 EP=0 IP=57 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS VDD DVSS
.ENDS
***************************************
.SUBCKT mc2_grounds_capl
** N=60 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS
.ENDS
***************************************
.SUBCKT ipplscp_dvss_sub
** N=1639 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ipplscp_dvss
** N=4628 EP=0 IP=2628 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD DVSS
.ENDS
***************************************
.SUBCKT bc_grounds_cnrl
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS pad
.ENDS
***************************************
.SUBCKT nc_grounds_capl
** N=1 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS
.ENDS
***************************************
.SUBCKT bc_grounds_l
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: pad vss_dvss_l1
.ENDS
***************************************
.SUBCKT mc2_grounds_l
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: pad vss_dvss_l1 DVDD
.ENDS
***************************************
.SUBCKT bc_grounds
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_l1 pad vss_dvss_r1
.ENDS
***************************************
.SUBCKT ICV_18
** N=3 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT nc_grounds
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_l1 pad vss_dvss_r1
.ENDS
***************************************
.SUBCKT ICV_17
** N=3 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT mc2_grounds
** N=5 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_l1 pad vss_dvss_r1
.ENDS
***************************************
.SUBCKT ICV_16
** N=4 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT bc_grounds_r
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_r1 pad
.ENDS
***************************************
.SUBCKT mc2_grounds_r
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: vss_dvss_r1 pad
.ENDS
***************************************
.SUBCKT PDVSS VSS DVSS DVDD VDD
** N=4 EP=4 IP=67 FDC=0
.ENDS
***************************************
.SUBCKT mc2_capl
** N=127 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD well_cntrl_res DVSS ng1 ng0 sdlow poff pg1 pg0
.ENDS
***************************************
.SUBCKT bc_cnrl
** N=21 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS ng1 ng0 pad sdlow
.ENDS
***************************************
.SUBCKT nct_capl
** N=240 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVSS VSS ng1 ng0 sdlow sdhigh
.ENDS
***************************************
.SUBCKT nct DVSS pad ntr0m2 ntr1m2 sdhigh 10 11
** N=144 EP=7 IP=0 FDC=6
*.CALIBRE ISOLATED NETS: sdlow ng1 ng0
M0 10 ntr0m2 DVSS DVSS dgnfet L=2.4e-07 W=1.642e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=370 $D=106
M1 13 sdhigh 10 DVSS dgnfet L=2.4e-07 W=1.642e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1220 $Y=370 $D=106
M2 11 sdhigh 14 DVSS dgnfet L=2.4e-07 W=1.642e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8540 $Y=370 $D=106
M3 DVSS ntr1m2 11 DVSS dgnfet L=2.4e-07 W=1.642e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9380 $Y=370 $D=106
X4 13 pad DVSS sblkndres w=1.642e-05 l=2e-06 r=9.64238 sbar=1 m=1 par=1 $X=2100 $Y=370 $D=350
X5 pad 14 DVSS sblkndres w=1.642e-05 l=2e-06 r=9.64238 sbar=1 m=1 par=1 $X=5900 $Y=370 $D=350
.ENDS
***************************************
.SUBCKT mc2l
** N=49 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD well_cntrl_res pad
.ENDS
***************************************
.SUBCKT bc
** N=10 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS pad
.ENDS
***************************************
.SUBCKT mc2
** N=53 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD well_cntrl_res pad
.ENDS
***************************************
.SUBCKT mc2r
** N=49 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD well_cntrl_res pad
.ENDS
***************************************
.SUBCKT mc2_capr
** N=124 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD well_cntrl_res ng0 ng1 pg0 pg1 sdhigh
.ENDS
***************************************
.SUBCKT nct_capr
** N=240 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVSS ng0 ng1 VSS DVDD sdhigh sdlow
.ENDS
***************************************
.SUBCKT bc_cnrr
** N=21 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS pad ng0 ng1 sdhigh
.ENDS
***************************************
.SUBCKT ICV_40 2 5 6 7 11
** N=2720 EP=5 IP=179 FDC=36
X3 2 7 6 5 11 12 13 nct $T=5000 121510 0 0 $X=3420 $Y=121360
X4 2 7 5 5 11 14 15 nct $T=15000 121510 0 0 $X=13420 $Y=121360
X5 2 7 5 5 11 16 17 nct $T=25000 121510 0 0 $X=23420 $Y=121360
X6 2 7 5 5 11 18 19 nct $T=35000 121510 0 0 $X=33420 $Y=121360
X7 2 7 5 5 11 20 21 nct $T=45000 121510 0 0 $X=43420 $Y=121360
X8 2 7 5 5 11 22 23 nct $T=55000 121510 0 0 $X=53420 $Y=121360
.ENDS
***************************************
.SUBCKT ppoly_res_250 1 2 3
** N=23 EP=3 IP=0 FDC=1
R0 1 2 249.937 L=2.6e-06 W=4e-06 sbar=1 m=1 par=1 bp=3 $SUB=3 $[opppcres] $X=0 $Y=590 $D=355
.ENDS
***************************************
.SUBCKT sc4 DVDD VSS sdlow well_cntrl_res poff oeb_3v3 n1_buf t3iR t3oR t2iR t2oR pgR t1oR t1iR t0iR t0oR ndisR psrc nsrc pg1
+ pg0 t3iL t3oL t2iL t2oL pgL t1iL t1oL t0iL t0oL ndisL sdhigh psupply pctrl VDD pad pd_en well_en_ pu_en_tol_ nctrl
+ plvl inxfr alow
** N=4232 EP=43 IP=6 FDC=94
*.CALIBRE ISOLATED NETS: ng0 ng1
M0 53 oeb_3v3 VSS VSS dgnfet L=8e-06 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-2380 $Y=20950 $D=106
M1 64 pd_en VSS VSS dgnfet L=8e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1530 $Y=19290 $D=106
M2 47 52 64 VSS dgnfet L=8e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-410 $Y=19290 $D=106
M3 65 52 51 VSS dgnfet L=1e-06 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3390 $Y=19290 $D=106
M4 VSS n1_buf 65 VSS dgnfet L=1e-06 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4690 $Y=19290 $D=106
M5 poff 52 52 VSS dgnfet L=2.4e-07 W=1.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7240 $Y=22290 $D=106
M6 t1iR sdhigh t1oR VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7410 $Y=19290 $D=106
M7 52 52 poff VSS dgnfet L=2.4e-07 W=1.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7940 $Y=22290 $D=106
M8 t0oR sdhigh t0iR VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9170 $Y=19290 $D=106
M9 nsrc nctrl ndisR VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10930 $Y=19290 $D=106
M10 ndisR nctrl nsrc VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11650 $Y=19290 $D=106
M11 nsrc nctrl ndisR VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12370 $Y=19290 $D=106
M12 57 57 53 VSS dgnfet L=6e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12940 $Y=25690 $D=106
M13 ndisR nctrl nsrc VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=13090 $Y=19290 $D=106
M14 48 48 57 VSS dgnfet L=2e-06 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=14270 $Y=25590 $D=106
M15 56 oeb_3v3 VSS VSS dgnfet L=1e-06 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15150 $Y=23470 $D=106
M16 nsrc nctrl ndisL VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15890 $Y=19290 $D=106
M17 ndisL nctrl nsrc VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16610 $Y=19290 $D=106
M18 54 57 56 VSS dgnfet L=2e-06 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17050 $Y=23470 $D=106
M19 nsrc nctrl ndisL VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17330 $Y=19290 $D=106
M20 ndisL nctrl nsrc VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18050 $Y=19290 $D=106
M21 60 oeb_3v3 VSS VSS dgnfet L=2.4e-07 W=7.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18630 $Y=21890 $D=106
M22 VSS oeb_3v3 60 VSS dgnfet L=2.4e-07 W=7.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19310 $Y=21890 $D=106
M23 t0iL sdhigh t0oL VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19810 $Y=19290 $D=106
M24 61 60 VSS VSS dgnfet L=2.4e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20310 $Y=21790 $D=106
M25 61 54 VSS VSS dgnfet L=2.4e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20920 $Y=23690 $D=106
M26 t1iL sdhigh t1oL VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=21570 $Y=19290 $D=106
M27 VSS 61 n1_buf VSS dgnfet L=2.4e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=22660 $Y=23350 $D=106
M28 psupply sdhigh 55 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23530 $Y=19290 $D=106
M29 62 n1_buf VSS VSS dgnfet L=2.4e-07 W=1.6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23600 $Y=22450 $D=106
M30 46 62 50 VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=25360 $Y=19050 $D=106
M31 50 62 46 VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26060 $Y=19050 $D=106
M32 inxfr sdhigh 47 VSS dgnfet L=2.4e-07 W=4.94e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=28000 $Y=19110 $D=106
M33 47 sdhigh inxfr VSS dgnfet L=2.4e-07 W=4.94e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=28700 $Y=19110 $D=106
M34 63 n1_buf VSS VSS dgnfet L=3e-06 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30640 $Y=19110 $D=106
M35 63 oeb_3v3 pctrl VSS dgnfet L=3e-06 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30640 $Y=20640 $D=106
M36 poff 46 47 well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-2990 $Y=7990 $D=193
M37 48 49 48 48 dgpfet L=1e-06 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-2800 $Y=24870 $D=193
M38 47 46 poff well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-2290 $Y=7990 $D=193
M39 48 49 48 48 dgpfet L=1e-06 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1340 $Y=24870 $D=193
M40 DVDD well_en_ well_cntrl_res well_cntrl_res dgpfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-450 $Y=8820 $D=193
M41 48 VSS 48 48 dgpfet L=1e-06 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=120 $Y=24870 $D=193
M42 well_cntrl_res well_en_ DVDD well_cntrl_res dgpfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=250 $Y=8820 $D=193
M43 48 VSS 48 48 dgpfet L=1e-06 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1580 $Y=24870 $D=193
M44 47 46 well_en_ well_cntrl_res dgpfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2090 $Y=10990 $D=193
M45 52 pctrl poff well_cntrl_res dgpfet L=2.4e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2840 $Y=8520 $D=193
M46 51 46 47 well_cntrl_res dgpfet L=2.4e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3030 $Y=11990 $D=193
M47 66 51 47 well_cntrl_res dgpfet L=2.4e-07 W=1.1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4870 $Y=11890 $D=193
M48 DVDD pu_en_tol_ 66 well_cntrl_res dgpfet L=2.4e-07 W=1.1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5570 $Y=11890 $D=193
M49 t3oR sdlow t3iR well_cntrl_res dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7410 $Y=9990 $D=193
M50 58 58 49 49 dgpfet L=1e-06 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7900 $Y=27560 $D=193
M51 t2oR sdlow t2iR well_cntrl_res dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9170 $Y=9990 $D=193
M52 psrc pctrl pgR well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10930 $Y=6990 $D=193
M53 pgR pctrl psrc well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11650 $Y=6990 $D=193
M54 psrc pctrl pgR well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12370 $Y=6990 $D=193
M55 pgR pctrl psrc well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=13090 $Y=6990 $D=193
M56 48 48 58 58 dgpfet L=2e-06 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=13610 $Y=28770 $D=193
M57 psrc pctrl pgL well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15890 $Y=6990 $D=193
M58 pgL pctrl psrc well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16610 $Y=6990 $D=193
M59 psrc pctrl pgL well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17330 $Y=6990 $D=193
M60 pgL pctrl psrc well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18050 $Y=6990 $D=193
M61 t2iL sdlow t2oL well_cntrl_res dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19810 $Y=9990 $D=193
M62 DVDD 58 54 DVDD dgpfet L=3e-07 W=1.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19970 $Y=26570 $D=193
M63 DVDD pg1 DVDD DVDD dgpfet L=2.4e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19970 $Y=29330 $D=193
M64 59 60 DVDD DVDD dgpfet L=2.4e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20950 $Y=26570 $D=193
M65 60 oeb_3v3 DVDD DVDD dgpfet L=2.4e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20950 $Y=28090 $D=193
M66 t3iL sdlow t3oL well_cntrl_res dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=21570 $Y=9990 $D=193
M67 61 54 59 DVDD dgpfet L=2.4e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=21870 $Y=26570 $D=193
M68 55 sdhigh 47 well_cntrl_res dgpfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=22060 $Y=6630 $D=193
M69 DVDD 61 n1_buf DVDD dgpfet L=2.4e-07 W=1.4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=22660 $Y=28150 $D=193
M70 62 n1_buf DVDD DVDD dgpfet L=2.4e-07 W=3.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23600 $Y=26570 $D=193
M71 67 47 DVDD well_cntrl_res dgpfet L=2.4e-07 W=6.4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23830 $Y=6630 $D=193
M72 pctrl plvl 67 well_cntrl_res dgpfet L=2.4e-07 W=6.4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=24370 $Y=6630 $D=193
M73 68 plvl pctrl well_cntrl_res dgpfet L=2.4e-07 W=6.4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=25070 $Y=6630 $D=193
M74 46 62 DVDD DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=25360 $Y=26570 $D=193
M75 DVDD 47 68 well_cntrl_res dgpfet L=2.4e-07 W=6.4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=25610 $Y=6630 $D=193
M76 DVDD 62 46 DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26060 $Y=26570 $D=193
M77 psupply 47 DVDD well_cntrl_res dgpfet L=2.4e-07 W=6.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26550 $Y=6230 $D=193
M78 46 62 DVDD DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26760 $Y=26570 $D=193
M79 DVDD 47 psupply well_cntrl_res dgpfet L=2.4e-07 W=6.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=27250 $Y=6230 $D=193
M80 psupply 47 DVDD well_cntrl_res dgpfet L=2.4e-07 W=6.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=27950 $Y=6230 $D=193
M81 DVDD 47 psupply well_cntrl_res dgpfet L=2.4e-07 W=6.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=28650 $Y=6230 $D=193
M82 psupply 47 DVDD well_cntrl_res dgpfet L=2.4e-07 W=6.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=29350 $Y=6230 $D=193
M83 47 46 pg1 well_cntrl_res dgpfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=31190 $Y=7030 $D=193
M84 pg0 46 47 well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=32150 $Y=8030 $D=193
M85 VDD alow 50 VDD dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=32720 $Y=24420 $D=193
M86 47 46 pg0 well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=32850 $Y=8030 $D=193
M87 pctrl 46 47 well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=33620 $Y=8030 $D=193
M88 47 46 pctrl well_cntrl_res dgpfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=34320 $Y=8030 $D=193
R89 52 DVDD 1000.61 L=8.42e-06 W=3e-06 sbar=1 m=1 par=1 bp=3 $SUB=VSS $[opppcres] $X=39720 $Y=6590 $D=355
D90 VSS 47 esdndsx areac=1.71799e-11 pjc=2.68627e-05 nf=1 bp=3 t3well=0 $X=42010 $Y=19800 $D=542
D91 VSS 47 esdndsx areac=1.71799e-11 pjc=2.68627e-05 nf=1 bp=3 t3well=0 $X=42010 $Y=24200 $D=542
X92 47 pad VSS ppoly_res_250 $T=50980 11940 0 270 $X=50680 $Y=7640
X93 pad 49 VSS ppoly_res_250 $T=55260 11940 0 270 $X=54960 $Y=7640
.ENDS
***************************************
.SUBCKT ICV_29 1 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25
** N=3052 EP=24 IP=45 FDC=94
X0 2 1 4 20 12 17 18 4 4 4 4 8 8 8 9 8 5 10 11 8
+ 9 4 4 11 5 9 8 8 10 9 5 6 19 23 25 7 13 14 15 16
+ 21 22 24
+ sc4 $T=0 0 0 0 $X=-5250 $Y=-2
.ENDS
***************************************
.SUBCKT ipplie DVSS pu pd ie oe y VDD VSS DVDD inxfr inp1 pd_en inn1 well_en_ pu_en_tol_ nctrl sdhigh oeb_3v3 psrc nsrc
+ n1_buf psupply pctrl alow sdlow puhi hic pdhi iehi oehi scmp scmn plvl nand nor
** N=3197 EP=35 IP=0 FDC=122
*.CALIBRE ISOLATED NETS: d
M0 inn1 inxfr VSS VSS dgnfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1980 $Y=16260 $D=106
M1 38 37 inn1 VSS dgnfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1300 $Y=16260 $D=106
M2 59 39 VSS VSS dgnfet L=2.4e-07 W=5.76e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1000 $Y=16260 $D=106
M3 VSS 39 59 VSS dgnfet L=2.4e-07 W=5.76e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1680 $Y=16260 $D=106
M4 60 38 scmn VSS dgnfet L=6.2e-07 W=4.86e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3580 $Y=16260 $D=106
M5 37 39 inxfr VSS dgnfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5860 $Y=16260 $D=106
M6 VSS VSS VSS VSS dgnfet L=6.2e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7460 $Y=21020 $D=106
M7 VSS 40 37 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7700 $Y=16260 $D=106
M8 41 38 VSS VSS dgnfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8660 $Y=16260 $D=106
M9 VSS 42 39 VSS dgnfet L=2.4e-07 W=8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12080 $Y=11540 $D=106
M10 40 iehi VSS VSS dgnfet L=2.4e-07 W=8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12760 $Y=11540 $D=106
M11 VSS 44 43 VSS dgnfet L=2.4e-07 W=4.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=14600 $Y=11540 $D=106
M12 45 sdhigh VSS VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15080 $Y=17020 $D=106
M13 61 puhi VSS VSS dgnfet L=2.4e-07 W=4.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15280 $Y=11540 $D=106
M14 VSS sdhigh 45 VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15760 $Y=17020 $D=106
M15 46 63 VSS VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16440 $Y=17020 $D=106
M16 VSS 53 pd_en VSS dgnfet L=2.4e-07 W=4.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17120 $Y=11540 $D=106
M17 VSS 63 46 VSS dgnfet L=2.4e-07 W=5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17120 $Y=17020 $D=106
M18 70 n1_buf VSS VSS dgnfet L=5e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18070 $Y=18960 $D=106
M19 62 pdhi VSS VSS dgnfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18080 $Y=11540 $D=106
M20 well_en_ 63 70 VSS dgnfet L=5e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18870 $Y=18960 $D=106
M21 66 48 VSS VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19920 $Y=11540 $D=106
M22 VSS 48 66 VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20600 $Y=11540 $D=106
M23 plvl 49 VSS VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=21280 $Y=11540 $D=106
M24 VSS 49 plvl VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=21960 $Y=11540 $D=106
M25 71 plvl pctrl VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23940 $Y=11540 $D=106
M26 VSS 64 71 VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=24480 $Y=11540 $D=106
M27 VSS 50 64 VSS dgnfet L=2.4e-07 W=5.66e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26320 $Y=11540 $D=106
M28 oeb_3v3 oehi VSS VSS dgnfet L=2.4e-07 W=8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=27280 $Y=11540 $D=106
M29 VSS 51 67 VSS dgnfet L=2.4e-07 W=8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=29120 $Y=11540 $D=106
M30 65 52 VSS VSS dgnfet L=2.4e-07 W=4.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30080 $Y=11540 $D=106
M31 DVSS 65 nctrl VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=31920 $Y=11540 $D=106
M32 DVSS 66 psrc VSS dgnfet L=2.4e-07 W=4.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=31920 $Y=17280 $D=106
M33 nsrc 67 DVSS VSS dgnfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=32880 $Y=11540 $D=106
M34 DVSS 67 nsrc VSS dgnfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=33560 $Y=11540 $D=106
M35 VSS 43 pu_en_tol_ VSS dgnfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=35400 $Y=11540 $D=106
M36 69 41 VSS VSS dgnfet L=2.4e-07 W=6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=59140 $Y=16260 $D=106
M37 58 38 69 VSS dgnfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=60100 $Y=16260 $D=106
M38 VSS puhi 44 VSS lpnfet w=1e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=41620 $Y=16260 $D=103
M39 pulow pu VSS VSS lpnfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=42460 $Y=16260 $D=103
M40 VSS pulow VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=42460 $Y=18440 $D=103
M41 VSS pdhi 53 VSS lpnfet w=1e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=44180 $Y=16260 $D=103
M42 pdlow pd VSS VSS lpnfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=45020 $Y=16260 $D=103
M43 VSS pdlow VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=45020 $Y=18440 $D=103
M44 VSS ie ielow VSS lpnfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=46740 $Y=16260 $D=103
M45 VSS ielow VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=46740 $Y=18660 $D=103
M46 42 iehi VSS VSS lpnfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=47560 $Y=16260 $D=103
M47 VSS oehi 50 VSS lpnfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=49300 $Y=16260 $D=103
M48 oelow oe VSS VSS lpnfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=50140 $Y=16260 $D=103
M49 VSS oelow VSS VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=50140 $Y=18660 $D=103
M50 VSS 51 52 VSS lpnfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=51860 $Y=16260 $D=103
M51 49 48 VSS VSS lpnfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=52700 $Y=16260 $D=103
M52 72 nand 48 VSS lpnfet w=1e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=54440 $Y=16260 $D=103
M53 VSS oehi 72 VSS lpnfet w=1e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=54840 $Y=16260 $D=103
M54 51 nor VSS VSS lpnfet w=4e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=56000 $Y=16260 $D=103
M55 VSS 68 51 VSS lpnfet w=4e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=56580 $Y=16260 $D=103
M56 68 oehi VSS VSS lpnfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=57420 $Y=16260 $D=103
M57 y 69 VSS VSS lpnfet w=5.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=61980 $Y=16260 $D=103
M58 VSS 69 y VSS lpnfet w=5.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=62540 $Y=16260 $D=103
M59 psupply inxfr inp1 DVDD dgpfet L=2.4e-07 W=8.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-2660 $Y=4320 $D=193
M60 inp1 inxfr psupply DVDD dgpfet L=2.4e-07 W=8.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1980 $Y=4320 $D=193
M61 38 inxfr inp1 DVDD dgpfet L=2.4e-07 W=8.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-1300 $Y=4320 $D=193
M62 inp1 inxfr 38 DVDD dgpfet L=2.4e-07 W=8.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=-620 $Y=4320 $D=193
M63 59 38 scmp DVDD dgpfet L=3.8e-07 W=5.76e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1220 $Y=7060 $D=193
M64 scmp 38 59 DVDD dgpfet L=3.8e-07 W=5.76e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2040 $Y=7060 $D=193
M65 60 40 DVDD DVDD dgpfet L=2.4e-07 W=4.86e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4020 $Y=7960 $D=193
M66 37 40 inxfr DVDD dgpfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5860 $Y=8820 $D=193
M67 DVDD DVDD DVDD DVDD dgpfet L=3.8e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6360 $Y=7060 $D=193
M68 41 38 DVDD DVDD dgpfet L=2.4e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7700 $Y=8800 $D=193
M69 DVDD 39 38 DVDD dgpfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7700 $Y=10820 $D=193
M70 DVDD 40 39 DVDD dgpfet L=2.4e-07 W=3.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12080 $Y=4900 $D=193
M71 40 39 DVDD DVDD dgpfet L=2.4e-07 W=3.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12760 $Y=4900 $D=193
M72 DVDD 61 43 DVDD dgpfet L=2.4e-07 W=1.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=14600 $Y=6300 $D=193
M73 61 43 DVDD DVDD dgpfet L=2.4e-07 W=1.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15280 $Y=6300 $D=193
M74 sdhigh 47 DVDD DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=15560 $Y=1840 $D=193
M75 DVDD 47 sdhigh DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16240 $Y=1840 $D=193
M76 sdhigh 47 DVDD DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16920 $Y=1840 $D=193
M77 DVDD 62 pd_en DVDD dgpfet L=2.4e-07 W=1.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17120 $Y=6300 $D=193
M78 DVDD 47 sdhigh DVDD dgpfet L=2.4e-07 W=2.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=17600 $Y=1840 $D=193
M79 62 pd_en DVDD DVDD dgpfet L=2.4e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18080 $Y=7100 $D=193
M80 63 47 DVDD DVDD dgpfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=18560 $Y=1840 $D=193
M81 DVDD 47 63 DVDD dgpfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19240 $Y=1840 $D=193
M82 DVDD plvl 66 DVDD dgpfet L=2.4e-07 W=3.6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=19920 $Y=4500 $D=193
M83 plvl 66 DVDD DVDD dgpfet L=2.4e-07 W=3.6e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=20600 $Y=4500 $D=193
M84 psrc 66 DVDD DVDD dgpfet L=2.4e-07 W=6.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=22440 $Y=1840 $D=193
M85 DVDD 66 psrc DVDD dgpfet L=2.4e-07 W=6.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23120 $Y=1840 $D=193
M86 psrc 66 DVDD DVDD dgpfet L=2.4e-07 W=6.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=23800 $Y=1840 $D=193
M87 DVDD 66 psrc DVDD dgpfet L=2.4e-07 W=6.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=24480 $Y=1840 $D=193
M88 DVDD oeb_3v3 64 DVDD dgpfet L=2.4e-07 W=2.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=26320 $Y=5840 $D=193
M89 oeb_3v3 64 DVDD DVDD dgpfet L=2.4e-07 W=3.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=27280 $Y=4900 $D=193
M90 DVDD 65 67 DVDD dgpfet L=2.4e-07 W=3.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=29120 $Y=4900 $D=193
M91 65 67 DVDD DVDD dgpfet L=2.4e-07 W=1.8e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30080 $Y=6300 $D=193
M92 DVDD 65 nctrl DVDD dgpfet L=2.4e-07 W=4.5e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=31920 $Y=3600 $D=193
M93 nsrc nctrl DVDD DVDD dgpfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=32880 $Y=4100 $D=193
M94 DVDD nctrl nsrc DVDD dgpfet L=2.4e-07 W=4e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=33560 $Y=4100 $D=193
M95 pu_en_tol_ 43 DVDD DVDD dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=34520 $Y=5100 $D=193
M96 69 41 VDD VDD dgpfet L=2.4e-07 W=3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=59140 $Y=9820 $D=193
M97 VDD 47 hic VDD lppfet w=4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=39900 $Y=8820 $D=192
M98 VDD puhi 44 VDD lppfet w=3e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=41620 $Y=9820 $D=192
M99 pulow pu VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=42460 $Y=9820 $D=192
M100 VDD pdhi 53 VDD lppfet w=3e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=44180 $Y=9820 $D=192
M101 pdlow pd VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=45020 $Y=9820 $D=192
M102 VDD ie ielow VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=46740 $Y=9820 $D=192
M103 42 iehi VDD VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=47560 $Y=7820 $D=192
M104 VDD iehi 42 VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=48140 $Y=7820 $D=192
M105 50 oehi VDD VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=48720 $Y=7820 $D=192
M106 VDD oehi 50 VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=49300 $Y=7820 $D=192
M107 oelow oe VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=50140 $Y=9820 $D=192
M108 VDD 51 52 VDD lppfet w=4e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=51860 $Y=8820 $D=192
M109 49 48 VDD VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=52700 $Y=7820 $D=192
M110 VDD 48 49 VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=53280 $Y=7820 $D=192
M111 48 nand VDD VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=53860 $Y=7820 $D=192
M112 VDD oehi 48 VDD lppfet w=5e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=54440 $Y=7820 $D=192
M113 73 nor 51 VDD lppfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=56180 $Y=10820 $D=192
M114 VDD 68 73 VDD lppfet w=2e-06 l=1.4e-07 m=1 par=1 nf=1 ngcon=1 $X=56580 $Y=10820 $D=192
M115 68 oehi VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=57420 $Y=9820 $D=192
M116 VDD alow 58 VDD lppfet w=7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=61160 $Y=5820 $D=192
M117 y 69 VDD VDD lppfet w=7.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=61980 $Y=5620 $D=192
M118 VDD 69 y VDD lppfet w=7.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=62540 $Y=5620 $D=192
R119 47 VSS 1000.61 L=8.42e-06 W=3e-06 sbar=1 m=1 par=1 bp=3 $SUB=VSS $[opppcres] $X=35870 $Y=19640 $D=355
R120 sdlow 45 1000.61 L=8.42e-06 W=3e-06 sbar=1 m=1 par=1 bp=3 $SUB=VSS $[opppcres] $X=39210 $Y=2660 $D=355
R121 alow 46 1000.61 L=8.42e-06 W=3e-06 sbar=1 m=1 par=1 bp=3 $SUB=VSS $[opppcres] $X=49410 $Y=2660 $D=355
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21
** N=1800 EP=21 IP=36 FDC=122
X0 1 4 4 5 4 6 2 3 8 20 22 9 23 10 11 12 17 13 14 15
+ 16 18 21 4 7 4 24 4 5 4 22 23 19 4 24
+ ipplie $T=5000 223260 0 0 $X=180 $Y=223260
.ENDS
***************************************
.SUBCKT MVNSX_1AS_ARTI 1 2
** N=1248 EP=2 IP=0 FDC=5
D0 2 1 esdndsx areac=7.1024e-11 pjc=0.000103783 nf=1 bp=3 t3well=0 $X=4000 $Y=3360 $D=542
D1 2 1 esdndsx areac=7.1024e-11 pjc=0.000103783 nf=1 bp=3 t3well=0 $X=8400 $Y=3360 $D=542
D2 2 1 esdndsx areac=7.1024e-11 pjc=0.000103783 nf=1 bp=3 t3well=0 $X=12800 $Y=3360 $D=542
D3 2 1 esdndsx areac=7.1024e-11 pjc=0.000103783 nf=1 bp=3 t3well=0 $X=17200 $Y=3360 $D=542
D4 2 1 esdndsx areac=7.1024e-11 pjc=0.000103783 nf=1 bp=3 t3well=0 $X=21600 $Y=3360 $D=542
.ENDS
***************************************
.SUBCKT MSVSXBAR_B
** N=331 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MSVSXBAR_A
** N=253 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MVBIT5_1AS_ARTI
** N=358 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT bp_i pad VSS
** N=3523 EP=2 IP=13 FDC=5
*.CALIBRE ISOLATED NETS: DVDD
X0 pad VSS MVNSX_1AS_ARTI $T=64980 89040 1 270 $X=5020 $Y=54020
.ENDS
***************************************
.SUBCKT ICV_38 1 3
** N=3 EP=2 IP=3 FDC=5
X0 1 3 bp_i $T=0 0 0 0 $X=-140 $Y=0
.ENDS
***************************************
.SUBCKT pct_capl
** N=661 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVSS VSS ng1 ng0 DVDD sdlow poff pg1 pg0 well_cntrl_res
.ENDS
***************************************
.SUBCKT ICV_37
** N=145 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT pct pad DVDD ptr0m2 ptr1m2 well_cntrl_res
** N=264 EP=5 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: poff pg0 pg1
M0 pad ptr0m2 DVDD well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=620 $D=193
M1 DVDD ptr1m2 pad well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9380 $Y=620 $D=193
.ENDS
***************************************
.SUBCKT ICV_36 1 3 4 5 7
** N=415 EP=5 IP=11 FDC=2
X0 3 1 4 5 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT pct2 pad DVDD ptr0m2 ptr1m2 well_cntrl_res
** N=262 EP=5 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: pg0 pg1 poff
M0 pad ptr0m2 DVDD well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=620 $D=193
M1 DVDD ptr1m2 pad well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9380 $Y=620 $D=193
.ENDS
***************************************
.SUBCKT ICV_35 1 3 4 7
** N=449 EP=4 IP=9 FDC=2
X0 3 1 4 4 7 pct2 $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT pct2_tap pad DVDD ptr0m2 well_cntrl_res ptr1m2
** N=426 EP=5 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: pg0 pg1 poff
M0 pad ptr0m2 DVDD well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=620 $D=193
M1 DVDD ptr1m2 pad well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9380 $Y=620 $D=193
.ENDS
***************************************
.SUBCKT ICV_34 1 3 4 6
** N=415 EP=4 IP=9 FDC=2
X0 3 1 4 6 4 pct2_tap $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_33 1 3 4 7
** N=449 EP=4 IP=11 FDC=2
X0 3 1 4 4 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT pct_tap pad DVDD ptr0m2 well_cntrl_res ptr1m2
** N=426 EP=5 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: poff pg0 pg1
M0 pad ptr0m2 DVDD well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=620 $D=193
M1 DVDD ptr1m2 pad well_cntrl_res dgpfet L=2.4e-07 W=3.544e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9380 $Y=620 $D=193
.ENDS
***************************************
.SUBCKT ICV_32 1 3 4 5
** N=415 EP=4 IP=9 FDC=2
X0 3 1 4 5 4 pct_tap $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_31 1 3 4 7
** N=483 EP=4 IP=11 FDC=2
X0 3 1 4 4 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT pct_capr
** N=660 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVDD ng0 ng1 VSS pg0 pg1 sdhigh poff well_cntrl_res
.ENDS
***************************************
.SUBCKT ICV_30
** N=247 EP=0 IP=9 FDC=0
.ENDS
***************************************
.SUBCKT PICS DVSS VSS DVDD VDD IE Y P
** N=27 EP=7 IP=120 FDC=269
X0 DVSS 8 9 P 13 ICV_40 $T=0 0 0 0 $X=-250 $Y=117000
X1 VSS DVDD 8 9 13 P 11 12 19 20 10 14 15 16 17 18 21 22 23 24
+ 25 26 27 VDD
+ ICV_29 $T=5000 192280 0 0 $X=-250 $Y=192278
X2 DVSS VDD VSS 27 IE Y 8 DVDD 14 15 16 17 18 19 20 21 13 22 24 25
+ 26
+ ICV_39 $T=0 0 0 0 $X=-250 $Y=223260
X3 P VSS ICV_38 $T=0 0 0 0 $X=-140 $Y=0
X5 DVDD P 11 10 23 ICV_36 $T=5000 151580 0 0 $X=3020 $Y=151300
X6 DVDD P 10 23 ICV_35 $T=15000 151580 0 0 $X=13020 $Y=151300
X7 DVDD P 10 23 ICV_34 $T=25000 151580 0 0 $X=23020 $Y=151300
X8 DVDD P 10 23 ICV_33 $T=35000 151580 0 0 $X=33020 $Y=151300
X9 DVDD P 10 23 ICV_32 $T=45000 151580 0 0 $X=43020 $Y=151300
X10 DVDD P 10 23 ICV_31 $T=55000 151580 0 0 $X=53020 $Y=151300
.ENDS
***************************************
.SUBCKT vddbp_i 1 VSS 4
** N=2305 EP=3 IP=32 FDC=24
X0 15 9 10 16 4 VSS ICV_152 $T=33550 79300 0 90 $X=7070 $Y=78980
X1 21 26 27 22 1 VSS ICV_152 $T=36450 79300 1 90 $X=36150 $Y=78980
X2 11 5 6 12 7 13 8 14 9 VSS ICV_153 $T=33550 56900 0 90 $X=7070 $Y=56580
X3 17 5 23 18 24 19 25 20 26 VSS ICV_153 $T=36450 56900 1 90 $X=36150 $Y=56580
.ENDS
***************************************
.SUBCKT ipplscp_vdd VSS VDD 5
** N=17055 EP=3 IP=0 FDC=196
*.CALIBRE ISOLATED NETS: DVSS DVDD
M0 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=5370 $D=106
M1 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=6050 $D=106
M2 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=6730 $D=106
M3 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=7410 $D=106
M4 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=8090 $D=106
M5 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=8770 $D=106
M6 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=9450 $D=106
M7 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=10130 $D=106
M8 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=10810 $D=106
M9 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=11490 $D=106
M10 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=12170 $D=106
M11 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=12850 $D=106
M12 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=13530 $D=106
M13 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=14210 $D=106
M14 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=14890 $D=106
M15 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=17910 $D=106
M16 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=18590 $D=106
M17 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=19270 $D=106
M18 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=19950 $D=106
M19 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=20630 $D=106
M20 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=21310 $D=106
M21 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=21990 $D=106
M22 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=22670 $D=106
M23 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=23350 $D=106
M24 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=24030 $D=106
M25 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=24710 $D=106
M26 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=25390 $D=106
M27 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=26070 $D=106
M28 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=26750 $D=106
M29 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=27430 $D=106
M30 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=30450 $D=106
M31 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=31130 $D=106
M32 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=31810 $D=106
M33 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=32490 $D=106
M34 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=33170 $D=106
M35 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=33850 $D=106
M36 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=34530 $D=106
M37 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=35210 $D=106
M38 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=35890 $D=106
M39 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=36570 $D=106
M40 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=37250 $D=106
M41 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=37930 $D=106
M42 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=38610 $D=106
M43 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=39290 $D=106
M44 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=39970 $D=106
M45 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=42990 $D=106
M46 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=43670 $D=106
M47 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=44350 $D=106
M48 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=45030 $D=106
M49 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=45710 $D=106
M50 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=46390 $D=106
M51 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=47070 $D=106
M52 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=47750 $D=106
M53 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=48430 $D=106
M54 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=49110 $D=106
M55 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=49790 $D=106
M56 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=50470 $D=106
M57 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=51150 $D=106
M58 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=51830 $D=106
M59 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=52510 $D=106
M60 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=55530 $D=106
M61 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=56210 $D=106
M62 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=56890 $D=106
M63 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=57570 $D=106
M64 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=58250 $D=106
M65 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=58930 $D=106
M66 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=59610 $D=106
M67 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=60290 $D=106
M68 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=60970 $D=106
M69 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=61650 $D=106
M70 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=62330 $D=106
M71 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=63010 $D=106
M72 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=63690 $D=106
M73 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=64370 $D=106
M74 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4810 $Y=65050 $D=106
M75 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=68810 $D=106
M76 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=69490 $D=106
M77 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=70170 $D=106
M78 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=30220 $Y=70850 $D=106
M79 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=5370 $D=106
M80 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=6050 $D=106
M81 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=6730 $D=106
M82 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=7410 $D=106
M83 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=8090 $D=106
M84 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=8770 $D=106
M85 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=9450 $D=106
M86 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=10130 $D=106
M87 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=10810 $D=106
M88 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=11490 $D=106
M89 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=12170 $D=106
M90 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=12850 $D=106
M91 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=13530 $D=106
M92 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=14210 $D=106
M93 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=14890 $D=106
M94 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=17910 $D=106
M95 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=18590 $D=106
M96 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=19270 $D=106
M97 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=19950 $D=106
M98 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=20630 $D=106
M99 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=21310 $D=106
M100 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=21990 $D=106
M101 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=22670 $D=106
M102 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=23350 $D=106
M103 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=24030 $D=106
M104 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=24710 $D=106
M105 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=25390 $D=106
M106 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=26070 $D=106
M107 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=26750 $D=106
M108 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=27430 $D=106
M109 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=30450 $D=106
M110 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=31130 $D=106
M111 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=31810 $D=106
M112 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=32490 $D=106
M113 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=33170 $D=106
M114 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=33850 $D=106
M115 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=34530 $D=106
M116 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=35210 $D=106
M117 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=35890 $D=106
M118 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=36570 $D=106
M119 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=37250 $D=106
M120 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=37930 $D=106
M121 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=38610 $D=106
M122 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=39290 $D=106
M123 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=39970 $D=106
M124 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=42990 $D=106
M125 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=43670 $D=106
M126 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=44350 $D=106
M127 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=45030 $D=106
M128 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=45710 $D=106
M129 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=46390 $D=106
M130 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=47070 $D=106
M131 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=47750 $D=106
M132 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=48430 $D=106
M133 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=49110 $D=106
M134 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=49790 $D=106
M135 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=50470 $D=106
M136 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=51150 $D=106
M137 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=51830 $D=106
M138 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=52510 $D=106
M139 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=55530 $D=106
M140 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=56210 $D=106
M141 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=56890 $D=106
M142 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=57570 $D=106
M143 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=58250 $D=106
M144 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=58930 $D=106
M145 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=59610 $D=106
M146 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=60290 $D=106
M147 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=60970 $D=106
M148 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=61650 $D=106
M149 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=62330 $D=106
M150 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=63010 $D=106
M151 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=63690 $D=106
M152 VSS 6 VDD VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=64370 $D=106
M153 VDD 6 VSS VSS dgnfet L=2.4e-07 W=2.9e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=36190 $Y=65050 $D=106
M154 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=68810 $D=106
M155 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=69490 $D=106
M156 6 5 VSS VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=70170 $D=106
M157 VSS 5 6 VSS dgnfet L=2.4e-07 W=2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=37780 $Y=70850 $D=106
M158 6 5 VDD VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=68810 $D=193
M159 VDD 5 6 VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=69490 $D=193
M160 6 5 VDD VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=70170 $D=193
M161 VDD 5 6 VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=16940 $Y=70850 $D=193
M162 6 5 VDD VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=68810 $D=193
M163 VDD 5 6 VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=69490 $D=193
M164 6 5 VDD VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=70170 $D=193
M165 VDD 5 6 VDD dgpfet L=2.4e-07 W=1e-05 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43060 $Y=70850 $D=193
X166 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=76490 $D=397
X167 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=84470 $D=397
X168 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=92450 $D=397
X169 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=100430 $D=397
X170 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=108410 $D=397
X171 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=8560 $Y=116390 $D=397
X172 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=76490 $D=397
X173 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=84470 $D=397
X174 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=92450 $D=397
X175 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=100430 $D=397
X176 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=108410 $D=397
X177 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=19280 $Y=116390 $D=397
X178 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=76490 $D=397
X179 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=84470 $D=397
X180 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=92450 $D=397
X181 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=100430 $D=397
X182 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=108410 $D=397
X183 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=30000 $Y=116390 $D=397
X184 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=76490 $D=397
X185 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=84470 $D=397
X186 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=92450 $D=397
X187 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=100430 $D=397
X188 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=108410 $D=397
X189 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=40720 $Y=116390 $D=397
X190 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=76490 $D=397
X191 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=84470 $D=397
X192 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=92450 $D=397
X193 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=100430 $D=397
X194 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=108410 $D=397
X195 5 VSS VSS VSS dgncap w=1e-05 l=7.5e-06 m=1 pcrep=1 prxrep=1 $X=51440 $Y=116390 $D=397
.ENDS
***************************************
.SUBCKT ICV_165
** N=1220 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_164
** N=1409 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_163
** N=1570 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_162
** N=1394 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_161
** N=785 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_160
** N=1576 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_159
** N=1309 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_158
** N=1343 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT vdd_oly
** N=4 EP=0 IP=19 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS VDD DVSS
.ENDS
***************************************
.SUBCKT PVDD VSS DVSS DVDD VDD
** N=5 EP=4 IP=13 FDC=220
X0 VDD VSS 5 vddbp_i $T=0 0 0 0 $X=-140 $Y=0
X1 VSS VDD 5 ipplscp_vdd $T=0 117000 0 0 $X=-140 $Y=117000
.ENDS
***************************************
.SUBCKT vssbp_i
** N=1719 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: DVDD
.ENDS
***************************************
.SUBCKT ICV_173
** N=2104 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_172
** N=2291 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_171
** N=2162 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_170
** N=1394 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_169
** N=786 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_168
** N=2606 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_167
** N=1309 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_166
** N=1583 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT vss_oly
** N=92 EP=0 IP=200 FDC=0
*.CALIBRE ISOLATED NETS: DVDD VSS VDD DVSS
.ENDS
***************************************
.SUBCKT ipplscp_vss_sub
** N=1534 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ipplscp_vss
** N=4506 EP=0 IP=2460 FDC=0
*.CALIBRE ISOLATED NETS: VSS DVDD DVSS
.ENDS
***************************************
.SUBCKT PVSS VSS DVSS DVDD VDD
** N=4 EP=4 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_260 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=106 FDC=978
X9 1 2 3 4 PDVDD $T=845000 0 0 180 $X=774860 $Y=-247000
X20 1 2 3 4 PDVSS $T=920000 0 0 180 $X=849860 $Y=-247000
X21 2 1 3 4 4 6 5 PICS $T=995000 0 0 180 $X=924760 $Y=-247002
X22 2 1 3 4 4 8 7 PICS $T=1070000 0 0 180 $X=999760 $Y=-247002
X23 1 2 3 4 PVDD $T=1145000 0 0 180 $X=1074860 $Y=-247000
X24 1 2 3 4 PVSS $T=1220000 0 0 180 $X=1149860 $Y=-247000
.ENDS
***************************************
.SUBCKT ICV_259
** N=4 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_258
** N=4 EP=0 IP=32 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_257
** N=4 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_150
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_242
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_254 2 5 6 7 12
** N=2721 EP=5 IP=179 FDC=36
X3 2 7 6 5 12 13 14 nct $T=5000 121510 0 0 $X=3420 $Y=121360
X4 2 7 6 5 12 15 16 nct $T=15000 121510 0 0 $X=13420 $Y=121360
X5 2 7 6 5 12 17 18 nct $T=25000 121510 0 0 $X=23420 $Y=121360
X6 2 7 6 5 12 19 20 nct $T=35000 121510 0 0 $X=33420 $Y=121360
X7 2 7 6 5 12 21 22 nct $T=45000 121510 0 0 $X=43420 $Y=121360
X8 2 7 6 5 12 23 24 nct $T=55000 121510 0 0 $X=53420 $Y=121360
.ENDS
***************************************
.SUBCKT ICV_243 1 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26
** N=3053 EP=25 IP=45 FDC=94
X0 2 1 4 21 13 18 19 5 5 6 5 10 10 9 9 10 5 11 12 10
+ 9 6 6 12 6 9 9 9 11 9 6 7 20 24 26 8 14 15 16 17
+ 22 23 25
+ sc4 $T=0 0 0 0 $X=-5250 $Y=-2
.ENDS
***************************************
.SUBCKT ICV_253 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
** N=1800 EP=20 IP=36 FDC=122
X0 1 4 4 4 21 22 2 3 7 19 23 8 24 9 10 11 16 12 13 14
+ 15 17 20 4 6 4 21 4 4 21 3 7 18 5 5
+ ipplie $T=5000 223260 0 0 $X=180 $Y=223260
.ENDS
***************************************
.SUBCKT ICV_252 1 3
** N=3 EP=2 IP=3 FDC=5
X0 1 3 bp_i $T=0 0 0 0 $X=-140 $Y=0
.ENDS
***************************************
.SUBCKT ICV_251
** N=146 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_250 1 3 4 5 7
** N=415 EP=5 IP=11 FDC=2
X0 3 1 4 5 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_249 1 3 4 5 7
** N=449 EP=5 IP=9 FDC=2
X0 3 1 4 5 7 pct2 $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_248 1 3 4 5 6
** N=415 EP=5 IP=9 FDC=2
X0 3 1 4 5 6 pct2_tap $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_247 1 3 4 5 7
** N=449 EP=5 IP=11 FDC=2
X0 3 1 4 5 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_246 1 3 4 5 6
** N=415 EP=5 IP=9 FDC=2
X0 3 1 4 5 6 pct_tap $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_245 1 3 4 5 7
** N=483 EP=5 IP=11 FDC=2
X0 3 1 4 5 7 pct $T=0 0 0 0 $X=-1980 $Y=-280
.ENDS
***************************************
.SUBCKT ICV_244
** N=247 EP=0 IP=9 FDC=0
.ENDS
***************************************
.SUBCKT POC24A DVSS VSS DVDD VDD P A
** N=27 EP=6 IP=122 FDC=269
X0 DVSS 7 8 P 13 ICV_254 $T=0 0 0 0 $X=-250 $Y=117000
X1 VSS DVDD 9 7 8 13 P 12 11 19 20 10 14 15 16 17 18 21 22 23
+ 24 25 26 27 VDD
+ ICV_243 $T=5000 192280 0 0 $X=-250 $Y=192278
X2 DVSS VDD VSS 27 A 9 DVDD 14 15 16 17 18 19 20 21 13 22 24 25 26 ICV_253 $T=0 0 0 0 $X=-250 $Y=223260
X3 P VSS ICV_252 $T=0 0 0 0 $X=-140 $Y=0
X5 DVDD P 12 11 23 ICV_250 $T=5000 151580 0 0 $X=3020 $Y=151300
X6 DVDD P 12 11 23 ICV_249 $T=15000 151580 0 0 $X=13020 $Y=151300
X7 DVDD P 12 23 11 ICV_248 $T=25000 151580 0 0 $X=23020 $Y=151300
X8 DVDD P 12 11 23 ICV_247 $T=35000 151580 0 0 $X=33020 $Y=151300
X9 DVDD P 12 23 11 ICV_246 $T=45000 151580 0 0 $X=43020 $Y=151300
X10 DVDD P 12 11 23 ICV_245 $T=55000 151580 0 0 $X=53020 $Y=151300
.ENDS
***************************************
.SUBCKT ICV_255 1 2 3 4 5 6
** N=6 EP=6 IP=14 FDC=269
X2 2 1 3 4 5 6 POC24A $T=5000 0 0 0 $X=4750 $Y=0
.ENDS
***************************************
.SUBCKT ICV_256 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
** N=37 EP=36 IP=140 FDC=4744
X3 1 2 3 4 PDVDD $T=1605000 0 0 0 $X=1604860 $Y=0
X4 1 2 3 4 PVDD $T=255000 0 0 0 $X=254860 $Y=0
X5 1 2 3 4 PVSS $T=330000 0 0 0 $X=329860 $Y=0
X11 1 2 3 4 5 21 ICV_255 $T=400000 0 0 0 $X=399860 $Y=0
X12 1 2 3 4 6 22 ICV_255 $T=475000 0 0 0 $X=474860 $Y=0
X13 1 2 3 4 7 23 ICV_255 $T=550000 0 0 0 $X=549860 $Y=0
X14 1 2 3 4 8 24 ICV_255 $T=625000 0 0 0 $X=624860 $Y=0
X15 1 2 3 4 9 25 ICV_255 $T=700000 0 0 0 $X=699860 $Y=0
X16 1 2 3 4 10 26 ICV_255 $T=775000 0 0 0 $X=774860 $Y=0
X17 1 2 3 4 11 27 ICV_255 $T=850000 0 0 0 $X=849860 $Y=0
X18 1 2 3 4 12 28 ICV_255 $T=925000 0 0 0 $X=924860 $Y=0
X19 1 2 3 4 13 29 ICV_255 $T=1000000 0 0 0 $X=999860 $Y=0
X20 1 2 3 4 14 30 ICV_255 $T=1075000 0 0 0 $X=1074860 $Y=0
X21 1 2 3 4 15 31 ICV_255 $T=1150000 0 0 0 $X=1149860 $Y=0
X22 1 2 3 4 16 32 ICV_255 $T=1225000 0 0 0 $X=1224860 $Y=0
X23 1 2 3 4 17 33 ICV_255 $T=1300000 0 0 0 $X=1299860 $Y=0
X24 1 2 3 4 18 34 ICV_255 $T=1375000 0 0 0 $X=1374860 $Y=0
X25 1 2 3 4 19 35 ICV_255 $T=1450000 0 0 0 $X=1449860 $Y=0
X26 1 2 3 4 20 36 ICV_255 $T=1525000 0 0 0 $X=1524860 $Y=0
.ENDS
***************************************
.SUBCKT ICV_177
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_178
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_179 1 2 202 203 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857
** N=11136 EP=34 IP=217 FDC=4475
X3 1 202 203 2 PDVDD $T=345000 2000000 0 180 $X=274860 $Y=1753000
X5 1 202 203 2 PDVSS $T=420000 2000000 0 180 $X=349860 $Y=1753000
X6 202 1 203 2 2 829 828 PICS $T=495000 2000000 0 180 $X=424760 $Y=1752998
X7 202 1 203 2 2 831 830 PICS $T=570000 2000000 0 180 $X=499760 $Y=1752998
X8 202 1 203 2 2 833 832 PICS $T=645000 2000000 0 180 $X=574760 $Y=1752998
X9 202 1 203 2 2 835 834 PICS $T=720000 2000000 0 180 $X=649760 $Y=1752998
X10 202 1 203 2 2 837 836 PICS $T=795000 2000000 0 180 $X=724760 $Y=1752998
X11 202 1 203 2 2 839 838 PICS $T=870000 2000000 0 180 $X=799760 $Y=1752998
X12 202 1 203 2 2 841 840 PICS $T=945000 2000000 0 180 $X=874760 $Y=1752998
X13 202 1 203 2 2 843 842 PICS $T=1020000 2000000 0 180 $X=949760 $Y=1752998
X14 202 1 203 2 2 845 844 PICS $T=1095000 2000000 0 180 $X=1024760 $Y=1752998
X15 202 1 203 2 2 847 846 PICS $T=1170000 2000000 0 180 $X=1099760 $Y=1752998
X16 202 1 203 2 2 849 848 PICS $T=1245000 2000000 0 180 $X=1174760 $Y=1752998
X17 202 1 203 2 2 851 850 PICS $T=1320000 2000000 0 180 $X=1249760 $Y=1752998
X18 202 1 203 2 2 853 852 PICS $T=1395000 2000000 0 180 $X=1324760 $Y=1752998
X19 202 1 203 2 2 855 854 PICS $T=1470000 2000000 0 180 $X=1399760 $Y=1752998
X20 202 1 203 2 2 857 856 PICS $T=1545000 2000000 0 180 $X=1474760 $Y=1752998
X21 1 202 203 2 PVDD $T=1620000 2000000 0 180 $X=1549860 $Y=1753000
X22 1 202 203 2 PVSS $T=1695000 2000000 0 180 $X=1624860 $Y=1753000
.ENDS
***************************************
.SUBCKT FILL64TR
** N=148 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_182
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_189
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_198
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_199
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_200
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_190
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_191
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_193
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_194
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_240
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_183
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT FILL32TR
** N=74 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL4TR
** N=8 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL1TR
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_185
** N=2 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_236
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_237
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_238
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_241
** N=113979 EP=0 IP=104 FDC=0
.ENDS
***************************************
.SUBCKT ICV_201
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_195
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_196
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT FILL2TR
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT CLKBUFX2TR A VSS VDD Y
** N=18 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1110 $D=97
M1 Y 5 VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=830 $D=97
M2 VDD A 5 VDD pfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=580 $Y=1910 $D=189
M3 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1070 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT FILL16TR
** N=36 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL8TR
** N=18 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_239 1 2 1017 1383
** N=206627 EP=4 IP=124 FDC=4
X58 1017 1 2 1383 CLKBUFX2TR $T=1518600 547400 1 0 $X=1518260 $Y=543400
.ENDS
***************************************
.SUBCKT ICV_220
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX8TR A Y VDD VSS
** N=32 EP=4 IP=0 FDC=8
M0 Y A VSS VSS nfet L=1.2e-07 W=5.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=720 $D=97
M1 VSS A Y VSS nfet L=1.2e-07 W=5.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=930 $Y=720 $D=97
M2 Y A VSS VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1490 $Y=790 $D=97
M3 VSS A Y VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=790 $D=97
M4 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=1910 $D=189
M5 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=930 $Y=1910 $D=189
M6 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1410 $Y=1910 $D=189
M7 VDD A Y VDD pfet L=1.2e-07 W=1.16e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1890 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_226
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX20TR A Y VSS VDD
** N=54 EP=4 IP=0 FDC=20
M0 Y A VSS VSS nfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=700 $D=97
M1 VSS A Y VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=900 $Y=540 $D=97
M2 Y A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1380 $Y=540 $D=97
M3 VSS A Y VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1860 $Y=540 $D=97
M4 Y A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2340 $Y=540 $D=97
M5 VSS A Y VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2820 $Y=540 $D=97
M6 Y A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3300 $Y=540 $D=97
M7 VSS A Y VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3780 $Y=540 $D=97
M8 Y A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4260 $Y=540 $D=97
M9 VSS A Y VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4740 $Y=680 $D=97
M10 Y A VDD VDD pfet L=1.2e-07 W=1.04e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M11 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=900 $Y=1910 $D=189
M12 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1380 $Y=1910 $D=189
M13 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1860 $Y=1910 $D=189
M14 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2340 $Y=1910 $D=189
M15 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2820 $Y=1910 $D=189
M16 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3300 $Y=1910 $D=189
M17 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3780 $Y=1910 $D=189
M18 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4260 $Y=1910 $D=189
M19 VDD A Y VDD pfet L=1.2e-07 W=1.06e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4740 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_222
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_188
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_206
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_203
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_216
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_181
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_225
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_223
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_234
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT INVX1TR VSS VDD A Y
** N=14 EP=4 IP=0 FDC=2
M0 Y A VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=520 $Y=850 $D=97
M1 Y A VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=520 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_180
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT AND2X2TR A B VDD VSS Y
** N=26 EP=5 IP=0 FDC=6
M0 7 A 6 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=470 $Y=830 $D=97
M1 VSS B 7 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=810 $Y=830 $D=97
M2 Y 6 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=390 $D=97
M3 6 A VDD VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=470 $Y=1910 $D=189
M4 VDD B 6 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=910 $Y=1910 $D=189
M5 Y 6 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_211
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT DLY3X1TR A VSS VDD Y
** N=43 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=790 $D=97
M1 6 5 VSS VSS nfet L=4.4e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1020 $Y=790 $D=97
M2 VSS 6 7 VSS nfet L=4.4e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=780 $D=97
M3 Y 7 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1060 $D=97
M4 VDD A 5 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M5 6 5 VDD VDD pfet L=4.4e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1020 $Y=1910 $D=189
M6 VDD 6 7 VDD pfet L=4.4e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=1910 $D=189
M7 Y 7 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DLY2X1TR A VSS VDD Y
** N=43 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1070 $D=97
M1 6 5 VSS VSS nfet L=2.4e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1220 $Y=790 $D=97
M2 VSS 6 7 VSS nfet L=2.4e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=780 $D=97
M3 Y 7 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1060 $D=97
M4 VDD A 5 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M5 6 5 VDD VDD pfet L=2.4e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1220 $Y=1910 $D=189
M6 VDD 6 7 VDD pfet L=2.4e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=1910 $D=189
M7 Y 7 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DLY1X1TR A VSS VDD Y
** N=43 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=790 $D=97
M1 6 5 VSS VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1120 $Y=790 $D=97
M2 VSS 6 7 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2670 $Y=780 $D=97
M3 Y 7 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1060 $D=97
M4 VDD A 5 VDD pfet L=1.2e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M5 6 5 VDD VDD pfet L=1.2e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1120 $Y=1910 $D=189
M6 VDD 6 7 VDD pfet L=1.2e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2670 $Y=1910 $D=189
M7 Y 7 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT CLKINVX2TR A VSS VDD Y
** N=14 EP=4 IP=0 FDC=2
M0 Y A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=630 $Y=830 $D=97
M1 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=630 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_212
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_224
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_228
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_231
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_232
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_233
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_229
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_230
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_227
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT AO22X1TR B1 B0 A0 A1 VDD VSS Y
** N=35 EP=7 IP=0 FDC=10
M0 10 B1 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=1070 $D=97
M1 9 B0 10 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=700 $Y=1070 $D=97
M2 11 A0 9 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1280 $Y=1030 $D=97
M3 VSS A1 11 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1680 $Y=1030 $D=97
M4 Y 9 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2270 $Y=810 $D=97
M5 VDD B1 8 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=1910 $D=189
M6 8 B0 VDD VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=790 $Y=1910 $D=189
M7 9 A0 8 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1280 $Y=1910 $D=189
M8 VDD 9 Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1540 $Y=3040 $D=189
M9 8 A1 9 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1760 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DLY4X1TR A VSS VDD Y
** N=37 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=790 $D=97
M1 6 5 VSS VSS nfet L=6e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=790 $D=97
M2 VSS 6 7 VSS nfet L=6e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=780 $D=97
M3 Y 7 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1060 $D=97
M4 VDD A 5 VDD pfet L=1.2e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M5 6 5 VDD VDD pfet L=6e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=1910 $D=189
M6 VDD 6 7 VDD pfet L=6e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=1910 $D=189
M7 Y 7 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3360 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT CLKAND2X2TR A B VSS VDD Y
** N=23 EP=5 IP=0 FDC=6
M0 7 A 6 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=560 $Y=990 $D=97
M1 VSS B 7 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=880 $Y=990 $D=97
M2 Y 6 VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=830 $D=97
M3 6 A VDD VDD pfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M4 VDD B 6 VDD pfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=1910 $D=189
M5 Y 6 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DFFRX1TR D CK RN QN VDD VSS Q
** N=85 EP=7 IP=0 FDC=33
M0 15 8 9 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1090 $D=97
M1 17 D 15 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=780 $Y=1090 $D=97
M2 VSS RN 17 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1100 $Y=1090 $D=97
M3 VSS CK 8 VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2080 $Y=840 $D=97
M4 11 8 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2590 $Y=940 $D=97
M5 19 11 9 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3610 $Y=1010 $D=97
M6 20 10 19 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3930 $Y=1010 $D=97
M7 VSS RN 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4250 $Y=1010 $D=97
M8 10 9 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4710 $Y=870 $D=97
M9 12 11 10 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5270 $Y=870 $D=97
M10 22 8 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5830 $Y=1110 $D=97
M11 VSS 14 22 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6150 $Y=1110 $D=97
M12 23 RN VSS VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6590 $Y=990 $D=97
M13 14 12 23 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6910 $Y=990 $D=97
M14 13 14 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7230 $Y=390 $D=97
M15 VSS 13 QN VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8190 $Y=850 $D=97
M16 Q 14 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8670 $Y=850 $D=97
M17 16 D VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=2640 $D=189
M18 9 11 16 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=780 $Y=2640 $D=189
M19 VDD RN 9 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1260 $Y=2640 $D=189
M20 VDD CK 8 VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1780 $Y=1910 $D=189
M21 11 8 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2290 $Y=1930 $D=189
M22 18 8 9 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2850 $Y=2410 $D=189
M23 VDD 10 18 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3170 $Y=2410 $D=189
M24 10 9 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3710 $Y=2410 $D=189
M25 12 8 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4540 $Y=2660 $D=189
M26 21 11 12 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5270 $Y=2660 $D=189
M27 VDD 14 21 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5600 $Y=2660 $D=189
M28 14 RN VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6060 $Y=2590 $D=189
M29 VDD 12 14 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6620 $Y=2880 $D=189
M30 13 14 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7230 $Y=2240 $D=189
M31 VDD 13 QN VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8170 $Y=1910 $D=189
M32 Q 14 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8670 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT OAI32X1TR VSS A2 A1 A0 B0 Y VDD B1
** N=35 EP=8 IP=0 FDC=10
M0 9 A2 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=390 $Y=710 $D=97
M1 VSS A1 9 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=870 $Y=710 $D=97
M2 9 A0 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1310 $Y=710 $D=97
M3 Y B0 9 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1790 $Y=710 $D=97
M4 9 B1 Y VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2270 $Y=710 $D=97
M5 10 A2 VDD VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=440 $Y=2030 $D=189
M6 11 A1 10 VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=760 $Y=2030 $D=189
M7 Y A0 11 VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1080 $Y=2030 $D=189
M8 12 B0 Y VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1630 $Y=2030 $D=189
M9 VDD B1 12 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1950 $Y=2030 $D=189
.ENDS
***************************************
.SUBCKT AOI2BB1X1TR A0N A1N B0 VDD Y VSS
** N=29 EP=6 IP=0 FDC=8
M0 7 A0N VSS VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=380 $Y=1060 $D=97
M1 VSS A1N 7 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=940 $Y=1060 $D=97
M2 Y B0 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1380 $Y=820 $D=97
M3 VSS 7 Y VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1860 $Y=820 $D=97
M4 8 A0N 7 VDD pfet L=1.2e-07 W=4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=540 $Y=2000 $D=189
M5 VDD A1N 8 VDD pfet L=1.2e-07 W=4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=2000 $D=189
M6 9 B0 VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=1910 $D=189
M7 Y 7 9 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1760 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT NAND2X1TR B VSS Y A VDD
** N=19 EP=5 IP=0 FDC=4
M0 6 B VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=710 $D=97
M1 Y A 6 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=800 $Y=710 $D=97
M2 Y B VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=1910 $D=189
M3 VDD A Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=960 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT NOR2X1TR B VDD A Y VSS
** N=20 EP=5 IP=0 FDC=4
M0 Y B VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=800 $D=97
M1 VSS A Y VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=960 $Y=800 $D=97
M2 6 B VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=560 $Y=1910 $D=189
M3 Y A 6 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=880 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT OAI21X1TR A1 VSS A0 B0 VDD Y
** N=24 EP=6 IP=0 FDC=6
M0 VSS A1 7 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=440 $Y=710 $D=97
M1 7 A0 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=920 $Y=710 $D=97
M2 Y B0 7 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1400 $Y=710 $D=97
M3 8 A1 VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=1970 $D=189
M4 Y A0 8 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=800 $Y=1970 $D=189
M5 VDD B0 Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1320 $Y=1970 $D=189
.ENDS
***************************************
.SUBCKT AOI21X1TR A1 A0 VDD B0 VSS Y
** N=24 EP=6 IP=0 FDC=6
M0 8 A1 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=490 $Y=710 $D=97
M1 Y A0 8 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=810 $Y=710 $D=97
M2 VSS B0 Y VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=850 $D=97
M3 VDD A1 7 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1920 $D=189
M4 7 A0 VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=1920 $D=189
M5 Y B0 7 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1370 $Y=1920 $D=189
.ENDS
***************************************
.SUBCKT AND2X1TR A B VSS VDD Y
** N=26 EP=5 IP=0 FDC=6
M0 7 A 6 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=950 $D=97
M1 VSS B 7 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=770 $Y=950 $D=97
M2 Y 6 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=850 $D=97
M3 6 A VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=2060 $D=189
M4 VDD B 6 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=900 $Y=2060 $D=189
M5 Y 6 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT BUFX3TR A Y VSS VDD
** N=21 EP=4 IP=0 FDC=6
M0 VSS A 5 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=750 $D=97
M1 Y 5 VSS VSS nfet L=1.2e-07 W=6.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=980 $Y=620 $D=97
M2 VSS 5 Y VSS nfet L=1.2e-07 W=6.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1460 $Y=620 $D=97
M3 VDD A 5 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M4 Y 5 VDD VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=980 $Y=1910 $D=189
M5 VDD 5 Y VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1460 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT AO22X2TR B1 B0 A0 A1 VSS Y VDD
** N=40 EP=7 IP=0 FDC=10
M0 10 B1 VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=770 $D=97
M1 8 B0 10 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=770 $Y=770 $D=97
M2 11 A0 8 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=770 $D=97
M3 VSS A1 11 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1730 $Y=770 $D=97
M4 Y 8 VSS VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2410 $Y=390 $D=97
M5 VDD B1 9 VDD pfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M6 9 B0 VDD VDD pfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=1910 $D=189
M7 8 A0 9 VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=1910 $D=189
M8 VDD 8 Y VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1520 $Y=3040 $D=189
M9 9 A1 8 VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1810 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT BUFX4TR A Y VSS VDD
** N=27 EP=4 IP=0 FDC=6
M0 VSS A 5 VSS nfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=520 $Y=630 $D=97
M1 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1080 $Y=390 $D=97
M2 VSS 5 Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1560 $Y=390 $D=97
M3 VDD A 5 VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=600 $Y=1930 $D=189
M4 Y 5 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1080 $Y=1930 $D=189
M5 VDD 5 Y VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1560 $Y=1930 $D=189
.ENDS
***************************************
.SUBCKT ICV_221
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_217
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_218
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_219
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_213
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_214
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_215
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_235 1 2 497 505 526 527 618 619 620 621 650 656 657 658 659 660 661 662 663 664
+ 709 711 714 715 719 721 722 723 724 727 728 729 731 733 734 735 736 738 742 744
+ 747 749 750 751 754 866 879 1001 1007 1061 1124 1125 1126 1127 1128 1132 1491 1493 1503 1532
+ 1535 1538 1539 1540 1541 1542 1566 1658 1659 1661 1662 1663 1664 1665 1666 1776 1973 2004 2005 2006
+ 2007 2008 2009 2010 2011 2012 2023 2038 2042 2043 2044 2049 2050 2062 2064 2067 2074 2083 2084 2088
+ 2096 2102 2103 2104 2105 2106 2107 2108 2109 2110 2111 2112 2113 2114 2115 2116 2118 2119 2218 2309
+ 2343 2387 2512 2662 2669 2724 2744 2748 2749 2784 2814 2815 3010 3011 3058
** N=256636 EP=135 IP=2815 FDC=1998
M0 229216 2218 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=265520 $Y=1000670 $D=97
M1 229238 229216 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=266950 $Y=1000820 $D=97
M2 1 229216 229238 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=267430 $Y=1000820 $D=97
M3 229303 229238 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=268860 $Y=1000930 $D=97
M4 1 229238 229303 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=269340 $Y=1000930 $D=97
M5 229303 229238 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=269900 $Y=1000930 $D=97
M6 1 229238 229303 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=270380 $Y=1000930 $D=97
M7 53417 229303 1 1 nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=271950 $Y=1000930 $D=97
M8 1 229303 53417 1 nfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=272430 $Y=1000670 $D=97
M9 53417 229303 1 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=272910 $Y=1000670 $D=97
M10 1 229303 53417 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=273390 $Y=1000670 $D=97
M11 53417 229303 1 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=273870 $Y=1000670 $D=97
M12 1 229303 53417 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=274350 $Y=1000670 $D=97
M13 53417 229303 1 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=274830 $Y=1000670 $D=97
M14 1 229303 53417 1 nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=275310 $Y=1000670 $D=97
M15 1001 101271 1 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=843110 $Y=763860 $D=97
M16 1 101271 1001 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=843590 $Y=763860 $D=97
M17 1001 101271 1 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=844070 $Y=763860 $D=97
M18 1 101271 1001 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=844550 $Y=763860 $D=97
M19 1001 101271 1 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=845110 $Y=763860 $D=97
M20 1 101271 1001 1 nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=845590 $Y=763860 $D=97
M21 1 239468 161683 1 nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1165160 $Y=720950 $D=97
M22 244639 113708 1 1 nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1165680 $Y=721110 $D=97
M23 244640 113728 244639 1 nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1166080 $Y=721110 $D=97
M24 239468 161723 244640 1 nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1166400 $Y=721110 $D=97
M25 239480 161733 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1171740 $Y=726090 $D=97
M26 1 161714 239480 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1172220 $Y=726090 $D=97
M27 239480 161723 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1172660 $Y=726090 $D=97
M28 209995 209994 239480 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1173140 $Y=726090 $D=97
M29 244643 210048 1 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185010 $Y=720890 $D=97
M30 161753 113839 244643 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185330 $Y=720890 $D=97
M31 244644 113708 161753 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185880 $Y=720890 $D=97
M32 1 113729 244644 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1186200 $Y=720890 $D=97
M33 244645 161782 1 1 nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1200750 $Y=713590 $D=97
M34 244646 113729 244645 1 nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201070 $Y=713590 $D=97
M35 161802 161786 244646 1 nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201390 $Y=713590 $D=97
M36 244647 210078 161802 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201910 $Y=713710 $D=97
M37 1 113729 244647 1 nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1202230 $Y=713710 $D=97
M38 229216 2218 2 2 pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=265520 $Y=1002270 $D=189
M39 229238 229216 2 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=266950 $Y=1002210 $D=189
M40 2 229216 229238 2 pfet L=1.2e-07 W=1.13e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=267430 $Y=1002210 $D=189
M41 229303 229238 2 2 pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=268860 $Y=1002190 $D=189
M42 2 229238 229303 2 pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=269340 $Y=1002190 $D=189
M43 229303 229238 2 2 pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=269820 $Y=1002190 $D=189
M44 2 229238 229303 2 pfet L=1.2e-07 W=1.08e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=270300 $Y=1002190 $D=189
M45 53417 229303 2 2 pfet L=1.2e-07 W=1.17e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=271950 $Y=1002190 $D=189
M46 2 229303 53417 2 pfet L=1.2e-07 W=1.17e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=272430 $Y=1002190 $D=189
M47 53417 229303 2 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=272910 $Y=1002190 $D=189
M48 2 229303 53417 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=273390 $Y=1002190 $D=189
M49 53417 229303 2 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=273870 $Y=1002190 $D=189
M50 2 229303 53417 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=274350 $Y=1002190 $D=189
M51 53417 229303 2 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=274830 $Y=1002190 $D=189
M52 2 229303 53417 2 pfet L=1.2e-07 W=1.21e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=275310 $Y=1002190 $D=189
M53 1001 101271 2 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=843190 $Y=765320 $D=189
M54 2 101271 1001 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=843670 $Y=765320 $D=189
M55 1001 101271 2 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=844150 $Y=765320 $D=189
M56 2 101271 1001 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=844630 $Y=765320 $D=189
M57 1001 101271 2 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=845110 $Y=765320 $D=189
M58 2 101271 1001 2 pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=845590 $Y=765320 $D=189
M59 2 239468 161683 2 pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1165040 $Y=722110 $D=189
M60 239468 113708 2 2 pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1165600 $Y=722110 $D=189
M61 2 113728 239468 2 pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1166080 $Y=722110 $D=189
M62 239468 161723 2 2 pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1166530 $Y=722110 $D=189
M63 244641 161733 2 2 pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1171900 $Y=724330 $D=189
M64 244642 161714 244641 2 pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1172220 $Y=724330 $D=189
M65 209995 161723 244642 2 pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1172540 $Y=724330 $D=189
M66 2 209994 209995 2 pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1173020 $Y=724710 $D=189
M67 2 210048 239505 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185010 $Y=722210 $D=189
M68 239505 113839 2 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185490 $Y=722210 $D=189
M69 161753 113708 239505 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1185970 $Y=722210 $D=189
M70 239505 113729 161753 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1186450 $Y=722210 $D=189
M71 239533 161782 2 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1200590 $Y=715050 $D=189
M72 2 113729 239533 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201070 $Y=715050 $D=189
M73 239533 161786 2 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201510 $Y=715050 $D=189
M74 161802 210078 239533 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1201990 $Y=715050 $D=189
M75 239533 113729 161802 2 pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1202470 $Y=715050 $D=189
X450 53417 1 2 58842 CLKBUFX2TR $T=493000 1001000 0 0 $X=492660 $Y=1000720
X451 2004 1 2 155638 CLKBUFX2TR $T=499000 871400 0 0 $X=498660 $Y=871120
X452 1124 1 2 193459 CLKBUFX2TR $T=647800 835400 1 0 $X=647460 $Y=831400
X453 1132 1 2 59120 CLKBUFX2TR $T=661800 965000 0 0 $X=661460 $Y=964720
X454 150107 1 2 2012 CLKBUFX2TR $T=663800 1145000 1 0 $X=663460 $Y=1141000
X455 2023 1 2 113509 CLKBUFX2TR $T=733400 957800 0 0 $X=733060 $Y=957520
X456 2038 1 2 59106 CLKBUFX2TR $T=808600 1058600 0 0 $X=808260 $Y=1058320
X457 155638 1 2 111502 CLKBUFX2TR $T=821800 749000 0 0 $X=821460 $Y=748720
X458 505 1 2 113398 CLKBUFX2TR $T=883000 1159400 1 0 $X=882660 $Y=1155400
X459 107645 1 2 59515 CLKBUFX2TR $T=939400 770600 1 0 $X=939060 $Y=766600
X460 57764 1 2 1658 CLKBUFX2TR $T=957400 1159400 1 0 $X=957060 $Y=1155400
X461 208907 1 2 161051 CLKBUFX2TR $T=988200 741800 0 0 $X=987860 $Y=741520
X462 2062 1 2 113735 CLKBUFX2TR $T=988200 1065800 1 0 $X=987860 $Y=1061800
X463 2064 1 2 113578 CLKBUFX2TR $T=988200 1173800 0 0 $X=987860 $Y=1173520
X464 58842 1 2 113808 CLKBUFX2TR $T=1009400 734600 0 0 $X=1009060 $Y=734320
X465 111502 1 2 113713 CLKBUFX2TR $T=1129400 734600 0 0 $X=1129060 $Y=734320
X466 115271 1 2 161655 CLKBUFX2TR $T=1186200 734600 0 180 $X=1184260 $Y=730600
X467 161765 1 2 161733 CLKBUFX2TR $T=1193000 720200 1 180 $X=1191060 $Y=719920
X468 161791 1 2 115271 CLKBUFX2TR $T=1203000 734600 0 0 $X=1202660 $Y=734320
X469 113713 1 2 115256 CLKBUFX2TR $T=1219800 734600 0 0 $X=1219460 $Y=734320
X470 2118 1 2 113966 CLKBUFX2TR $T=1475800 1159400 1 180 $X=1473860 $Y=1159120
X471 1776 1 2 111657 CLKBUFX2TR $T=1542200 698600 1 0 $X=1541860 $Y=694600
X472 866 1 2 58776 CLKBUFX2TR $T=1598600 749000 0 0 $X=1598260 $Y=748720
X562 879 61957 2 1 CLKINVX8TR $T=263000 878600 0 0 $X=262660 $Y=878320
X563 61957 137750 2 1 CLKINVX8TR $T=269800 921800 0 180 $X=266660 $Y=917800
X564 101271 113461 2 1 CLKINVX8TR $T=1135000 734600 0 0 $X=1134660 $Y=734320
X602 137750 63522 1 2 CLKINVX20TR $T=288600 921800 0 180 $X=282660 $Y=917800
X603 63522 100051 1 2 CLKINVX20TR $T=683800 835400 0 180 $X=677860 $Y=831400
X604 100051 101271 1 2 CLKINVX20TR $T=825400 763400 0 0 $X=825060 $Y=763120
X605 101271 527 1 2 CLKINVX20TR $T=1183800 734600 0 0 $X=1183460 $Y=734320
X745 1 2 53417 2005 INVX1TR $T=493400 1008200 0 0 $X=493060 $Y=1007920
X746 1 2 113713 161759 INVX1TR $T=1188200 734600 1 0 $X=1187860 $Y=730600
X747 1 2 161760 161758 INVX1TR $T=1192200 713000 1 180 $X=1190660 $Y=712720
X748 1 2 161808 161765 INVX1TR $T=1209800 720200 1 0 $X=1209460 $Y=716200
X769 1007 155638 2 1 2309 AND2X2TR $T=516600 756200 1 180 $X=514260 $Y=755920
X770 1061 155638 2 1 2343 AND2X2TR $T=564600 756200 1 180 $X=562260 $Y=755920
X771 650 155638 2 1 2387 AND2X2TR $T=641800 756200 1 180 $X=639460 $Y=755920
X772 709 111502 2 1 2512 AND2X2TR $T=825400 756200 1 180 $X=823060 $Y=755920
X773 661 111502 2 1 2043 AND2X2TR $T=840200 749000 0 180 $X=837860 $Y=745000
X774 714 111502 2 1 2044 AND2X2TR $T=846200 749000 1 180 $X=843860 $Y=748720
X775 722 111502 2 1 2662 AND2X2TR $T=1100600 734600 1 180 $X=1098260 $Y=734320
X776 2088 111502 2 1 2084 AND2X2TR $T=1124600 734600 1 180 $X=1122260 $Y=734320
X777 2102 115256 2 1 2724 AND2X2TR $T=1254600 734600 1 180 $X=1252260 $Y=734320
X778 2749 115256 2 1 2748 AND2X2TR $T=1298600 734600 1 180 $X=1296260 $Y=734320
X779 2104 115256 2 1 2784 AND2X2TR $T=1345800 734600 0 0 $X=1345460 $Y=734320
X780 2105 115256 2 1 2106 AND2X2TR $T=1397400 734600 0 0 $X=1397060 $Y=734320
X781 2110 115256 2 1 2115 AND2X2TR $T=1412200 749000 1 0 $X=1411860 $Y=745000
X782 751 115256 2 1 2814 AND2X2TR $T=1412200 756200 1 0 $X=1411860 $Y=752200
X816 193459 1 2 112307 DLY3X1TR $T=649400 835400 1 0 $X=649060 $Y=831400
X817 2042 1 2 155527 DLY3X1TR $T=822200 986600 1 0 $X=821860 $Y=982600
X818 161659 1 2 161674 DLY3X1TR $T=1145800 713000 0 0 $X=1145460 $Y=712720
X819 161692 1 2 161685 DLY3X1TR $T=1156600 713000 1 0 $X=1156260 $Y=709000
X820 161706 1 2 161699 DLY3X1TR $T=1161800 713000 0 0 $X=1161460 $Y=712720
X821 210033 1 2 161744 DLY3X1TR $T=1180200 713000 1 0 $X=1179860 $Y=709000
X822 161740 1 2 161734 DLY3X1TR $T=1181000 727400 0 0 $X=1180660 $Y=727120
X823 210047 1 2 161748 DLY3X1TR $T=1183800 741800 1 0 $X=1183460 $Y=737800
X824 210068 1 2 161789 DLY3X1TR $T=1199000 734600 1 0 $X=1198660 $Y=730600
X825 113917 1 2 161828 DLY3X1TR $T=1215800 741800 1 0 $X=1215460 $Y=737800
X826 161817 1 2 161827 DLY3X1TR $T=1216200 734600 1 0 $X=1215860 $Y=730600
X827 149685 1 2 58898 DLY2X1TR $T=650200 849800 0 0 $X=649860 $Y=849520
X828 149788 1 2 112800 DLY2X1TR $T=650200 857000 0 0 $X=649860 $Y=856720
X829 149916 1 2 58934 DLY2X1TR $T=650600 842600 0 0 $X=650260 $Y=842320
X830 149686 1 2 112417 DLY2X1TR $T=650600 849800 1 0 $X=650260 $Y=845800
X831 2009 1 2 149788 DLY2X1TR $T=650600 857000 1 0 $X=650260 $Y=853000
X832 1125 1 2 656 DLY2X1TR $T=651400 1145000 0 0 $X=651060 $Y=1144720
X833 1127 1 2 149685 DLY2X1TR $T=654200 849800 0 0 $X=653860 $Y=849520
X834 2011 1 2 149916 DLY2X1TR $T=654200 857000 0 0 $X=653860 $Y=856720
X835 1126 1 2 149686 DLY2X1TR $T=654600 849800 1 0 $X=654260 $Y=845800
X836 152692 1 2 152691 DLY2X1TR $T=738200 1029800 1 0 $X=737860 $Y=1025800
X837 660 1 2 155706 DLY2X1TR $T=821000 993800 0 0 $X=820660 $Y=993520
X838 662 1 2 2050 DLY2X1TR $T=929000 1130600 1 0 $X=928660 $Y=1126600
X839 113839 1 2 161775 DLY2X1TR $T=1193000 734600 1 0 $X=1192660 $Y=730600
X840 161826 1 2 161852 DLY2X1TR $T=1234200 734600 0 0 $X=1233860 $Y=734320
X841 657 1 2 1128 DLY1X1TR $T=653000 1130600 1 0 $X=652660 $Y=1126600
X842 497 1 2 107645 DLY1X1TR $T=724200 770600 1 0 $X=723860 $Y=766600
X843 155706 1 2 58355 DLY1X1TR $T=817000 993800 0 0 $X=816660 $Y=993520
X844 155527 1 2 58354 DLY1X1TR $T=818200 986600 1 0 $X=817860 $Y=982600
X845 659 1 2 57764 DLY1X1TR $T=822200 1065800 1 0 $X=821860 $Y=1061800
X846 663 1 2 2049 DLY1X1TR $T=925000 1130600 1 0 $X=924660 $Y=1126600
X847 2010 1 2 152692 CLKINVX2TR $T=655800 1022600 0 0 $X=655460 $Y=1022320
X848 2008 1 2 150083 CLKINVX2TR $T=655800 1044200 1 0 $X=655460 $Y=1040200
X849 150083 1 2 150107 CLKINVX2TR $T=663000 1044200 0 0 $X=662660 $Y=1043920
X850 152691 1 2 664 CLKINVX2TR $T=737000 1029800 1 0 $X=736660 $Y=1025800
X851 2007 1 2 113812 CLKINVX2TR $T=783800 1094600 1 0 $X=783460 $Y=1090600
X852 2006 1 2 113832 CLKINVX2TR $T=786600 1094600 0 0 $X=786260 $Y=1094320
X967 58355 161655 111502 58776 2 1 723 AO22X1TR $T=984600 849800 1 0 $X=984260 $Y=845800
X968 161051 161655 111502 2067 2 1 1491 AO22X1TR $T=985800 749000 0 0 $X=985460 $Y=748720
X969 58354 161655 111502 111657 2 1 721 AO22X1TR $T=986600 842600 1 0 $X=986260 $Y=838600
X970 112307 161655 111502 1493 2 1 2074 AO22X1TR $T=1021000 741800 1 0 $X=1020660 $Y=737800
X971 112417 161655 111502 58935 2 1 1503 AO22X1TR $T=1036600 741800 1 0 $X=1036260 $Y=737800
X972 58898 161655 111502 112801 2 1 711 AO22X1TR $T=1049800 741800 1 0 $X=1049460 $Y=737800
X973 58934 161655 111502 526 2 1 2083 AO22X1TR $T=1059800 741800 1 0 $X=1059460 $Y=737800
X974 112800 161655 111502 719 2 1 715 AO22X1TR $T=1078600 741800 1 0 $X=1078260 $Y=737800
X975 1532 113713 113510 161655 2 1 728 AO22X1TR $T=1139400 734600 0 0 $X=1139060 $Y=734320
X976 161686 161673 161683 161669 2 1 161645 AO22X1TR $T=1145000 720200 0 0 $X=1144660 $Y=719920
X977 113398 113713 161673 161655 2 1 733 AO22X1TR $T=1145400 734600 0 0 $X=1145060 $Y=734320
X978 161698 113597 113630 161689 2 1 161706 AO22X1TR $T=1157800 720200 1 180 $X=1154660 $Y=719920
X979 113578 113713 113597 161655 2 1 731 AO22X1TR $T=1155400 734600 0 0 $X=1155060 $Y=734320
X980 724 113713 161703 161655 2 1 1538 AO22X1TR $T=1159800 734600 0 0 $X=1159460 $Y=734320
X981 59106 113713 161723 161655 2 1 735 AO22X1TR $T=1164600 734600 0 0 $X=1164260 $Y=734320
X982 113509 113713 113728 161655 2 1 736 AO22X1TR $T=1170200 734600 0 0 $X=1169860 $Y=734320
X983 161724 113708 113728 161735 2 1 161727 AO22X1TR $T=1172200 713000 0 0 $X=1171860 $Y=712720
X984 59120 113713 113708 161655 2 1 738 AO22X1TR $T=1176200 734600 0 0 $X=1175860 $Y=734320
X985 113735 113713 161752 161655 2 1 2096 AO22X1TR $T=1183800 734600 1 180 $X=1180660 $Y=734320
X986 161754 161752 113818 161745 2 1 210047 AO22X1TR $T=1185800 727400 0 180 $X=1182660 $Y=723400
X987 161775 161759 113713 113812 2 1 1540 AO22X1TR $T=1192200 734600 1 180 $X=1189060 $Y=734320
X988 161775 161759 113713 113832 2 1 1542 AO22X1TR $T=1190200 734600 1 0 $X=1189860 $Y=730600
X989 734 113713 161792 115271 2 1 1539 AO22X1TR $T=1199000 734600 1 180 $X=1195860 $Y=734320
X990 161808 210107 113917 161760 2 1 161835 AO22X1TR $T=1210200 713000 1 180 $X=1207060 $Y=712720
X991 1541 113713 161815 115271 2 1 727 AO22X1TR $T=1210200 734600 1 180 $X=1207060 $Y=734320
X992 113966 113713 161828 115271 2 1 1535 AO22X1TR $T=1217000 734600 1 180 $X=1213860 $Y=734320
X993 161824 161826 161779 210134 2 1 161848 AO22X1TR $T=1217800 727400 0 0 $X=1217460 $Y=727120
X994 742 115256 161852 115271 2 1 729 AO22X1TR $T=1234200 734600 1 180 $X=1231060 $Y=734320
X995 1661 115271 115256 1659 2 1 754 AO22X1TR $T=1415000 1058600 1 180 $X=1411860 $Y=1058320
X996 658 1 2 208907 DLY4X1TR $T=985800 749000 1 0 $X=985460 $Y=745000
X997 161656 1 2 161646 DLY4X1TR $T=1133400 727400 0 0 $X=1133060 $Y=727120
X998 161654 1 2 161677 DLY4X1TR $T=1142200 734600 1 0 $X=1141860 $Y=730600
X999 161664 1 2 161670 DLY4X1TR $T=1144200 741800 1 0 $X=1143860 $Y=737800
X1000 161674 1 2 161673 DLY4X1TR $T=1145400 720200 1 0 $X=1145060 $Y=716200
X1001 161670 1 2 113510 DLY4X1TR $T=1146200 734600 1 0 $X=1145860 $Y=730600
X1002 161700 1 2 161682 DLY4X1TR $T=1151400 727400 0 0 $X=1151060 $Y=727120
X1003 161685 1 2 113597 DLY4X1TR $T=1152600 713000 1 0 $X=1152260 $Y=709000
X1004 209974 1 2 209975 DLY4X1TR $T=1159800 727400 0 0 $X=1159460 $Y=727120
X1005 161715 1 2 161703 DLY4X1TR $T=1160600 741800 1 0 $X=1160260 $Y=737800
X1006 161710 1 2 161723 DLY4X1TR $T=1164600 727400 0 0 $X=1164260 $Y=727120
X1007 161709 1 2 161715 DLY4X1TR $T=1164600 741800 1 0 $X=1164260 $Y=737800
X1008 161722 1 2 113728 DLY4X1TR $T=1165800 705800 0 0 $X=1165460 $Y=705520
X1009 161716 1 2 161722 DLY4X1TR $T=1166200 713000 0 0 $X=1165860 $Y=712720
X1010 161719 1 2 161710 DLY4X1TR $T=1168600 727400 0 0 $X=1168260 $Y=727120
X1011 209995 1 2 161732 DLY4X1TR $T=1172600 727400 0 0 $X=1172260 $Y=727120
X1012 161734 1 2 161752 DLY4X1TR $T=1177000 727400 0 0 $X=1176660 $Y=727120
X1013 161744 1 2 113708 DLY4X1TR $T=1179800 720200 1 0 $X=1179460 $Y=716200
X1014 210034 1 2 210048 DLY4X1TR $T=1180600 720200 0 0 $X=1180260 $Y=719920
X1015 161770 1 2 210060 DLY4X1TR $T=1187000 727400 0 0 $X=1186660 $Y=727120
X1016 210059 1 2 161782 DLY4X1TR $T=1188200 713000 1 0 $X=1187860 $Y=709000
X1017 161753 1 2 161761 DLY4X1TR $T=1188200 720200 1 0 $X=1187860 $Y=716200
X1018 161766 1 2 210062 DLY4X1TR $T=1193000 713000 0 0 $X=1192660 $Y=712720
X1019 161767 1 2 161774 DLY4X1TR $T=1193000 720200 0 0 $X=1192660 $Y=719920
X1020 161776 1 2 161780 DLY4X1TR $T=1194600 713000 1 0 $X=1194260 $Y=709000
X1021 113856 1 2 161760 DLY4X1TR $T=1196600 720200 1 0 $X=1196260 $Y=716200
X1022 161781 1 2 210078 DLY4X1TR $T=1198600 713000 1 0 $X=1198260 $Y=709000
X1023 161789 1 2 161792 DLY4X1TR $T=1200200 727400 0 0 $X=1199860 $Y=727120
X1024 161790 1 2 161781 DLY4X1TR $T=1202600 713000 1 0 $X=1202260 $Y=709000
X1025 161793 1 2 161786 DLY4X1TR $T=1203800 720200 1 0 $X=1203460 $Y=716200
X1026 161799 1 2 161803 DLY4X1TR $T=1204200 727400 0 0 $X=1203860 $Y=727120
X1027 161802 1 2 161798 DLY4X1TR $T=1207000 705800 0 0 $X=1206660 $Y=705520
X1028 161811 1 2 161818 DLY4X1TR $T=1208600 727400 0 0 $X=1208260 $Y=727120
X1029 161809 1 2 161807 DLY4X1TR $T=1210200 727400 1 0 $X=1209860 $Y=723400
X1030 161827 1 2 161815 DLY4X1TR $T=1212200 734600 1 0 $X=1211860 $Y=730600
X1031 210113 1 2 113917 DLY4X1TR $T=1213000 713000 1 0 $X=1212660 $Y=709000
X1032 161835 1 2 161833 DLY4X1TR $T=1222200 713000 0 0 $X=1221860 $Y=712720
X1033 161848 1 2 161838 DLY4X1TR $T=1225000 720200 1 0 $X=1224660 $Y=716200
X1034 210188 1 2 161826 DLY4X1TR $T=1233800 720200 0 0 $X=1233460 $Y=719920
X1035 744 111502 1 2 2669 CLKAND2X2TR $T=1115800 734600 1 180 $X=1113460 $Y=734320
X1036 2103 115256 1 2 2744 CLKAND2X2TR $T=1289800 734600 1 180 $X=1287460 $Y=734320
X1037 161646 113461 113808 161654 2 1 161664 DFFRX1TR $T=1133000 734600 1 0 $X=1132660 $Y=730600
X1038 161645 113461 113808 244632 2 1 161659 DFFRX1TR $T=1134200 720200 0 0 $X=1133860 $Y=719920
X1039 161682 113461 113808 209974 2 1 161709 DFFRX1TR $T=1151800 734600 1 0 $X=1151460 $Y=730600
X1040 161699 113461 113808 244633 2 1 161692 DFFRX1TR $T=1161800 713000 1 180 $X=1152260 $Y=712720
X1041 161732 113461 113808 244634 2 1 161719 DFFRX1TR $T=1172600 734600 0 180 $X=1163060 $Y=730600
X1042 161727 113461 113808 244635 2 1 161716 DFFRX1TR $T=1173800 713000 0 180 $X=1164260 $Y=709000
X1043 161748 113461 113808 244636 2 1 161740 DFFRX1TR $T=1184600 734600 0 180 $X=1175060 $Y=730600
X1044 161761 113461 113808 210034 2 1 210033 DFFRX1TR $T=1189000 713000 1 180 $X=1179460 $Y=712720
X1045 161758 113461 113808 210059 2 1 161766 DFFRX1TR $T=1180200 705800 0 0 $X=1179860 $Y=705520
X1046 210060 113461 113808 161809 2 1 210068 DFFRX1TR $T=1191000 727400 0 0 $X=1190660 $Y=727120
X1047 161798 113461 113808 161790 2 1 161776 DFFRX1TR $T=1207000 705800 1 180 $X=1197460 $Y=705520
X1048 161803 113461 113808 161811 2 1 161817 DFFRX1TR $T=1203000 734600 1 0 $X=1202660 $Y=730600
X1049 161833 113461 113808 244637 2 1 210113 DFFRX1TR $T=1222200 713000 1 180 $X=1212660 $Y=712720
X1050 161838 113461 113808 244638 2 1 210188 DFFRX1TR $T=1224600 720200 0 0 $X=1224260 $Y=719920
X1051 1 161733 161678 113510 161663 161656 2 161677 OAI32X1TR $T=1143800 727400 1 180 $X=1140660 $Y=727120
X1052 1 161733 161697 161703 161694 161700 2 209975 OAI32X1TR $T=1159000 727400 1 0 $X=1158660 $Y=723400
X1053 1 161765 161774 161792 161757 161770 2 161807 OAI32X1TR $T=1193400 727400 1 0 $X=1193060 $Y=723400
X1054 1 113839 161797 161815 161819 161799 2 161818 OAI32X1TR $T=1204600 727400 1 0 $X=1204260 $Y=723400
X1055 161733 161673 161686 2 161663 1 AOI2BB1X1TR $T=1146600 727400 0 180 $X=1143860 $Y=723400
X1056 161733 113597 161698 2 161694 1 AOI2BB1X1TR $T=1155400 727400 1 0 $X=1155060 $Y=723400
X1057 161733 161752 161754 2 161757 1 AOI2BB1X1TR $T=1187400 727400 1 0 $X=1187060 $Y=723400
X1058 161765 161826 161824 2 161819 1 AOI2BB1X1TR $T=1215000 720200 1 180 $X=1212260 $Y=719920
X1059 161673 1 161678 161683 2 NAND2X1TR $T=1145800 727400 0 0 $X=1145460 $Y=727120
X1060 113597 1 161697 113630 2 NAND2X1TR $T=1157000 727400 1 180 $X=1155060 $Y=727120
X1061 113708 1 161714 113728 2 NAND2X1TR $T=1165800 727400 1 0 $X=1165460 $Y=723400
X1062 161752 1 161767 113818 2 NAND2X1TR $T=1190600 727400 1 0 $X=1190260 $Y=723400
X1063 161780 1 113839 161782 2 NAND2X1TR $T=1200200 720200 0 0 $X=1199860 $Y=719920
X1064 210078 1 113729 161782 2 NAND2X1TR $T=1202200 720200 0 180 $X=1200260 $Y=716200
X1065 161826 1 161797 161779 2 NAND2X1TR $T=1214200 727400 1 180 $X=1212260 $Y=727120
X1066 161733 2 161673 161669 1 NOR2X1TR $T=1147800 720200 0 0 $X=1147460 $Y=719920
X1067 161677 2 161678 113630 1 NOR2X1TR $T=1149800 727400 0 0 $X=1149460 $Y=727120
X1068 161733 2 113597 161689 1 NOR2X1TR $T=1151800 720200 1 0 $X=1151460 $Y=716200
X1069 209975 2 161697 113818 1 NOR2X1TR $T=1162600 727400 1 0 $X=1162260 $Y=723400
X1070 161733 2 113728 161724 1 NOR2X1TR $T=1168200 720200 0 0 $X=1167860 $Y=719920
X1071 161733 2 161752 161745 1 NOR2X1TR $T=1177400 727400 1 0 $X=1177060 $Y=723400
X1072 161807 2 161774 161779 1 NOR2X1TR $T=1197400 727400 1 0 $X=1197060 $Y=723400
X1073 113839 2 113713 161791 1 NOR2X1TR $T=1200600 734600 0 0 $X=1200260 $Y=734320
X1074 161786 2 113839 161808 1 NOR2X1TR $T=1205000 720200 0 0 $X=1204660 $Y=719920
X1075 161818 2 161797 210107 1 NOR2X1TR $T=1208600 727400 1 0 $X=1208260 $Y=723400
X1076 161765 2 161826 210134 1 NOR2X1TR $T=1219000 720200 1 0 $X=1218660 $Y=716200
X1077 161733 1 161683 113729 2 161686 OAI21X1TR $T=1151800 720200 0 0 $X=1151460 $Y=719920
X1078 161733 1 113630 113729 2 161698 OAI21X1TR $T=1158600 720200 0 0 $X=1158260 $Y=719920
X1079 161735 1 161724 161723 2 209994 OAI21X1TR $T=1174200 720200 1 180 $X=1171860 $Y=719920
X1080 161733 1 113708 113729 2 161735 OAI21X1TR $T=1177000 720200 0 0 $X=1176660 $Y=719920
X1081 161733 1 113818 113729 2 161754 OAI21X1TR $T=1187800 720200 0 0 $X=1187460 $Y=719920
X1082 161765 1 161779 113729 2 161824 OAI21X1TR $T=1203000 727400 0 180 $X=1200660 $Y=723400
X1083 161780 161786 2 210062 1 113856 AOI21X1TR $T=1199000 713000 1 180 $X=1196660 $Y=712720
X1084 113917 210107 1 2 161793 AND2X1TR $T=1209800 720200 0 180 $X=1207460 $Y=716200
X1085 2108 58935 1 2 BUFX3TR $T=1412200 943400 0 0 $X=1411860 $Y=943120
X1086 2109 115271 115256 2114 1 620 2 AO22X2TR $T=1412200 1065800 1 0 $X=1411860 $Y=1061800
X1087 59515 115271 115256 1662 1 747 2 AO22X2TR $T=1412600 993800 0 0 $X=1412260 $Y=993520
X1088 2112 115271 115256 1665 1 1566 2 AO22X2TR $T=1413000 1044200 1 0 $X=1412660 $Y=1040200
X1089 1658 115271 115256 1666 1 619 2 AO22X2TR $T=1413000 1051400 0 0 $X=1412660 $Y=1051120
X1090 2113 115271 115256 1663 1 749 2 AO22X2TR $T=1413800 1022600 0 0 $X=1413460 $Y=1022320
X1091 2111 115271 115256 2116 1 750 2 AO22X2TR $T=1413800 1029800 1 0 $X=1413460 $Y=1025800
X1092 618 115271 115256 1664 1 621 2 AO22X2TR $T=1413800 1029800 0 0 $X=1413460 $Y=1029520
X1093 2107 526 1 2 BUFX4TR $T=1412200 1188200 0 0 $X=1411860 $Y=1187920
X1094 2815 719 1 2 BUFX4TR $T=1414600 1188200 0 0 $X=1414260 $Y=1187920
X1095 2119 112801 1 2 BUFX4TR $T=1708600 749000 0 0 $X=1708260 $Y=748720
X1096 1973 3058 1 2 BUFX4TR $T=1734600 1188200 1 0 $X=1734260 $Y=1184200
X1097 3010 3011 1 2 BUFX4TR $T=1734600 1217000 0 0 $X=1734260 $Y=1216720
.ENDS
***************************************
.SUBCKT ICV_207
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_208
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_209
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_184
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_204
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_205
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_186
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_187
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT BUFX20TR A Y VDD VSS
** N=73 EP=4 IP=0 FDC=28
M0 5 A VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=390 $D=97
M1 VSS A 5 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=390 $D=97
M2 5 A VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1370 $Y=390 $D=97
M3 VSS A 5 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1850 $Y=390 $D=97
M4 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2330 $Y=390 $D=97
M5 VSS 5 Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2810 $Y=390 $D=97
M6 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3290 $Y=390 $D=97
M7 VSS 5 Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3770 $Y=390 $D=97
M8 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4250 $Y=390 $D=97
M9 VSS 5 Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4730 $Y=390 $D=97
M10 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5210 $Y=390 $D=97
M11 VSS 5 Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5690 $Y=390 $D=97
M12 Y 5 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6170 $Y=390 $D=97
M13 VSS 5 Y VSS nfet L=1.2e-07 W=6.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6690 $Y=650 $D=97
M14 5 A VDD VDD pfet L=1.2e-07 W=1.22e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M15 VDD A 5 VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=1910 $D=189
M16 5 A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1370 $Y=1910 $D=189
M17 VDD A 5 VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1850 $Y=1910 $D=189
M18 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2330 $Y=1910 $D=189
M19 VDD 5 Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2810 $Y=1910 $D=189
M20 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3290 $Y=1910 $D=189
M21 VDD 5 Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3770 $Y=1910 $D=189
M22 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4250 $Y=1910 $D=189
M23 VDD 5 Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4730 $Y=1910 $D=189
M24 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5210 $Y=1910 $D=189
M25 VDD 5 Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5690 $Y=1910 $D=189
M26 Y 5 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6170 $Y=1910 $D=189
M27 VDD 5 Y VDD pfet L=1.2e-07 W=1.04e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6650 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_210 1 2 347 424 426 434 435 476 477 478 834 847 850 919 980 983 1025 1026 1027 1028
+ 1030 1143 1353 1356 1357 1359 1361 1362 1368 1369 1370 1371 1372 1378 1395 1403 1858
** N=131371 EP=37 IP=596 FDC=109
M0 1 1378 125073 1 nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1734880 $Y=1309370 $D=97
M1 1371 125073 1 1 nfet L=1.2e-07 W=7.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1735440 $Y=1309290 $D=97
M2 1 125073 1371 1 nfet L=1.2e-07 W=7.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1735920 $Y=1309290 $D=97
M3 2 1378 125073 2 pfet L=1.2e-07 W=1.16e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1734960 $Y=1307530 $D=189
M4 1371 125073 2 2 pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1735440 $Y=1307410 $D=189
M5 2 125073 1371 2 pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1735920 $Y=1307410 $D=189
M6 1371 125073 2 2 pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1736400 $Y=1307410 $D=189
X171 426 1 2 834 CLKBUFX2TR $T=879000 1260200 0 0 $X=878660 $Y=1259920
X172 424 1 2 477 CLKBUFX2TR $T=883800 1267400 1 0 $X=883460 $Y=1263400
X173 847 1 2 478 CLKBUFX2TR $T=925000 1260200 0 0 $X=924660 $Y=1259920
X174 850 1 2 476 CLKBUFX2TR $T=928600 1260200 0 0 $X=928260 $Y=1259920
X175 347 1 2 1028 CLKBUFX2TR $T=939400 1260200 0 0 $X=939060 $Y=1259920
X176 1353 1 2 1858 CLKBUFX2TR $T=958600 1317800 0 0 $X=958260 $Y=1317520
X177 919 1 2 1027 CLKBUFX2TR $T=988200 1281800 1 0 $X=987860 $Y=1277800
X178 1357 1 2 435 CLKBUFX2TR $T=1076600 1346600 1 0 $X=1076260 $Y=1342600
X179 1025 1 2 1359 CLKBUFX2TR $T=1386200 1281800 0 0 $X=1385860 $Y=1281520
X180 1026 1 2 1362 CLKBUFX2TR $T=1387800 1281800 0 0 $X=1387460 $Y=1281520
X181 1030 1 2 1361 CLKBUFX2TR $T=1397400 1346600 0 0 $X=1397060 $Y=1346320
X231 980 1356 1 2 BUFX3TR $T=1131400 1325000 0 0 $X=1131060 $Y=1324720
X232 983 434 1 2 BUFX3TR $T=1207800 1289000 1 0 $X=1207460 $Y=1285000
X233 1143 1370 1 2 BUFX3TR $T=1542600 1397000 1 0 $X=1542260 $Y=1393000
X234 1368 1369 1 2 BUFX4TR $T=1530200 1325000 1 0 $X=1529860 $Y=1321000
X235 1395 1372 1 2 BUFX4TR $T=1734600 1281800 1 0 $X=1734260 $Y=1277800
X287 1372 1403 2 1 BUFX20TR $T=1729400 1346600 0 0 $X=1729060 $Y=1346320
.ENDS
***************************************
.SUBCKT ICV_197
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_192
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_202 1 2 221 1495 1838 1841 1858 1862 1895 1948 1949 1950 1951 1967 1968 1969 1975 1976 1977 1978
+ 1984 1987 1988 1995 1998 2007 2014 2027 2045 2224 2225 2226 2505 2663 2664 2665 2671 2713 2714 2788
+ 2790 2822 2823
** N=210263 EP=43 IP=550 FDC=274
X149 221 1 2 2045 CLKBUFX2TR $T=263000 1735400 1 0 $X=262660 $Y=1731400
X150 1495 1 2 2505 CLKBUFX2TR $T=1181800 1454600 0 0 $X=1181460 $Y=1454320
X182 1895 1 2 2224 CLKINVX2TR $T=634200 1706600 1 0 $X=633860 $Y=1702600
X183 2225 1 2 2226 CLKINVX2TR $T=636600 1692200 0 0 $X=636260 $Y=1691920
X184 2663 2664 1 2 BUFX3TR $T=1413400 1663400 0 0 $X=1413060 $Y=1663120
X185 1858 1984 1 2 BUFX3TR $T=1716200 1490600 0 0 $X=1715860 $Y=1490320
X186 2007 2027 1 2 BUFX3TR $T=1735000 1620200 1 0 $X=1734660 $Y=1616200
X187 2665 1950 1 2 BUFX4TR $T=1415800 1699400 1 0 $X=1415460 $Y=1695400
X188 2713 1949 1 2 BUFX4TR $T=1467800 1735400 1 0 $X=1467460 $Y=1731400
X189 2788 1968 1 2 BUFX4TR $T=1614200 1670600 0 0 $X=1613860 $Y=1670320
X190 1838 1975 1 2 BUFX4TR $T=1692200 1548200 0 0 $X=1691860 $Y=1547920
X191 1841 1976 1 2 BUFX4TR $T=1693800 1562600 0 0 $X=1693460 $Y=1562320
X192 2823 1978 1 2 BUFX4TR $T=1698200 1613000 0 0 $X=1697860 $Y=1612720
X193 1998 2014 1 2 BUFX4TR $T=1734600 1447400 0 0 $X=1734260 $Y=1447120
X194 1862 1995 1 2 BUFX4TR $T=1734600 1505000 0 0 $X=1734260 $Y=1504720
X217 2014 1948 2 1 BUFX20TR $T=1401000 1663400 0 0 $X=1400660 $Y=1663120
X218 1995 1951 2 1 BUFX20TR $T=1446200 1735400 1 0 $X=1445860 $Y=1731400
X219 2714 2671 2 1 BUFX20TR $T=1470200 1735400 1 0 $X=1469860 $Y=1731400
X220 2027 1967 2 1 BUFX20TR $T=1605800 1735400 1 0 $X=1605460 $Y=1731400
X221 2790 1969 2 1 BUFX20TR $T=1624200 1735400 1 0 $X=1623860 $Y=1731400
X222 2822 1977 2 1 BUFX20TR $T=1695400 1483400 0 0 $X=1695060 $Y=1483120
X223 1988 1987 2 1 BUFX20TR $T=1729400 1706600 1 0 $X=1729060 $Y=1702600
.ENDS
***************************************
.SUBCKT CLKINVX16TR A VSS Y VDD
** N=34 EP=4 IP=0 FDC=14
M0 Y A VSS VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=680 $D=97
M1 VSS A Y VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1340 $Y=680 $D=97
M2 Y A VSS VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1900 $Y=680 $D=97
M3 VSS A Y VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2380 $Y=680 $D=97
M4 Y A VSS VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2940 $Y=680 $D=97
M5 VSS A Y VSS nfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3420 $Y=680 $D=97
M6 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=900 $Y=1910 $D=189
M7 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1380 $Y=1910 $D=189
M8 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1860 $Y=1910 $D=189
M9 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2340 $Y=1910 $D=189
M10 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2820 $Y=1910 $D=189
M11 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3300 $Y=1910 $D=189
M12 Y A VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3780 $Y=1910 $D=189
M13 VDD A Y VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4260 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_267
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_266
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT DFFHQX8TR CK D VDD VSS Q
** N=118 EP=5 IP=0 FDC=47
M0 VSS CK 6 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=770 $D=97
M1 9 CK VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=830 $D=97
M2 VSS D 7 VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1920 $Y=870 $D=97
M3 11 6 VSS VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=590 $D=97
M4 15 9 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3540 $Y=710 $D=97
M5 8 7 15 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3860 $Y=710 $D=97
M6 17 7 8 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4500 $Y=500 $D=97
M7 VSS 9 17 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4820 $Y=500 $D=97
M8 20 11 8 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5700 $Y=900 $D=97
M9 VSS 10 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6020 $Y=900 $D=97
M10 10 8 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6420 $Y=390 $D=97
M11 VSS 8 10 VSS nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6900 $Y=670 $D=97
M12 13 11 10 VSS nfet L=1.2e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7910 $Y=600 $D=97
M13 10 11 13 VSS nfet L=1.2e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8390 $Y=600 $D=97
M14 21 9 13 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9370 $Y=600 $D=97
M15 VSS 12 21 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9710 $Y=600 $D=97
M16 VSS 13 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10270 $Y=1110 $D=97
M17 Q 13 VSS VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10670 $Y=570 $D=97
M18 VSS 13 Q VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11150 $Y=570 $D=97
M19 Q 13 VSS VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11630 $Y=570 $D=97
M20 VSS 13 Q VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12110 $Y=570 $D=97
M21 Q 13 VSS VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12590 $Y=570 $D=97
M22 VDD CK 6 VDD pfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1910 $D=189
M23 14 CK VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=1910 $D=189
M24 9 11 14 VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1180 $Y=1910 $D=189
M25 VDD D 7 VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2000 $Y=1910 $D=189
M26 11 6 VDD VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=1910 $D=189
M27 VDD 6 11 VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2920 $Y=1910 $D=189
M28 16 7 8 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3860 $Y=2140 $D=189
M29 VDD 11 16 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4180 $Y=2140 $D=189
M30 18 11 VDD VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4740 $Y=2140 $D=189
M31 8 7 18 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5060 $Y=2140 $D=189
M32 19 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5590 $Y=1930 $D=189
M33 VDD 10 19 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5940 $Y=1930 $D=189
M34 10 8 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6420 $Y=1930 $D=189
M35 VDD 8 10 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6900 $Y=1930 $D=189
M36 13 9 10 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7910 $Y=1960 $D=189
M37 10 9 13 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8390 $Y=1960 $D=189
M38 13 9 10 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8870 $Y=1960 $D=189
M39 22 11 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9390 $Y=2620 $D=189
M40 VDD 12 22 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9710 $Y=2620 $D=189
M41 VDD 13 12 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10270 $Y=1910 $D=189
M42 Q 13 VDD VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10670 $Y=1910 $D=189
M43 VDD 13 Q VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11150 $Y=1910 $D=189
M44 Q 13 VDD VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11630 $Y=1910 $D=189
M45 VDD 13 Q VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12110 $Y=1910 $D=189
M46 Q 13 VDD VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12590 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DFFHQX4TR CK D Q VSS VDD
** N=104 EP=5 IP=0 FDC=41
M0 VSS CK 6 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=770 $D=97
M1 9 CK VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=830 $D=97
M2 VSS D 7 VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1830 $Y=870 $D=97
M3 11 6 VSS VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2430 $Y=590 $D=97
M4 15 9 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3450 $Y=710 $D=97
M5 8 7 15 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3770 $Y=710 $D=97
M6 17 7 8 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4410 $Y=500 $D=97
M7 VSS 9 17 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4730 $Y=500 $D=97
M8 20 11 8 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5610 $Y=900 $D=97
M9 VSS 10 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5930 $Y=900 $D=97
M10 10 8 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6330 $Y=390 $D=97
M11 VSS 8 10 VSS nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6810 $Y=670 $D=97
M12 13 11 10 VSS nfet L=1.2e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7820 $Y=600 $D=97
M13 10 11 13 VSS nfet L=1.2e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8300 $Y=600 $D=97
M14 21 9 13 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9280 $Y=600 $D=97
M15 VSS 12 21 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9620 $Y=600 $D=97
M16 VSS 13 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10180 $Y=1110 $D=97
M17 Q 13 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10580 $Y=390 $D=97
M18 VSS 13 Q VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11060 $Y=390 $D=97
M19 VDD CK 6 VDD pfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M20 14 CK VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=1910 $D=189
M21 9 11 14 VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1170 $Y=1910 $D=189
M22 VDD D 7 VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1990 $Y=1910 $D=189
M23 11 6 VDD VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2430 $Y=1910 $D=189
M24 VDD 6 11 VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2910 $Y=1910 $D=189
M25 16 7 8 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3770 $Y=2140 $D=189
M26 VDD 11 16 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4090 $Y=2140 $D=189
M27 18 11 VDD VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4650 $Y=2140 $D=189
M28 8 7 18 VDD pfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4970 $Y=2140 $D=189
M29 19 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5500 $Y=1930 $D=189
M30 VDD 10 19 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5850 $Y=1930 $D=189
M31 10 8 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6330 $Y=1930 $D=189
M32 VDD 8 10 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6810 $Y=1930 $D=189
M33 13 9 10 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7820 $Y=1960 $D=189
M34 10 9 13 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8300 $Y=1960 $D=189
M35 13 9 10 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8780 $Y=1960 $D=189
M36 22 11 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9300 $Y=2620 $D=189
M37 VDD 12 22 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9620 $Y=2620 $D=189
M38 VDD 13 12 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10180 $Y=1910 $D=189
M39 Q 13 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10580 $Y=1910 $D=189
M40 VDD 13 Q VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11060 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DFFSX2TR D CK SN VSS Q VDD QN
** N=88 EP=7 IP=0 FDC=31
M0 16 D VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=950 $D=97
M1 8 9 16 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=650 $Y=950 $D=97
M2 18 11 8 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1210 $Y=930 $D=97
M3 VSS 10 18 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1530 $Y=930 $D=97
M4 9 CK VSS VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=530 $D=97
M5 12 8 10 VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2490 $Y=1010 $D=97
M6 11 9 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3350 $Y=1020 $D=97
M7 13 11 10 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4370 $Y=700 $D=97
M8 20 9 13 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4930 $Y=1050 $D=97
M9 12 14 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5250 $Y=1050 $D=97
M10 VSS SN 12 VSS nfet L=1.2e-07 W=4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5690 $Y=850 $D=97
M11 14 13 VSS VSS nfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6130 $Y=990 $D=97
M12 15 14 VSS VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6450 $Y=390 $D=97
M13 VSS 14 Q VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7310 $Y=390 $D=97
M14 QN 15 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=390 $D=97
M15 17 D VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=2180 $D=189
M16 8 11 17 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=650 $Y=2180 $D=189
M17 19 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1210 $Y=2180 $D=189
M18 VDD 10 19 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1530 $Y=2180 $D=189
M19 9 CK VDD VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=2470 $D=189
M20 VDD 8 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2580 $Y=1910 $D=189
M21 11 9 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3020 $Y=2110 $D=189
M22 13 9 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4040 $Y=1910 $D=189
M23 VDD SN 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4120 $Y=2850 $D=189
M24 13 SN VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4680 $Y=2610 $D=189
M25 21 11 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5240 $Y=2610 $D=189
M26 VDD 14 21 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5560 $Y=2610 $D=189
M27 14 13 VDD VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6390 $Y=1910 $D=189
M28 15 14 VDD VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6430 $Y=2910 $D=189
M29 VDD 14 Q VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7310 $Y=1930 $D=189
M30 QN 15 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=1930 $D=189
.ENDS
***************************************
.SUBCKT ICV_265
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ADDFHX2TR A B CI CO VSS VDD S
** N=111 EP=7 IP=0 FDC=46
M0 9 A VSS VSS nfet L=1.2e-07 W=5.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=560 $D=97
M1 VSS A 9 VSS nfet L=1.2e-07 W=5.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=560 $D=97
M2 8 A VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=670 $D=97
M3 VSS 8 10 VSS nfet L=1.2e-07 W=5.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2370 $Y=620 $D=97
M4 10 8 VSS VSS nfet L=1.2e-07 W=5.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2930 $Y=620 $D=97
M5 11 B 10 VSS nfet L=1.2e-07 W=5.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3410 $Y=620 $D=97
M6 10 B 11 VSS nfet L=1.2e-07 W=5.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3970 $Y=620 $D=97
M7 11 12 9 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4910 $Y=710 $D=97
M8 9 12 11 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5390 $Y=710 $D=97
M9 14 B 9 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5870 $Y=710 $D=97
M10 9 B 14 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6350 $Y=710 $D=97
M11 10 12 14 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7390 $Y=760 $D=97
M12 14 12 10 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7950 $Y=760 $D=97
M13 VSS B 12 VSS nfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9140 $Y=480 $D=97
M14 12 B VSS VSS nfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9800 $Y=480 $D=97
M15 13 11 12 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10280 $Y=640 $D=97
M16 16 14 13 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10800 $Y=710 $D=97
M17 17 11 16 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11280 $Y=710 $D=97
M18 15 14 17 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11760 $Y=710 $D=97
M19 VSS 16 15 VSS nfet L=1.2e-07 W=6.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12240 $Y=650 $D=97
M20 16 CI VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12800 $Y=390 $D=97
M21 VSS 13 CO VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=13760 $Y=390 $D=97
M22 S 17 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=14240 $Y=390 $D=97
M23 9 A VDD VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M24 VDD A 9 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=1910 $D=189
M25 8 A VDD VDD pfet L=1.2e-07 W=6.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=1910 $D=189
M26 VDD 8 10 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2170 $Y=2240 $D=189
M27 10 8 VDD VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2650 $Y=2240 $D=189
M28 11 12 10 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3130 $Y=2240 $D=189
M29 10 12 11 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3610 $Y=2240 $D=189
M30 11 B 9 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4550 $Y=1920 $D=189
M31 9 B 11 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5030 $Y=1920 $D=189
M32 14 12 9 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5510 $Y=1920 $D=189
M33 9 12 14 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5990 $Y=1920 $D=189
M34 14 B 10 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6850 $Y=2240 $D=189
M35 10 B 14 VDD pfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7330 $Y=2240 $D=189
M36 VDD B 12 VDD pfet L=1.2e-07 W=1.06e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8390 $Y=2150 $D=189
M37 12 B VDD VDD pfet L=1.2e-07 W=1.06e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9140 $Y=2150 $D=189
M38 13 14 12 VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9950 $Y=2260 $D=189
M39 16 11 13 VDD pfet L=1.2e-07 W=9.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=10610 $Y=1950 $D=189
M40 17 14 16 VDD pfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11120 $Y=2290 $D=189
M41 15 11 17 VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=11600 $Y=2090 $D=189
M42 VDD 16 15 VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12160 $Y=2090 $D=189
M43 16 CI VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=12720 $Y=1910 $D=189
M44 VDD 13 CO VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=13760 $Y=1910 $D=189
M45 S 17 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=14240 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_263
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_264
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ADDFX2TR B A CI CO VSS VDD S
** N=88 EP=7 IP=0 FDC=29
M0 VSS B 10 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=390 $D=97
M1 8 10 VSS VSS nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=670 $D=97
M2 12 9 8 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=770 $D=97
M3 9 8 12 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=950 $D=97
M4 VSS A 9 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2450 $Y=750 $D=97
M5 9 A VSS VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2890 $Y=950 $D=97
M6 13 10 9 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3370 $Y=950 $D=97
M7 10 9 13 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3860 $Y=850 $D=97
M8 14 13 10 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4750 $Y=1030 $D=97
M9 11 12 14 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5230 $Y=1030 $D=97
M10 VSS CI 11 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5750 $Y=730 $D=97
M11 15 CI 12 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6610 $Y=790 $D=97
M12 13 11 15 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7090 $Y=790 $D=97
M13 VSS 14 CO VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8090 $Y=390 $D=97
M14 S 15 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8570 $Y=390 $D=97
M15 VDD B 10 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M16 8 10 VDD VDD pfet L=1.2e-07 W=9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=1910 $D=189
M17 13 9 8 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=1910 $D=189
M18 9 8 13 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=1910 $D=189
M19 VDD A 9 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2550 $Y=1910 $D=189
M20 12 10 9 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3370 $Y=1990 $D=189
M21 10 9 12 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3860 $Y=1990 $D=189
M22 14 12 10 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4340 $Y=2450 $D=189
M23 11 13 14 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4820 $Y=2450 $D=189
M24 VDD CI 11 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5400 $Y=3030 $D=189
M25 15 11 12 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6510 $Y=1910 $D=189
M26 13 CI 15 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6990 $Y=2130 $D=189
M27 VDD 14 CO VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8090 $Y=1910 $D=189
M28 S 15 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8570 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT NOR2X2TR A B Y VSS VDD
** N=26 EP=5 IP=0 FDC=6
M0 Y A VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=390 $D=97
M1 VSS B Y VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1340 $Y=390 $D=97
M2 6 B VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=430 $Y=2030 $D=189
M3 Y A 6 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=750 $Y=2030 $D=189
M4 7 A Y VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1230 $Y=2030 $D=189
M5 VDD B 7 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1550 $Y=2030 $D=189
.ENDS
***************************************
.SUBCKT DFFSX1TR D CK SN VSS Q VDD
** N=83 EP=6 IP=0 FDC=31
M0 16 D VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=950 $D=97
M1 7 8 16 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=650 $Y=950 $D=97
M2 18 10 7 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1210 $Y=930 $D=97
M3 VSS 9 18 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1530 $Y=930 $D=97
M4 8 CK VSS VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=530 $D=97
M5 11 7 9 VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2580 $Y=1010 $D=97
M6 10 8 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3440 $Y=1020 $D=97
M7 12 10 9 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4460 $Y=700 $D=97
M8 20 8 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5020 $Y=1110 $D=97
M9 11 13 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5340 $Y=1110 $D=97
M10 VSS SN 11 VSS nfet L=1.2e-07 W=4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5840 $Y=480 $D=97
M11 13 12 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6280 $Y=1110 $D=97
M12 14 13 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6600 $Y=390 $D=97
M13 VSS 13 Q VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7370 $Y=850 $D=97
M14 QN 14 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=850 $D=97
M15 17 D VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=330 $Y=2180 $D=189
M16 7 10 17 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=650 $Y=2180 $D=189
M17 19 8 7 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1210 $Y=2180 $D=189
M18 VDD 9 19 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1530 $Y=2180 $D=189
M19 8 CK VDD VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=2470 $D=189
M20 VDD 7 9 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2580 $Y=1910 $D=189
M21 10 8 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3020 $Y=2110 $D=189
M22 12 8 9 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4040 $Y=1910 $D=189
M23 VDD SN 9 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4120 $Y=2850 $D=189
M24 12 SN VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4680 $Y=2610 $D=189
M25 21 10 12 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5240 $Y=2610 $D=189
M26 VDD 13 21 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5560 $Y=2610 $D=189
M27 13 12 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6390 $Y=1910 $D=189
M28 14 13 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6430 $Y=2860 $D=189
M29 VDD 13 Q VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7370 $Y=2340 $D=189
M30 QN 14 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=1940 $D=189
.ENDS
***************************************
.SUBCKT DFFHQX1TR D CK VSS VDD Q
** N=81 EP=5 IP=0 FDC=29
M0 VSS D 7 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1060 $D=97
M1 VSS CK 9 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1480 $Y=860 $D=97
M2 6 CK VSS VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1920 $Y=780 $D=97
M3 VSS 6 11 VSS nfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2810 $Y=500 $D=97
M4 16 9 VSS VSS nfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3260 $Y=650 $D=97
M5 8 7 16 VSS nfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3580 $Y=650 $D=97
M6 18 11 8 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4140 $Y=910 $D=97
M7 VSS 10 18 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4460 $Y=910 $D=97
M8 10 8 VSS VSS nfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4930 $Y=720 $D=97
M9 12 11 10 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5470 $Y=720 $D=97
M10 20 9 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6090 $Y=570 $D=97
M11 VSS 13 20 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6410 $Y=570 $D=97
M12 VSS 12 13 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6970 $Y=1080 $D=97
M13 Q 12 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7470 $Y=820 $D=97
M14 VDD D 7 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1910 $D=189
M15 6 CK VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=1910 $D=189
M16 14 CK VDD VDD pfet L=1.2e-07 W=7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=2370 $D=189
M17 9 11 14 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=2500 $D=189
M18 VDD 6 11 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2490 $Y=1910 $D=189
M19 15 11 VDD VDD pfet L=1.2e-07 W=5.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3050 $Y=1910 $D=189
M20 8 7 15 VDD pfet L=1.2e-07 W=5.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3370 $Y=1910 $D=189
M21 17 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3890 $Y=2110 $D=189
M22 VDD 10 17 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4210 $Y=2110 $D=189
M23 10 8 VDD VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4740 $Y=2110 $D=189
M24 12 9 10 VDD pfet L=1.2e-07 W=9.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5250 $Y=2110 $D=189
M25 19 11 12 VDD pfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5770 $Y=2290 $D=189
M26 VDD 13 19 VDD pfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6090 $Y=2290 $D=189
M27 VDD 12 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7040 $Y=2280 $D=189
M28 Q 12 VDD VDD pfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7440 $Y=2280 $D=189
.ENDS
***************************************
.SUBCKT XOR2X1TR A B Y VDD VSS
** N=30 EP=5 IP=0 FDC=10
M0 VSS A 6 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=1040 $D=97
M1 8 B VSS VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1010 $Y=720 $D=97
M2 Y A 8 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1490 $Y=720 $D=97
M3 7 6 Y VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=710 $D=97
M4 VSS 8 7 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2630 $Y=710 $D=97
M5 VDD A 6 VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=2000 $D=189
M6 8 B VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1010 $Y=2000 $D=189
M7 Y 6 8 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1490 $Y=2000 $D=189
M8 7 A Y VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=2240 $D=189
M9 VDD 8 7 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2630 $Y=2240 $D=189
.ENDS
***************************************
.SUBCKT DFFQX1TR D CK VSS VDD Q
** N=63 EP=5 IP=0 FDC=25
M0 12 D VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=390 $Y=1010 $D=97
M1 6 9 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=710 $Y=1010 $D=97
M2 15 7 6 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1270 $Y=1010 $D=97
M3 VSS 8 15 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1590 $Y=1010 $D=97
M4 9 CK VSS VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2030 $Y=960 $D=97
M5 8 6 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2890 $Y=1090 $D=97
M6 VSS 9 7 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3610 $Y=710 $D=97
M7 10 7 8 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4490 $Y=1110 $D=97
M8 17 9 10 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5150 $Y=1000 $D=97
M9 VSS 11 Q VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5470 $Y=390 $D=97
M10 VSS 11 17 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5470 $Y=1000 $D=97
M11 11 10 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5910 $Y=1110 $D=97
M12 Q 11 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6230 $Y=520 $D=97
M13 13 D VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=390 $Y=2390 $D=189
M14 6 7 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=780 $Y=2390 $D=189
M15 14 9 6 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1260 $Y=2390 $D=189
M16 VDD 8 14 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1580 $Y=2390 $D=189
M17 VDD CK 9 VDD pfet L=1.2e-07 W=3.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2440 $Y=2450 $D=189
M18 8 6 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2890 $Y=2450 $D=189
M19 VDD 9 7 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3780 $Y=1990 $D=189
M20 10 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4640 $Y=2290 $D=189
M21 16 7 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5080 $Y=2290 $D=189
M22 VDD 11 16 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5400 $Y=2290 $D=189
M23 11 10 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5860 $Y=1950 $D=189
M24 Q 11 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6260 $Y=2570 $D=189
.ENDS
***************************************
.SUBCKT NOR2BX1TR AN B VDD Y VSS
** N=25 EP=5 IP=0 FDC=6
M0 VSS AN 6 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1090 $D=97
M1 Y B VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=850 $D=97
M2 VSS 6 Y VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1520 $Y=850 $D=97
M3 VDD AN 6 VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1940 $D=189
M4 7 B VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=1940 $D=189
M5 Y 6 7 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1360 $Y=1940 $D=189
.ENDS
***************************************
.SUBCKT CMPR32X2TR B A C CO VSS VDD S
** N=81 EP=7 IP=0 FDC=29
M0 VSS B 10 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=390 $D=97
M1 8 10 VSS VSS nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=670 $D=97
M2 12 9 8 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=770 $D=97
M3 9 8 12 VSS nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=970 $D=97
M4 VSS A 9 VSS nfet L=1.2e-07 W=5.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2450 $Y=730 $D=97
M5 9 A VSS VSS nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2890 $Y=970 $D=97
M6 14 10 9 VSS nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3410 $Y=970 $D=97
M7 10 9 14 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3890 $Y=770 $D=97
M8 13 14 10 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4570 $Y=1040 $D=97
M9 11 12 13 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5050 $Y=1040 $D=97
M10 VSS C 11 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5570 $Y=390 $D=97
M11 15 C 12 VSS nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6290 $Y=900 $D=97
M12 14 11 15 VSS nfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6770 $Y=900 $D=97
M13 VSS 13 CO VSS nfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7690 $Y=400 $D=97
M14 S 15 VSS VSS nfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8170 $Y=400 $D=97
M15 VDD B 10 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1930 $D=189
M16 8 10 VDD VDD pfet L=1.2e-07 W=9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=1910 $D=189
M17 14 9 8 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1330 $Y=1910 $D=189
M18 9 8 14 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1970 $Y=1910 $D=189
M19 VDD A 9 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2450 $Y=1910 $D=189
M20 12 10 9 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3270 $Y=2030 $D=189
M21 10 9 12 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3750 $Y=2030 $D=189
M22 13 12 10 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4230 $Y=2500 $D=189
M23 11 14 13 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4710 $Y=2500 $D=189
M24 VDD C 11 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5430 $Y=2500 $D=189
M25 15 11 12 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6390 $Y=2240 $D=189
M26 14 C 15 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6870 $Y=2240 $D=189
M27 VDD 13 CO VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7690 $Y=1910 $D=189
M28 S 15 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8170 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT OR2X2TR A B VSS VDD Y
** N=26 EP=5 IP=0 FDC=6
M0 6 A VSS VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=790 $D=97
M1 VSS B 6 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=970 $Y=790 $D=97
M2 Y 6 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=390 $D=97
M3 7 A 6 VDD pfet L=1.2e-07 W=6.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=1910 $D=189
M4 VDD B 7 VDD pfet L=1.2e-07 W=6.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=800 $Y=1910 $D=189
M5 Y 6 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT INVX2TR A VSS VDD Y
** N=14 EP=4 IP=0 FDC=2
M0 Y A VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=520 $Y=390 $D=97
M1 Y A VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=520 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT DFFHQX2TR D CK VDD VSS Q
** N=87 EP=5 IP=0 FDC=31
M0 VSS D 7 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=910 $D=97
M1 VSS CK 9 VSS nfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1520 $Y=710 $D=97
M2 6 CK VSS VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1960 $Y=650 $D=97
M3 VSS 6 11 VSS nfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2900 $Y=650 $D=97
M4 16 9 VSS VSS nfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3420 $Y=390 $D=97
M5 8 7 16 VSS nfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3740 $Y=390 $D=97
M6 18 11 8 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4300 $Y=770 $D=97
M7 VSS 10 18 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4620 $Y=770 $D=97
M8 10 8 VSS VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5580 $Y=410 $D=97
M9 12 11 10 VSS nfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6150 $Y=450 $D=97
M10 19 9 12 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6900 $Y=580 $D=97
M11 VSS 13 19 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7220 $Y=580 $D=97
M12 VSS 12 13 VSS nfet L=1.2e-07 W=1.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=1090 $D=97
M13 Q 12 VSS VSS nfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8270 $Y=390 $D=97
M14 VDD D 7 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=460 $Y=1910 $D=189
M15 6 CK VDD VDD pfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1080 $Y=1750 $D=189
M16 14 CK VDD VDD pfet L=1.2e-07 W=9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1080 $Y=2250 $D=189
M17 9 11 14 VDD pfet L=1.2e-07 W=6.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1480 $Y=2470 $D=189
M18 VDD 6 11 VDD pfet L=1.2e-07 W=1.18e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2400 $Y=1890 $D=189
M19 15 11 VDD VDD pfet L=1.2e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2960 $Y=1890 $D=189
M20 8 7 15 VDD pfet L=1.2e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3280 $Y=1890 $D=189
M21 17 9 8 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3800 $Y=2110 $D=189
M22 VDD 10 17 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4120 $Y=2110 $D=189
M23 10 8 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4560 $Y=2110 $D=189
M24 VDD 8 10 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5040 $Y=2110 $D=189
M25 10 9 12 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5900 $Y=1990 $D=189
M26 12 9 10 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6380 $Y=1990 $D=189
M27 20 11 12 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6900 $Y=2490 $D=189
M28 VDD 13 20 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7220 $Y=2490 $D=189
M29 VDD 12 13 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7870 $Y=1910 $D=189
M30 Q 12 VDD VDD pfet L=1.2e-07 W=1.3e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8270 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ADDFHX1TR A B CI CO VSS VDD S
** N=77 EP=7 IP=0 FDC=32
M0 VSS A 9 VSS nfet L=1.2e-07 W=5.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=730 $D=97
M1 8 A VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=870 $Y=1070 $D=97
M2 10 8 VSS VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1730 $Y=710 $D=97
M3 11 B 10 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2210 $Y=710 $D=97
M4 9 13 11 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2690 $Y=710 $D=97
M5 12 B 9 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3170 $Y=710 $D=97
M6 10 13 12 VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3650 $Y=710 $D=97
M7 13 B VSS VSS nfet L=1.2e-07 W=8.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5260 $Y=390 $D=97
M8 14 11 13 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5800 $Y=850 $D=97
M9 16 12 14 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6280 $Y=850 $D=97
M10 17 11 16 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6760 $Y=850 $D=97
M11 15 12 17 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7240 $Y=850 $D=97
M12 VSS 16 15 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7720 $Y=850 $D=97
M13 16 CI VSS VSS nfet L=1.2e-07 W=5.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=8160 $Y=570 $D=97
M14 VSS 14 CO VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9010 $Y=850 $D=97
M15 S 17 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9450 $Y=850 $D=97
M16 VDD A 9 VDD pfet L=1.2e-07 W=8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=1940 $D=189
M17 8 A VDD VDD pfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=850 $Y=1940 $D=189
M18 10 8 VDD VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1410 $Y=2450 $D=189
M19 11 13 10 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1890 $Y=2170 $D=189
M20 9 B 11 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2370 $Y=2170 $D=189
M21 12 13 9 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2850 $Y=2220 $D=189
M22 10 B 12 VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3330 $Y=2220 $D=189
M23 13 B VDD VDD pfet L=1.2e-07 W=1.14e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4500 $Y=1960 $D=189
M24 14 12 13 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4980 $Y=2420 $D=189
M25 16 11 14 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=5960 $Y=2190 $D=189
M26 17 12 16 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6440 $Y=2190 $D=189
M27 15 11 17 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=6920 $Y=2190 $D=189
M28 VDD 16 15 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7550 $Y=2190 $D=189
M29 16 CI VDD VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7990 $Y=2190 $D=189
M30 VDD 14 CO VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9010 $Y=1910 $D=189
M31 S 17 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=9450 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT INVX4TR A Y VSS VDD
** N=19 EP=4 IP=0 FDC=4
M0 Y A VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=390 $D=97
M1 VSS A Y VSS nfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=530 $D=97
M2 Y A VDD VDD pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=410 $Y=1960 $D=189
M3 VDD A Y VDD pfet L=1.2e-07 W=1.1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=890 $Y=1960 $D=189
.ENDS
***************************************
.SUBCKT OAI2BB1X1TR A1N A0N B0 VSS Y VDD
** N=26 EP=6 IP=0 FDC=8
M0 8 A1N 7 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=560 $Y=970 $D=97
M1 VSS A0N 8 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=880 $Y=970 $D=97
M2 9 B0 VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1440 $Y=650 $D=97
M3 Y 7 9 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1760 $Y=650 $D=97
M4 7 A1N VDD VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=1970 $D=189
M5 VDD A0N 7 VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=940 $Y=1970 $D=189
M6 Y B0 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1400 $Y=1970 $D=189
M7 VDD 7 Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1840 $Y=1970 $D=189
.ENDS
***************************************
.SUBCKT ADDHX1TR S B A CO VDD VSS
** N=47 EP=6 IP=0 FDC=18
M0 VSS 9 8 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=440 $Y=390 $D=97
M1 7 B VSS VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1000 $Y=830 $D=97
M2 S 7 8 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2180 $Y=390 $D=97
M3 9 B S VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2660 $Y=390 $D=97
M4 VSS A 9 VSS nfet L=1.2e-07 W=8.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3140 $Y=390 $D=97
M5 11 A VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3700 $Y=390 $D=97
M6 9 A VSS VSS nfet L=1.2e-07 W=4.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3700 $Y=810 $D=97
M7 10 B 11 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4170 $Y=390 $D=97
M8 VSS 10 CO VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4750 $Y=850 $D=97
M9 VDD 9 8 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=440 $Y=1930 $D=189
M10 7 B VDD VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=990 $Y=2250 $D=189
M11 S B 8 VDD pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1940 $Y=1970 $D=189
M12 9 7 S VDD pfet L=1.2e-07 W=1.24e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2420 $Y=1970 $D=189
M13 VDD A 9 VDD pfet L=1.2e-07 W=1.15e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3140 $Y=2060 $D=189
M14 9 A VDD VDD pfet L=1.2e-07 W=6.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3700 $Y=2060 $D=189
M15 10 A VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3700 $Y=2870 $D=189
M16 VDD B 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4310 $Y=2870 $D=189
M17 VDD 10 CO VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4750 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ADDHXLTR S A B VSS VDD CO
** N=48 EP=6 IP=0 FDC=16
M0 VSS 9 7 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=500 $Y=950 $D=97
M1 8 B VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=940 $Y=990 $D=97
M2 S 8 7 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1570 $Y=410 $D=97
M3 9 B S VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2110 $Y=820 $D=97
M4 VSS A 9 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2660 $Y=900 $D=97
M5 11 A VSS VSS nfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3270 $Y=880 $D=97
M6 10 B 11 VSS nfet L=1.2e-07 W=2.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3590 $Y=880 $D=97
M7 CO 10 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4220 $Y=420 $D=97
M8 VDD 9 7 VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=500 $Y=2250 $D=189
M9 8 B VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=940 $Y=2250 $D=189
M10 S B 7 VDD pfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1850 $Y=2250 $D=189
M11 9 8 S VDD pfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2350 $Y=2060 $D=189
M12 VDD A 9 VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2830 $Y=2060 $D=189
M13 10 A VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3270 $Y=2060 $D=189
M14 VDD B 10 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3830 $Y=2060 $D=189
M15 CO 10 VDD VDD pfet L=1.2e-07 W=4.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=4270 $Y=2060 $D=189
.ENDS
***************************************
.SUBCKT NAND2BX1TR AN B VSS Y VDD
** N=22 EP=5 IP=0 FDC=6
M0 VSS AN 6 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=560 $Y=1050 $D=97
M1 7 B VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1100 $Y=650 $D=97
M2 Y 6 7 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1420 $Y=650 $D=97
M3 VDD AN 6 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=2040 $D=189
M4 Y B VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=940 $Y=2040 $D=189
M5 VDD 6 Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1420 $Y=2040 $D=189
.ENDS
***************************************
.SUBCKT ICV_268 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=6
X0 1 2 3 4 5 AND2X2TR $T=1200 0 0 0 $X=860 $Y=-280
.ENDS
***************************************
.SUBCKT OAI21X2TR A0 A1 VSS B0 Y VDD
** N=45 EP=6 IP=0 FDC=12
M0 VSS A1 7 VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=480 $Y=700 $D=97
M1 7 A0 VSS VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=700 $D=97
M2 VSS A0 7 VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1520 $Y=700 $D=97
M3 7 A1 VSS VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2080 $Y=700 $D=97
M4 Y B0 7 VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2560 $Y=700 $D=97
M5 7 B0 Y VSS nfet L=1.2e-07 W=6.1e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3040 $Y=700 $D=97
M6 8 A1 VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=720 $Y=1910 $D=189
M7 Y A0 8 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1040 $Y=1910 $D=189
M8 9 A0 Y VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1520 $Y=1910 $D=189
M9 VDD A1 9 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1840 $Y=1910 $D=189
M10 Y B0 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2520 $Y=1910 $D=189
M11 VDD B0 Y VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=3000 $Y=1910 $D=189
.ENDS
***************************************
.SUBCKT ICV_269 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=6
X1 3 4 2 1 5 AND2X2TR $T=1600 0 0 0 $X=1260 $Y=-280
.ENDS
***************************************
.SUBCKT NAND2X2TR VSS A B Y VDD
** N=26 EP=5 IP=0 FDC=6
M0 6 B VSS VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=360 $Y=670 $D=97
M1 Y A 6 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=680 $Y=670 $D=97
M2 7 A Y VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1160 $Y=670 $D=97
M3 VSS B 7 VSS nfet L=1.2e-07 W=6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1480 $Y=670 $D=97
M4 Y A VDD VDD pfet L=1.2e-07 W=1.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=950 $Y=1950 $D=189
M5 VDD B Y VDD pfet L=1.2e-07 W=1.26e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1430 $Y=1950 $D=189
.ENDS
***************************************
.SUBCKT XNOR2X1TR B A Y VDD VSS
** N=31 EP=5 IP=0 FDC=10
M0 VSS A 6 VSS nfet L=1.2e-07 W=2.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=450 $Y=1090 $D=97
M1 8 B VSS VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=970 $Y=750 $D=97
M2 Y 6 8 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1450 $Y=750 $D=97
M3 7 A Y VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1930 $Y=750 $D=97
M4 VSS 8 7 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2570 $Y=750 $D=97
M5 VDD A 6 VDD pfet L=1.2e-07 W=3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=2170 $D=189
M6 8 B VDD VDD pfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=950 $Y=2170 $D=189
M7 Y A 8 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1430 $Y=2290 $D=189
M8 7 6 Y VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1910 $Y=2100 $D=189
M9 VDD 8 7 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=2570 $Y=2100 $D=189
.ENDS
***************************************
.SUBCKT ICV_1 VDD VSS clk signature<0> signature<4> signature<5> signature<7> signature<8> signature<9> signature<13> signature<15> reset signature<2> signature<6> signature<1> signature<3> signature<10> signature<11> signature<12> signature<14>
** N=5433 EP=20 IP=3332 FDC=7185
M0 2201 reset VSS VSS nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43500 $Y=131880 $D=97
M1 VSS reset 2201 VSS nfet L=1.2e-07 W=4.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43980 $Y=131880 $D=97
M2 2581 2144 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=69360 $Y=102890 $D=97
M3 VSS 4351 2581 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=69840 $Y=102890 $D=97
M4 4351 2180 VSS VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=70400 $Y=102910 $D=97
M5 VSS 4357 3828 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72210 $Y=52490 $D=97
M6 4356 4364 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72410 $Y=66890 $D=97
M7 VSS 4364 4356 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72890 $Y=66890 $D=97
M8 VSS 3848 4366 VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73200 $Y=52520 $D=97
M9 4355 3847 VSS VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73450 $Y=66890 $D=97
M10 4366 3848 VSS VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73680 $Y=52520 $D=97
M11 VSS 3848 4366 VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74160 $Y=52520 $D=97
M12 4356 4355 2584 VSS nfet L=1.2e-07 W=8.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74550 $Y=66980 $D=97
M13 4463 3848 VSS VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74600 $Y=52520 $D=97
M14 4357 2585 4463 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74920 $Y=52520 $D=97
M15 2584 4355 4356 VSS nfet L=1.2e-07 W=8.3e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75030 $Y=66980 $D=97
M16 VSS 2607 4367 VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75420 $Y=88490 $D=97
M17 4364 3847 2584 VSS nfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75510 $Y=66930 $D=97
M18 4358 4367 VSS VSS nfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75860 $Y=88490 $D=97
M19 2584 3847 4364 VSS nfet L=1.2e-07 W=8.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75990 $Y=66930 $D=97
M20 4366 2585 2255 VSS nfet L=1.2e-07 W=8.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76040 $Y=52520 $D=97
M21 4370 4361 4358 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76340 $Y=88490 $D=97
M22 2255 2585 4366 VSS nfet L=1.2e-07 W=8.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76520 $Y=52520 $D=97
M23 4464 3847 4363 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76930 $Y=66920 $D=97
M24 4361 4358 4370 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76980 $Y=88490 $D=97
M25 4365 4362 2255 VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77000 $Y=52550 $D=97
M26 VSS 2580 4464 VSS nfet L=1.2e-07 W=4.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77250 $Y=66920 $D=97
M27 VSS 2608 4361 VSS nfet L=1.2e-07 W=5.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77460 $Y=88490 $D=97
M28 2255 4362 4365 VSS nfet L=1.2e-07 W=8.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77480 $Y=52550 $D=97
M29 4364 2580 VSS VSS nfet L=1.2e-07 W=8.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77690 $Y=66920 $D=97
M30 4361 2608 VSS VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77900 $Y=88490 $D=97
M31 VSS 2580 4364 VSS nfet L=1.2e-07 W=8.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78170 $Y=66920 $D=97
M32 4372 4367 4361 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78380 $Y=88490 $D=97
M33 VSS 2585 4362 VSS nfet L=1.2e-07 W=7.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78660 $Y=52670 $D=97
M34 4364 2580 VSS VSS nfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78730 $Y=66920 $D=97
M35 4367 4361 4372 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78860 $Y=88490 $D=97
M36 4365 4366 VSS VSS nfet L=1.2e-07 W=8.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79180 $Y=52520 $D=97
M37 VSS 4366 4365 VSS nfet L=1.2e-07 W=8.9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79660 $Y=52520 $D=97
M38 2616 4363 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79670 $Y=66890 $D=97
M39 4373 4372 4367 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79760 $Y=88410 $D=97
M40 4368 4370 4373 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=80240 $Y=88410 $D=97
M41 VSS 3881 4368 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=80760 $Y=88710 $D=97
M42 4374 3881 4370 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=81620 $Y=88700 $D=97
M43 4372 4368 4374 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=82100 $Y=88700 $D=97
M44 VSS 4373 2216 VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=83100 $Y=88490 $D=97
M45 2629 4374 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=83580 $Y=88490 $D=97
M46 4465 2648 4377 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87090 $Y=59920 $D=97
M47 VSS 2593 4465 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87410 $Y=59920 $D=97
M48 2689 4377 VSS VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87970 $Y=59690 $D=97
M49 4387 2676 VSS VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=95770 $Y=119360 $D=97
M50 VSS 2676 4387 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=96250 $Y=119360 $D=97
M51 4385 4387 VSS VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=96690 $Y=119360 $D=97
M52 VSS 4387 4385 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=97230 $Y=119360 $D=97
M53 4383 3985 VSS VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=97670 $Y=119470 $D=97
M54 2698 2691 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=98370 $Y=18870 $D=97
M55 4385 4383 2312 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=98630 $Y=119340 $D=97
M56 2312 4383 4385 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99110 $Y=119340 $D=97
M57 4391 2649 VSS VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99430 $Y=11360 $D=97
M58 4387 3985 2312 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99590 $Y=119250 $D=97
M59 VSS 2649 4391 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99910 $Y=11360 $D=97
M60 2312 3985 4387 VSS nfet L=1.2e-07 W=5.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100070 $Y=119250 $D=97
M61 4389 4391 VSS VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100350 $Y=11360 $D=97
M62 VSS 4391 4389 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100830 $Y=11360 $D=97
M63 4388 2693 VSS VSS nfet L=1.2e-07 W=4.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=101270 $Y=11310 $D=97
M64 4389 2693 3996 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=102230 $Y=11200 $D=97
M65 3996 2693 4389 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=102710 $Y=11200 $D=97
M66 4391 4388 3996 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=103190 $Y=11200 $D=97
M67 3996 4388 4391 VSS nfet L=1.2e-07 W=5.5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=103670 $Y=11200 $D=97
M68 4466 4049 VSS VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=110480 $Y=68790 $D=97
M69 4467 2744 4466 VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=110800 $Y=68790 $D=97
M70 4064 2748 4467 VSS nfet L=1.2e-07 W=7.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=111120 $Y=68790 $D=97
M71 4468 4090 VSS VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=115860 $Y=83520 $D=97
M72 4402 2766 4468 VSS nfet L=1.2e-07 W=2.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=116180 $Y=83520 $D=97
M73 VSS 4103 4402 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=116740 $Y=83560 $D=97
M74 4118 4402 VSS VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=117270 $Y=83450 $D=97
M75 2759 4407 VSS VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=123420 $Y=103490 $D=97
M76 VSS 4407 2759 VSS nfet L=1.2e-07 W=3.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=123900 $Y=103490 $D=97
M77 VSS 4409 4407 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=124220 $Y=102890 $D=97
M78 4469 4407 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=124660 $Y=103000 $D=97
M79 2759 4407 VSS VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=124660 $Y=103530 $D=97
M80 4409 4414 4469 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=125010 $Y=103000 $D=97
M81 4413 4411 4409 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=125650 $Y=102890 $D=97
M82 4411 4414 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=126510 $Y=103290 $D=97
M83 VSS 4415 4413 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=127190 $Y=102910 $D=97
M84 VSS 2202 4414 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=128050 $Y=102960 $D=97
M85 4471 4413 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=128490 $Y=102990 $D=97
M86 4415 4411 4471 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=128810 $Y=102990 $D=97
M87 4474 4414 4415 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=129370 $Y=102990 $D=97
M88 VSS 2810 4474 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=129690 $Y=102990 $D=97
M89 2812 4420 VSS VSS nfet L=1.2e-07 W=9.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=134610 $Y=90190 $D=97
M90 VSS 4420 2812 VSS nfet L=1.2e-07 W=4.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=135090 $Y=90190 $D=97
M91 VSS 4421 4420 VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=135820 $Y=90750 $D=97
M92 2812 4420 VSS VSS nfet L=1.2e-07 W=3.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=136260 $Y=90190 $D=97
M93 4475 4420 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=136260 $Y=90860 $D=97
M94 4421 4426 4475 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=136610 $Y=90860 $D=97
M95 4425 4423 4421 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=137250 $Y=90910 $D=97
M96 4423 4426 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=138110 $Y=90510 $D=97
M97 VSS 4427 4425 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=138820 $Y=90890 $D=97
M98 VSS 2202 4426 VSS nfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=139680 $Y=90760 $D=97
M99 4477 4425 VSS VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=140120 $Y=90810 $D=97
M100 4427 4423 4477 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=140440 $Y=90810 $D=97
M101 4479 4426 4427 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=141000 $Y=90810 $D=97
M102 VSS 2861 4479 VSS nfet L=1.2e-07 W=2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=141320 $Y=90810 $D=97
M103 2201 reset VDD VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43500 $Y=129820 $D=189
M104 VDD reset 2201 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=43980 $Y=129820 $D=189
M105 4461 2144 VDD VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=69200 $Y=101260 $D=189
M106 2581 4351 4461 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=69520 $Y=101260 $D=189
M107 4462 4351 2581 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=70000 $Y=101260 $D=189
M108 VDD 2144 4462 VDD pfet L=1.2e-07 W=8.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=70320 $Y=101260 $D=189
M109 4351 2180 VDD VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=70800 $Y=101480 $D=189
M110 VDD 4357 3828 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72210 $Y=50610 $D=189
M111 4356 4364 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72410 $Y=64990 $D=189
M112 VDD 4364 4356 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=72890 $Y=64990 $D=189
M113 VDD 3848 4366 VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73200 $Y=50660 $D=189
M114 4355 3847 VDD VDD pfet L=1.2e-07 W=1.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73450 $Y=65250 $D=189
M115 4366 3848 VDD VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=73680 $Y=50660 $D=189
M116 VDD 3848 4366 VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74160 $Y=50660 $D=189
M117 4356 3847 2584 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74390 $Y=64990 $D=189
M118 4357 3848 VDD VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74600 $Y=51360 $D=189
M119 2584 3847 4356 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=74870 $Y=64990 $D=189
M120 VDD 2585 4357 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75140 $Y=51360 $D=189
M121 4364 4355 2584 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75400 $Y=64990 $D=189
M122 VDD 2607 4367 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75420 $Y=86610 $D=189
M123 4358 4367 VDD VDD pfet L=1.2e-07 W=9e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75860 $Y=86990 $D=189
M124 2584 4355 4364 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=75880 $Y=64990 $D=189
M125 4366 4362 2255 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76240 $Y=50590 $D=189
M126 4372 4361 4358 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76340 $Y=87130 $D=189
M127 2255 4362 4366 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76720 $Y=50590 $D=189
M128 4363 3847 VDD VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76740 $Y=65740 $D=189
M129 4361 4358 4372 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=76980 $Y=87390 $D=189
M130 4365 2585 2255 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77240 $Y=50590 $D=189
M131 VDD 2580 4363 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77250 $Y=65740 $D=189
M132 VDD 2608 4361 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77560 $Y=86610 $D=189
M133 4364 2580 VDD VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77660 $Y=65040 $D=189
M134 2255 2585 4365 VDD pfet L=1.2e-07 W=1.27e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=77720 $Y=50590 $D=189
M135 VDD 2580 4364 VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78140 $Y=65040 $D=189
M136 4370 4367 4361 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78380 $Y=87310 $D=189
M137 4364 2580 VDD VDD pfet L=1.2e-07 W=1.2e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78620 $Y=65040 $D=189
M138 VDD 2585 4362 VDD pfet L=1.2e-07 W=1e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78740 $Y=50910 $D=189
M139 4367 4361 4370 VDD pfet L=1.2e-07 W=7.6e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=78860 $Y=87050 $D=189
M140 4365 4366 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79180 $Y=50610 $D=189
M141 4373 4370 4367 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79340 $Y=86900 $D=189
M142 2616 4363 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79640 $Y=65010 $D=189
M143 VDD 4366 4365 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79660 $Y=50610 $D=189
M144 4368 4372 4373 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=79820 $Y=86900 $D=189
M145 4368 3881 VDD VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=80370 $Y=86700 $D=189
M146 4374 4368 4370 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=81540 $Y=87390 $D=189
M147 4372 3881 4374 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=82020 $Y=87220 $D=189
M148 VDD 4373 2216 VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=83140 $Y=87250 $D=189
M149 2629 4374 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=83580 $Y=87250 $D=189
M150 4377 2648 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87010 $Y=58260 $D=189
M151 VDD 2593 4377 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87490 $Y=58260 $D=189
M152 2689 4377 VDD VDD pfet L=1.2e-07 W=9.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=87970 $Y=58120 $D=189
M153 VDD 4377 2689 VDD pfet L=1.2e-07 W=9.7e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=88450 $Y=58120 $D=189
M154 4387 2676 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=95770 $Y=120630 $D=189
M155 VDD 2676 4387 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=96250 $Y=120630 $D=189
M156 4385 4387 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=96690 $Y=120630 $D=189
M157 VDD 4387 4385 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=97230 $Y=120630 $D=189
M158 4383 3985 VDD VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=97670 $Y=120630 $D=189
M159 2698 2691 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=98370 $Y=19710 $D=189
M160 4385 3985 2312 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=98630 $Y=120770 $D=189
M161 2312 3985 4385 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99110 $Y=120770 $D=189
M162 4391 2649 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99430 $Y=12510 $D=189
M163 4387 4383 2312 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99590 $Y=120770 $D=189
M164 VDD 2649 4391 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=99910 $Y=12510 $D=189
M165 2312 4383 4387 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100070 $Y=120770 $D=189
M166 4389 4391 VDD VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100350 $Y=12510 $D=189
M167 VDD 4391 4389 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=100830 $Y=12510 $D=189
M168 4388 2693 VDD VDD pfet L=1.2e-07 W=6.2e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=101270 $Y=12510 $D=189
M169 4389 4388 3996 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=102230 $Y=12710 $D=189
M170 3996 4388 4389 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=102710 $Y=12710 $D=189
M171 4391 2693 3996 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=103190 $Y=12730 $D=189
M172 3996 2693 4391 VDD pfet L=1.2e-07 W=7.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=103670 $Y=12730 $D=189
M173 4064 4049 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=110240 $Y=70250 $D=189
M174 VDD 2744 4064 VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=110720 $Y=70250 $D=189
M175 4064 2748 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=111240 $Y=70250 $D=189
M176 VDD 4090 4399 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=115820 $Y=84510 $D=189
M177 4399 2766 VDD VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=116340 $Y=84510 $D=189
M178 4402 4103 4399 VDD pfet L=1.2e-07 W=3.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=116820 $Y=84510 $D=189
M179 VDD 4402 4118 VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=116830 $Y=85640 $D=189
M180 2759 4407 VDD VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=123420 $Y=100990 $D=189
M181 VDD 4407 2759 VDD pfet L=1.2e-07 W=6.4e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=123900 $Y=100990 $D=189
M182 VDD 4409 4407 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=124220 $Y=101970 $D=189
M183 4470 4407 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=124680 $Y=101630 $D=189
M184 4409 4411 4470 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=125000 $Y=101630 $D=189
M185 4413 4414 4409 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=125440 $Y=101630 $D=189
M186 4411 4414 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=126300 $Y=101930 $D=189
M187 VDD 4415 4413 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=127190 $Y=101470 $D=189
M188 4414 2202 VDD VDD pfet L=1.2e-07 W=3.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=127640 $Y=101370 $D=189
M189 4472 4413 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=128500 $Y=101530 $D=189
M190 4415 4414 4472 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=128820 $Y=101530 $D=189
M191 4473 4411 4415 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=129300 $Y=101530 $D=189
M192 VDD 2810 4473 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=129690 $Y=101530 $D=189
M193 2812 4420 VDD VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=134610 $Y=91730 $D=189
M194 VDD 4420 2812 VDD pfet L=1.2e-07 W=1.28e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=135090 $Y=91730 $D=189
M195 VDD 4421 4420 VDD pfet L=1.2e-07 W=5e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=135940 $Y=91750 $D=189
M196 4476 4420 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=136390 $Y=92090 $D=189
M197 4421 4423 4476 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=136710 $Y=92090 $D=189
M198 4425 4426 4421 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=137150 $Y=92090 $D=189
M199 4423 4426 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=138010 $Y=91790 $D=189
M200 VDD 4427 4425 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=138900 $Y=92250 $D=189
M201 4426 2202 VDD VDD pfet L=1.2e-07 W=3.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=139340 $Y=92250 $D=189
M202 4478 4425 VDD VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=140200 $Y=92190 $D=189
M203 4427 4426 4478 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=140520 $Y=92190 $D=189
M204 4480 4423 4427 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=141000 $Y=92190 $D=189
M205 VDD 2861 4480 VDD pfet L=1.2e-07 W=2.8e-07 m=1 par=1 nf=1 ngcon=1 psp=0 $X=141320 $Y=92190 $D=189
X356 2808 VSS VDD 2810 CLKBUFX2TR $T=126200 82600 0 0 $X=125860 $Y=82320
X357 2179 VSS VDD 2861 CLKBUFX2TR $T=138600 39400 0 0 $X=138260 $Y=39120
X415 clk 2442 VDD VSS CLKINVX8TR $T=9800 17800 0 180 $X=6660 $Y=13800
X416 2055 2172 VSS VDD CLKINVX20TR $T=51400 68200 0 0 $X=51060 $Y=67920
X417 2172 2202 VSS VDD CLKINVX20TR $T=103800 104200 0 180 $X=97860 $Y=100200
X418 2172 2305 VSS VDD CLKINVX20TR $T=99000 68200 0 0 $X=98660 $Y=67920
X442 VSS VDD 2690 3981 INVX1TR $T=97400 111400 0 0 $X=97060 $Y=111120
X443 VSS VDD 2343 4104 INVX1TR $T=115800 53800 0 0 $X=115460 $Y=53520
X491 2592 2180 VDD VSS 2570 AND2X2TR $T=70600 53800 1 180 $X=68260 $Y=53520
X492 2630 2642 VDD VSS 2702 AND2X2TR $T=87800 17800 1 0 $X=87460 $Y=13800
X493 2661 2666 VDD VSS 2715 AND2X2TR $T=101800 118600 1 0 $X=101460 $Y=114600
X494 2718 2734 VDD VSS 2741 AND2X2TR $T=107800 32200 1 0 $X=107460 $Y=28200
X495 2755 2759 VDD VSS 2763 AND2X2TR $T=113800 111400 0 0 $X=113460 $Y=111120
X496 4087 2749 VDD VSS 2788 AND2X2TR $T=115000 89800 1 0 $X=114660 $Y=85800
X497 4113 2808 VDD VSS 2792 AND2X2TR $T=117800 10600 0 0 $X=117460 $Y=10320
X498 2753 2759 VDD VSS 2794 AND2X2TR $T=117800 111400 1 0 $X=117460 $Y=107400
X499 2796 2808 VDD VSS 2769 AND2X2TR $T=121000 25000 1 180 $X=118660 $Y=24720
X500 2798 2364 VDD VSS 4154 AND2X2TR $T=120200 32200 0 0 $X=119860 $Y=31920
X501 2792 2716 VDD VSS 4141 AND2X2TR $T=120600 10600 0 0 $X=120260 $Y=10320
X502 4137 2808 VDD VSS 4150 AND2X2TR $T=121400 17800 1 0 $X=121060 $Y=13800
X503 4129 2808 VDD VSS 4151 AND2X2TR $T=121400 25000 1 0 $X=121060 $Y=21000
X504 2800 2759 VDD VSS 2804 AND2X2TR $T=121800 82600 1 0 $X=121460 $Y=78600
X505 2801 2759 VDD VSS 2805 AND2X2TR $T=122200 89800 1 0 $X=121860 $Y=85800
X506 2802 4152 VDD VSS 4160 AND2X2TR $T=122200 97000 0 0 $X=121860 $Y=96720
X507 4141 2179 VDD VSS 4159 AND2X2TR $T=122600 10600 0 0 $X=122260 $Y=10320
X508 2364 2759 VDD VSS 4152 AND2X2TR $T=125000 89800 1 180 $X=122660 $Y=89520
X509 4170 2364 VDD VSS 4167 AND2X2TR $T=125800 53800 1 180 $X=123460 $Y=53520
X510 2816 2808 VDD VSS 4174 AND2X2TR $T=124200 25000 0 0 $X=123860 $Y=24720
X511 4166 2364 VDD VSS 4183 AND2X2TR $T=124200 46600 1 0 $X=123860 $Y=42600
X512 4163 4196 VDD VSS 2811 AND2X2TR $T=124600 118600 1 0 $X=124260 $Y=114600
X513 2806 4196 VDD VSS 4184 AND2X2TR $T=125400 111400 0 0 $X=125060 $Y=111120
X514 2809 2759 VDD VSS 4170 AND2X2TR $T=127800 53800 1 180 $X=125460 $Y=53520
X515 4174 2716 VDD VSS 4185 AND2X2TR $T=126600 25000 0 0 $X=126260 $Y=24720
X516 4171 2716 VDD VSS 2807 AND2X2TR $T=126600 32200 0 0 $X=126260 $Y=31920
X517 4186 2759 VDD VSS 4166 AND2X2TR $T=129400 46600 0 180 $X=127060 $Y=42600
X518 4178 4196 VDD VSS 4188 AND2X2TR $T=127800 125800 1 0 $X=127460 $Y=121800
X519 4175 2179 VDD VSS 4192 AND2X2TR $T=128600 17800 1 0 $X=128260 $Y=13800
X520 4176 2179 VDD VSS 4193 AND2X2TR $T=128600 25000 1 0 $X=128260 $Y=21000
X521 4185 2179 VDD VSS 2819 AND2X2TR $T=129000 25000 0 0 $X=128660 $Y=24720
X522 2807 2179 VDD VSS 4195 AND2X2TR $T=129400 32200 0 0 $X=129060 $Y=31920
X523 2832 2810 VDD VSS 2840 AND2X2TR $T=130200 82600 0 0 $X=129860 $Y=82320
X524 4190 2810 VDD VSS 2831 AND2X2TR $T=130200 104200 0 0 $X=129860 $Y=103920
X525 4188 2810 VDD VSS 4198 AND2X2TR $T=130200 125800 1 0 $X=129860 $Y=121800
X526 4194 4196 VDD VSS 4199 AND2X2TR $T=130600 68200 1 0 $X=130260 $Y=64200
X527 4199 2808 VDD VSS 2857 AND2X2TR $T=131000 61000 0 0 $X=130660 $Y=60720
X528 2826 2808 VDD VSS 2839 AND2X2TR $T=131000 75400 0 0 $X=130660 $Y=75120
X529 4197 2808 VDD VSS 2830 AND2X2TR $T=131400 61000 1 0 $X=131060 $Y=57000
X530 4198 2812 VDD VSS 2855 AND2X2TR $T=131400 125800 0 0 $X=131060 $Y=125520
X531 2831 2812 VDD VSS 2837 AND2X2TR $T=132600 104200 1 0 $X=132260 $Y=100200
X532 2840 2812 VDD VSS 2842 AND2X2TR $T=134200 82600 0 0 $X=133860 $Y=82320
X533 2857 2812 VDD VSS 4212 AND2X2TR $T=139400 61000 0 180 $X=137060 $Y=57000
X586 2210 VSS VDD 2644 CLKINVX2TR $T=87400 53800 0 0 $X=87060 $Y=53520
X587 2651 VSS VDD 2723 CLKINVX2TR $T=105400 125800 1 180 $X=103860 $Y=125520
X588 4013 VSS VDD 4022 CLKINVX2TR $T=105800 25000 0 0 $X=105460 $Y=24720
X589 2786 VSS VDD 4087 CLKINVX2TR $T=114600 89800 0 0 $X=114260 $Y=89520
X638 4184 2810 VSS VDD 2365 CLKAND2X2TR $T=128600 118600 0 180 $X=126260 $Y=114600
X639 2821 2810 VSS VDD 2835 CLKAND2X2TR $T=130200 118600 0 0 $X=129860 $Y=118320
X640 2526 2175 2179 2555 VDD VSS 3745 DFFRX1TR $T=46600 32200 0 0 $X=46260 $Y=31920
X641 3817 2175 2179 2591 VDD VSS 3832 DFFRX1TR $T=63800 25000 1 0 $X=63460 $Y=21000
X642 signature<15> 2202 2201 4444 VDD VSS 2875 DFFRX1TR $T=133800 118600 1 0 $X=133460 $Y=114600
X643 3811 VSS 2609 3806 VDD NAND2X1TR $T=68200 125800 1 180 $X=66260 $Y=125520
X644 2588 VSS 2601 2573 VDD NAND2X1TR $T=71800 125800 1 0 $X=71460 $Y=121800
X645 2622 VSS 3883 2617 VDD NAND2X1TR $T=80600 111400 1 180 $X=78660 $Y=111120
X646 3899 VSS 2642 3903 VDD NAND2X1TR $T=84200 17800 1 0 $X=83860 $Y=13800
X647 2627 VSS 2655 2663 VDD NAND2X1TR $T=85000 111400 1 0 $X=84660 $Y=107400
X648 2281 VSS 2712 3931 VDD NAND2X1TR $T=92200 125800 1 180 $X=90260 $Y=125520
X649 2647 VSS 2691 2664 VDD NAND2X1TR $T=92200 17800 0 0 $X=91860 $Y=17520
X650 2660 VSS 2695 3962 VDD NAND2X1TR $T=95000 17800 1 0 $X=94660 $Y=13800
X651 3957 VSS 2682 2667 VDD NAND2X1TR $T=95000 25000 1 0 $X=94660 $Y=21000
X652 2690 VSS 2676 2666 VDD NAND2X1TR $T=97800 118600 1 0 $X=97460 $Y=114600
X653 2691 VSS 2693 2695 VDD NAND2X1TR $T=98200 17800 1 0 $X=97860 $Y=13800
X654 2701 VSS 2710 2678 VDD NAND2X1TR $T=101000 97000 1 0 $X=100660 $Y=93000
X655 2318 VSS 4015 2323 VDD NAND2X1TR $T=104200 89800 0 180 $X=102260 $Y=85800
X656 2651 VSS 2722 2711 VDD NAND2X1TR $T=104600 125800 0 180 $X=102660 $Y=121800
X657 4036 VSS 2733 4022 VDD NAND2X1TR $T=107000 25000 0 180 $X=105060 $Y=21000
X658 2719 VSS 2785 2731 VDD NAND2X1TR $T=109000 39400 1 0 $X=108660 $Y=35400
X659 2740 VSS 4049 4065 VDD NAND2X1TR $T=112200 68200 0 180 $X=110260 $Y=64200
X660 4064 VSS 2754 4056 VDD NAND2X1TR $T=112200 75400 1 180 $X=110260 $Y=75120
X661 2745 VSS 2793 2735 VDD NAND2X1TR $T=113000 104200 0 180 $X=111060 $Y=100200
X662 4070 VSS 2761 2739 VDD NAND2X1TR $T=113400 25000 1 180 $X=111460 $Y=24720
X663 2742 VSS 2744 4065 VDD NAND2X1TR $T=113400 68200 1 180 $X=111460 $Y=67920
X664 2742 VSS 2748 2740 VDD NAND2X1TR $T=112200 68200 1 0 $X=111860 $Y=64200
X665 4075 VSS 2757 2726 VDD NAND2X1TR $T=114200 46600 1 180 $X=112260 $Y=46320
X666 2747 VSS 2751 2752 VDD NAND2X1TR $T=113000 53800 1 0 $X=112660 $Y=49800
X667 2768 VSS 2778 4090 VDD NAND2X1TR $T=117000 82600 0 180 $X=115060 $Y=78600
X668 2762 VSS 2789 2773 VDD NAND2X1TR $T=115400 97000 0 0 $X=115060 $Y=96720
X669 2766 VSS 2773 2735 VDD NAND2X1TR $T=116600 97000 1 0 $X=116260 $Y=93000
X670 4107 VSS 2783 2343 VDD NAND2X1TR $T=117400 46600 0 0 $X=117060 $Y=46320
X671 2785 VSS 2799 2787 VDD NAND2X1TR $T=118600 39400 1 0 $X=118260 $Y=35400
X672 2757 VSS 4132 2783 VDD NAND2X1TR $T=119400 46600 0 0 $X=119060 $Y=46320
X673 2751 VSS 4146 4139 VDD NAND2X1TR $T=121400 53800 1 0 $X=121060 $Y=49800
X674 2208 VDD 2203 2538 VSS NOR2X1TR $T=50600 82600 1 0 $X=50260 $Y=78600
X675 2181 VDD 2197 2145 VSS NOR2X1TR $T=58200 75400 1 180 $X=56260 $Y=75120
X676 2210 VDD 2197 2537 VSS NOR2X1TR $T=58200 89800 1 180 $X=56260 $Y=89520
X677 2203 VDD 2185 2561 VSS NOR2X1TR $T=59000 82600 0 0 $X=58660 $Y=82320
X678 2551 VDD 2560 3788 VSS NOR2X1TR $T=59400 68200 1 0 $X=59060 $Y=64200
X679 2210 VDD 2185 3776 VSS NOR2X1TR $T=62600 89800 1 180 $X=60660 $Y=89520
X680 2566 VDD 2567 2212 VSS NOR2X1TR $T=62200 125800 0 0 $X=61860 $Y=125520
X681 2144 VDD 2209 2554 VSS NOR2X1TR $T=65000 82600 1 180 $X=63060 $Y=82320
X682 2198 VDD 2209 3823 VSS NOR2X1TR $T=71400 82600 1 180 $X=69460 $Y=82320
X683 2198 VDD 2205 2182 VSS NOR2X1TR $T=71800 68200 1 180 $X=69860 $Y=67920
X684 2243 VDD 2197 2578 VSS NOR2X1TR $T=71800 75400 1 0 $X=71460 $Y=71400
X685 2588 VDD 2573 2590 VSS NOR2X1TR $T=71800 118600 0 0 $X=71460 $Y=118320
X686 2243 VDD 2205 2603 VSS NOR2X1TR $T=74200 32200 1 180 $X=72260 $Y=31920
X687 2197 VDD 2598 2597 VSS NOR2X1TR $T=72600 61000 1 0 $X=72260 $Y=57000
X688 2198 VDD 2185 3835 VSS NOR2X1TR $T=74200 104200 0 180 $X=72260 $Y=100200
X689 2210 VDD 2208 2614 VSS NOR2X1TR $T=75400 82600 1 0 $X=75060 $Y=78600
X690 2210 VDD 2248 2608 VSS NOR2X1TR $T=75400 82600 0 0 $X=75060 $Y=82320
X691 2144 VDD 2185 3850 VSS NOR2X1TR $T=77000 104200 0 180 $X=75060 $Y=100200
X692 2208 VDD 2181 2611 VSS NOR2X1TR $T=75800 75400 1 0 $X=75460 $Y=71400
X693 2622 VDD 2617 3862 VSS NOR2X1TR $T=76200 111400 0 0 $X=75860 $Y=111120
X694 2198 VDD 2197 2612 VSS NOR2X1TR $T=77000 104200 1 0 $X=76660 $Y=100200
X695 2208 VDD 2598 2618 VSS NOR2X1TR $T=77400 39400 1 0 $X=77060 $Y=35400
X696 2247 VDD 2244 2596 VSS NOR2X1TR $T=79400 32200 0 180 $X=77460 $Y=28200
X697 2181 VDD 2209 3873 VSS NOR2X1TR $T=77800 39400 0 0 $X=77460 $Y=39120
X698 2208 VDD 2244 2626 VSS NOR2X1TR $T=78600 46600 1 0 $X=78260 $Y=42600
X699 2144 VDD 2197 2622 VSS NOR2X1TR $T=78600 104200 1 0 $X=78260 $Y=100200
X700 2197 VDD 2244 3881 VSS NOR2X1TR $T=79400 82600 1 0 $X=79060 $Y=78600
X701 2243 VDD 2208 2621 VSS NOR2X1TR $T=81800 53800 0 180 $X=79860 $Y=49800
X702 2247 VDD 2598 3903 VSS NOR2X1TR $T=80600 17800 0 0 $X=80260 $Y=17520
X703 2598 VDD 2209 2631 VSS NOR2X1TR $T=81000 32200 1 0 $X=80660 $Y=28200
X704 2185 VDD 2598 2266 VSS NOR2X1TR $T=82600 53800 1 180 $X=80660 $Y=53520
X705 2248 VDD 2598 2273 VSS NOR2X1TR $T=81800 46600 1 0 $X=81460 $Y=42600
X706 2185 VDD 2244 3892 VSS NOR2X1TR $T=81800 82600 1 0 $X=81460 $Y=78600
X707 2243 VDD 2185 2275 VSS NOR2X1TR $T=82200 68200 0 0 $X=81860 $Y=67920
X708 2247 VDD 2181 2272 VSS NOR2X1TR $T=82600 39400 0 0 $X=82260 $Y=39120
X709 2243 VDD 2228 3899 VSS NOR2X1TR $T=85000 17800 1 180 $X=83060 $Y=17520
X710 2627 VDD 2663 3912 VSS NOR2X1TR $T=85000 104200 0 0 $X=84660 $Y=103920
X711 2243 VDD 2209 2635 VSS NOR2X1TR $T=86200 39400 1 0 $X=85860 $Y=35400
X712 2228 VDD 2598 2316 VSS NOR2X1TR $T=86600 17800 0 0 $X=86260 $Y=17520
X713 2205 VDD 2244 2641 VSS NOR2X1TR $T=87000 32200 1 0 $X=86660 $Y=28200
X714 2205 VDD 2598 2640 VSS NOR2X1TR $T=87400 25000 1 0 $X=87060 $Y=21000
X715 2244 VDD 2209 2643 VSS NOR2X1TR $T=87400 46600 1 0 $X=87060 $Y=42600
X716 2210 VDD 2228 3927 VSS NOR2X1TR $T=87800 46600 0 0 $X=87460 $Y=46320
X717 2228 VDD 2244 2647 VSS NOR2X1TR $T=88200 25000 0 0 $X=87860 $Y=24720
X718 2210 VDD 2209 3944 VSS NOR2X1TR $T=91000 68200 0 0 $X=90660 $Y=67920
X719 3957 VDD 2667 2679 VSS NOR2X1TR $T=94200 25000 0 0 $X=93860 $Y=24720
X720 2678 VDD 2701 2650 VSS NOR2X1TR $T=96600 104200 0 180 $X=94660 $Y=100200
X721 2323 VDD 2318 4019 VSS NOR2X1TR $T=102600 97000 1 0 $X=102260 $Y=93000
X722 4064 VDD 4056 4040 VSS NOR2X1TR $T=112200 82600 0 180 $X=110260 $Y=78600
X723 4075 VDD 2726 2775 VSS NOR2X1TR $T=114200 46600 0 0 $X=113860 $Y=46320
X724 2790 VDD 4084 4088 VSS NOR2X1TR $T=117000 104200 1 180 $X=115060 $Y=103920
X725 2775 VDD 2770 2767 VSS NOR2X1TR $T=118200 53800 0 180 $X=116260 $Y=49800
X726 2797 VDD 2793 2790 VSS NOR2X1TR $T=120600 104200 0 180 $X=118660 $Y=100200
X727 3823 VSS 2582 3818 VDD 2579 OAI21X1TR $T=71400 89800 1 180 $X=69060 $Y=89520
X728 2635 VSS 2646 2641 VDD 3948 OAI21X1TR $T=91800 32200 0 0 $X=91460 $Y=31920
X729 2680 VSS 2677 2658 VDD 2674 OAI21X1TR $T=97400 89800 0 180 $X=95060 $Y=85800
X730 2721 VSS 2665 2697 VDD 2717 OAI21X1TR $T=106200 104200 1 180 $X=103860 $Y=103920
X731 4013 VSS 2736 4036 VDD 2760 OAI21X1TR $T=107400 25000 1 0 $X=107060 $Y=21000
X732 2330 VSS 2762 2721 VDD 4084 OAI21X1TR $T=113400 104200 1 0 $X=113060 $Y=100200
X733 2757 VSS 2770 2751 VDD 2765 OAI21X1TR $T=114600 53800 1 0 $X=114260 $Y=49800
X734 2649 2695 VDD 2698 VSS 3992 AOI21X1TR $T=99000 17800 0 0 $X=98660 $Y=17520
X735 2666 2656 VDD 3981 VSS 2311 AOI21X1TR $T=102600 111400 1 180 $X=100260 $Y=111120
X736 2661 4039 VDD 2656 VSS 3985 AOI21X1TR $T=102600 118600 1 180 $X=100260 $Y=118320
X737 2711 4039 VDD 2723 VSS 2732 AOI21X1TR $T=107000 125800 0 0 $X=106660 $Y=125520
X738 2324 2728 VDD 2717 VSS 4037 AOI21X1TR $T=109400 104200 1 180 $X=107060 $Y=103920
X739 2739 2760 VDD 2741 VSS 2756 AOI21X1TR $T=113000 32200 1 0 $X=112660 $Y=28200
X740 2343 2767 VDD 2765 VSS 4073 AOI21X1TR $T=115800 53800 1 180 $X=113460 $Y=53520
X741 2593 2263 VSS VDD 2278 AND2X1TR $T=83400 82600 1 0 $X=83060 $Y=78600
X742 2316 2716 VSS VDD 2743 AND2X1TR $T=111000 17800 0 0 $X=110660 $Y=17520
X743 2812 2716 VSS VDD BUFX3TR $T=129800 39400 0 180 $X=127460 $Y=35400
X744 2201 2179 VSS VDD BUFX4TR $T=71400 39400 1 0 $X=71060 $Y=35400
X745 2442 VSS 2055 VDD CLKINVX16TR $T=16200 17800 0 180 $X=11060 $Y=13800
X746 2172 VSS 2175 VDD CLKINVX16TR $T=59000 68200 0 0 $X=58660 $Y=67920
X772 2175 3617 VDD VSS 2203 DFFHQX8TR $T=37000 68200 0 0 $X=36660 $Y=67920
X773 2202 2258 VDD VSS 2709 DFFHQX8TR $T=91400 89800 0 0 $X=91060 $Y=89520
X774 2202 4098 VDD VSS 4178 DFFHQX8TR $T=114600 125800 1 0 $X=114260 $Y=121800
X775 2175 2143 2198 VSS VDD DFFHQX4TR $T=37000 75400 1 0 $X=36660 $Y=71400
X776 2175 2521 2210 VSS VDD DFFHQX4TR $T=37400 53800 0 0 $X=37060 $Y=53520
X777 2175 3668 2208 VSS VDD DFFHQX4TR $T=45000 39400 0 0 $X=44660 $Y=39120
X778 2175 3689 2185 VSS VDD DFFHQX4TR $T=45800 61000 1 0 $X=45460 $Y=57000
X779 2175 2547 2180 VSS VDD DFFHQX4TR $T=58200 53800 0 180 $X=46260 $Y=49800
X780 2175 3696 2205 VSS VDD DFFHQX4TR $T=47000 25000 1 0 $X=46660 $Y=21000
X781 2175 2551 2144 VSS VDD DFFHQX4TR $T=59400 68200 0 180 $X=47460 $Y=64200
X782 2175 2555 2209 VSS VDD DFFHQX4TR $T=56200 32200 0 0 $X=55860 $Y=31920
X783 2175 2559 2181 VSS VDD DFFHQX4TR $T=58200 46600 0 0 $X=57860 $Y=46320
X784 2175 2560 2228 VSS VDD DFFHQX4TR $T=58200 61000 1 0 $X=57860 $Y=57000
X785 2175 2196 2247 VSS VDD DFFHQX4TR $T=63400 32200 1 0 $X=63060 $Y=28200
X786 2175 3801 2243 VSS VDD DFFHQX4TR $T=63800 17800 0 0 $X=63460 $Y=17520
X787 2305 2694 2742 VSS VDD DFFHQX4TR $T=97400 68200 1 0 $X=97060 $Y=64200
X788 2305 2754 2768 VSS VDD DFFHQX4TR $T=112200 75400 0 0 $X=111860 $Y=75120
X789 2305 2812 2808 VSS VDD DFFHQX4TR $T=134600 75400 0 180 $X=122660 $Y=71400
X790 2553 2175 2201 VSS 2142 VDD 2521 DFFSX2TR $T=46600 53800 0 180 $X=37860 $Y=49800
X791 2142 2175 2201 VSS 2522 VDD 3617 DFFSX2TR $T=47000 61000 1 180 $X=38260 $Y=60720
X792 2522 2175 2201 VSS 2527 VDD 2143 DFFSX2TR $T=38600 68200 1 0 $X=38260 $Y=64200
X793 3745 2175 2201 VSS 3686 VDD 3668 DFFSX2TR $T=55000 39400 0 180 $X=46260 $Y=35400
X794 2547 2175 2201 VSS 2184 VDD 3689 DFFSX2TR $T=55400 46600 1 180 $X=46660 $Y=46320
X795 3755 2175 2179 VSS 3698 VDD 3696 DFFSX2TR $T=57000 25000 1 180 $X=48260 $Y=24720
X796 2527 2175 2201 VSS 2541 VDD 2551 DFFSX2TR $T=52200 61000 0 0 $X=51860 $Y=60720
X797 2558 2175 2179 VSS 3755 VDD 2196 DFFSX2TR $T=63000 32200 0 180 $X=54260 $Y=28200
X798 2541 2175 2201 VSS 2558 VDD 2560 DFFSX2TR $T=54600 53800 0 0 $X=54260 $Y=53520
X799 3808 2175 2201 VSS 2553 VDD 2559 DFFSX2TR $T=65000 46600 0 180 $X=56260 $Y=42600
X800 2184 2175 2201 VSS 2206 VDD 3775 DFFSX2TR $T=69400 39400 1 180 $X=60660 $Y=39120
X801 3800 2175 2179 VSS 2583 VDD 4445 DFFSX2TR $T=64200 25000 0 0 $X=63860 $Y=24720
X802 3832 2175 2179 VSS 3800 VDD 3801 DFFSX2TR $T=73000 17800 0 180 $X=64260 $Y=13800
X803 4191 2202 2201 VSS signature<15> VDD 4446 DFFSX2TR $T=130600 133000 1 0 $X=130260 $Y=129000
X804 4203 2305 2179 VSS signature<0> VDD 4447 DFFSX2TR $T=131400 10600 0 0 $X=131060 $Y=10320
X805 2866 2305 2179 VSS signature<1> VDD 4448 DFFSX2TR $T=139800 17800 0 180 $X=131060 $Y=13800
X806 2836 2305 2179 VSS signature<3> VDD 4449 DFFSX2TR $T=134200 32200 1 0 $X=133860 $Y=28200
X807 2854 2202 2861 VSS signature<11> VDD 4450 DFFSX2TR $T=134200 104200 0 0 $X=133860 $Y=103920
X808 2846 2202 2861 VSS 4221 VDD 4451 DFFSX2TR $T=134200 111400 1 0 $X=133860 $Y=107400
X809 2871 2202 2201 VSS signature<13> VDD 4452 DFFSX2TR $T=142600 125800 0 180 $X=133860 $Y=121800
X810 2872 2202 2201 VSS signature<14> VDD 4453 DFFSX2TR $T=142600 133000 1 180 $X=133860 $Y=132720
X811 4205 2305 2179 VSS signature<2> VDD 4454 DFFSX2TR $T=134600 17800 0 0 $X=134260 $Y=17520
X812 2860 2305 2861 VSS signature<4> VDD 4455 DFFSX2TR $T=134600 39400 1 0 $X=134260 $Y=35400
X813 2838 2305 2861 VSS signature<5> VDD 4456 DFFSX2TR $T=134600 46600 0 0 $X=134260 $Y=46320
X814 2845 2305 2861 VSS signature<6> VDD 4457 DFFSX2TR $T=134600 53800 0 0 $X=134260 $Y=53520
X815 4206 2305 2861 VSS signature<7> VDD 4458 DFFSX2TR $T=134600 68200 0 0 $X=134260 $Y=67920
X816 2853 2305 2861 VSS signature<8> VDD 4459 DFFSX2TR $T=134600 82600 1 0 $X=134260 $Y=78600
X817 2859 2202 2861 VSS signature<9> VDD 4460 DFFSX2TR $T=134600 89800 1 0 $X=134260 $Y=85800
X836 2548 2536 2145 2146 VSS VDD 2525 ADDFHX2TR $T=57800 89800 0 180 $X=42660 $Y=85800
X837 2534 2146 2552 2556 VSS VDD 2557 ADDFHX2TR $T=44600 104200 0 0 $X=44260 $Y=103920
X838 2546 2211 2199 3807 VSS VDD 2280 ADDFHX2TR $T=53800 104200 1 0 $X=53460 $Y=100200
X839 2538 2569 2183 3810 VSS VDD 3818 ADDFHX2TR $T=54600 82600 1 0 $X=54260 $Y=78600
X840 2570 2584 2597 2257 VSS VDD 2256 ADDFHX2TR $T=62600 61000 0 0 $X=62260 $Y=60720
X841 2612 3850 2615 2617 VSS VDD 2624 ADDFHX2TR $T=66200 104200 0 0 $X=65860 $Y=103920
X842 3828 3873 2626 2261 VSS VDD 2683 ADDFHX2TR $T=71400 46600 0 0 $X=71060 $Y=46320
X843 2596 2625 2631 2259 VSS VDD 2667 ADDFHX2TR $T=73000 25000 0 0 $X=72660 $Y=24720
X844 2616 2276 2277 2267 VSS VDD 2638 ADDFHX2TR $T=76600 75400 0 0 $X=76260 $Y=75120
X845 2605 3930 3923 3932 VSS VDD 2652 ADDFHX2TR $T=77000 97000 1 0 $X=76660 $Y=93000
X846 2611 3908 2275 2276 VSS VDD 2692 ADDFHX2TR $T=77800 75400 1 0 $X=77460 $Y=71400
X847 2623 3932 2280 2663 VSS VDD 2701 ADDFHX2TR $T=80200 104200 1 0 $X=79860 $Y=100200
X848 2621 3938 2255 3964 VSS VDD 3971 ADDFHX2TR $T=82200 53800 1 0 $X=81860 $Y=49800
X849 2706 2256 2261 2659 VSS VDD 2694 ADDFHX2TR $T=100600 61000 1 180 $X=85460 $Y=60720
X850 2274 2689 2707 2706 VSS VDD 2705 ADDFHX2TR $T=89400 61000 1 0 $X=89060 $Y=57000
X851 2696 4014 2703 4075 VSS VDD 2731 ADDFHX2TR $T=99400 39400 0 0 $X=99060 $Y=39120
X887 3680 2561 2537 2545 VSS VDD 2552 ADDFX2TR $T=45800 89800 0 0 $X=45460 $Y=89520
X888 2554 3776 3810 2572 VSS VDD 2571 ADDFX2TR $T=57800 97000 1 0 $X=57460 $Y=93000
X889 3892 2251 2278 2279 VSS VDD 2636 ADDFX2TR $T=83000 82600 0 0 $X=82660 $Y=82320
X890 2273 2643 2672 2704 VSS VDD 2654 ADDFX2TR $T=89800 46600 1 0 $X=89460 $Y=42600
X891 3980 2709 2652 2678 VSS VDD 2318 ADDFX2TR $T=101000 97000 0 180 $X=91460 $Y=93000
X892 2714 2317 2720 2323 VSS VDD 4056 ADDFX2TR $T=101400 82600 1 0 $X=101060 $Y=78600
X893 2208 2144 3680 VSS VDD NOR2X2TR $T=48600 82600 0 180 $X=46260 $Y=78600
X894 2208 2198 2536 VSS VDD NOR2X2TR $T=49800 82600 0 0 $X=49460 $Y=82320
X895 2205 2144 2569 VSS VDD NOR2X2TR $T=63800 68200 0 0 $X=63460 $Y=67920
X896 2248 2203 2548 VSS VDD NOR2X2TR $T=66200 82600 0 0 $X=65860 $Y=82320
X897 2248 2181 3803 VSS VDD NOR2X2TR $T=69000 75400 0 180 $X=66660 $Y=71400
X898 2205 2181 2585 VSS VDD NOR2X2TR $T=69800 53800 1 0 $X=69460 $Y=49800
X899 2205 2203 3847 VSS VDD NOR2X2TR $T=73400 68200 0 0 $X=73060 $Y=67920
X900 2228 2181 2606 VSS VDD NOR2X2TR $T=73800 39400 0 0 $X=73460 $Y=39120
X901 2228 2203 3848 VSS VDD NOR2X2TR $T=73800 53800 0 0 $X=73460 $Y=53520
X902 2247 2144 3876 VSS VDD NOR2X2TR $T=78200 68200 0 0 $X=77860 $Y=67920
X903 2248 2243 2274 VSS VDD NOR2X2TR $T=81000 61000 1 0 $X=80660 $Y=57000
X904 2228 2198 2282 VSS VDD NOR2X2TR $T=85400 68200 0 180 $X=83060 $Y=64200
X905 2198 2247 3908 VSS VDD NOR2X2TR $T=83800 68200 0 0 $X=83460 $Y=67920
X906 2243 2247 2634 VSS VDD NOR2X2TR $T=84600 25000 1 0 $X=84260 $Y=21000
X907 2205 2210 2673 VSS VDD NOR2X2TR $T=87800 68200 1 0 $X=87460 $Y=64200
X908 2212 2633 2661 VSS VDD NOR2X2TR $T=90600 118600 0 0 $X=90260 $Y=118320
X909 2330 2665 2324 VSS VDD NOR2X2TR $T=105800 104200 0 180 $X=103460 $Y=100200
X910 2731 2719 2725 VSS VDD NOR2X2TR $T=105400 39400 1 0 $X=105060 $Y=35400
X911 2752 2747 2770 VSS VDD NOR2X2TR $T=112200 53800 1 180 $X=109860 $Y=53520
X912 4076 2786 2735 VSS VDD NOR2X2TR $T=113400 97000 1 0 $X=113060 $Y=93000
X913 3686 2175 2201 VSS 2547 VDD DFFSX1TR $T=47000 46600 1 0 $X=46660 $Y=42600
X914 2851 2202 2861 VSS signature<10> VDD DFFSX1TR $T=134600 97000 0 0 $X=134260 $Y=96720
X915 2557 2202 VSS VDD 2528 DFFHQX1TR $T=55400 111400 0 180 $X=47060 $Y=107400
X916 2525 2202 VSS VDD 2546 DFFHQX1TR $T=48200 97000 0 0 $X=47860 $Y=96720
X917 3811 2202 VSS VDD 2566 DFFHQX1TR $T=67400 125800 0 180 $X=59060 $Y=121800
X918 3806 2202 VSS VDD 2567 DFFHQX1TR $T=67800 133000 0 180 $X=59460 $Y=129000
X919 3788 2175 VSS VDD 2580 DFFHQX1TR $T=62200 68200 1 0 $X=61860 $Y=64200
X920 2279 2202 VSS VDD 2605 DFFHQX1TR $T=82600 89800 1 180 $X=74260 $Y=89520
X921 2609 2202 VSS VDD 2651 DFFHQX1TR $T=77400 125800 1 0 $X=77060 $Y=121800
X922 2629 2202 VSS VDD 3930 DFFHQX1TR $T=82600 97000 0 0 $X=82260 $Y=96720
X923 2636 2202 VSS VDD 2658 DFFHQX1TR $T=85400 89800 1 0 $X=85060 $Y=85800
X924 3912 2202 VSS VDD 2665 DFFHQX1TR $T=86600 104200 0 0 $X=86260 $Y=103920
X925 2654 2305 VSS VDD 2703 DFFHQX1TR $T=91400 39400 0 0 $X=91060 $Y=39120
X926 2655 2202 VSS VDD 2697 DFFHQX1TR $T=91800 111400 1 0 $X=91460 $Y=107400
X927 2257 2202 VSS VDD 2677 DFFHQX1TR $T=93400 82600 1 0 $X=93060 $Y=78600
X928 2679 2305 VSS VDD 4013 DFFHQX1TR $T=96600 25000 0 0 $X=96260 $Y=24720
X929 2271 2305 VSS VDD 2718 DFFHQX1TR $T=96600 32200 1 0 $X=96260 $Y=28200
X930 2683 2305 VSS VDD 4012 DFFHQX1TR $T=97000 53800 1 0 $X=96660 $Y=49800
X931 2682 2305 VSS VDD 4036 DFFHQX1TR $T=97400 25000 1 0 $X=97060 $Y=21000
X932 2710 2202 VSS VDD 2721 DFFHQX1TR $T=99400 97000 0 0 $X=99060 $Y=96720
X933 2704 2305 VSS VDD 2699 DFFHQX1TR $T=108600 46600 0 180 $X=100260 $Y=42600
X934 2708 2305 VSS VDD 2680 DFFHQX1TR $T=101400 75400 0 0 $X=101060 $Y=75120
X935 2700 2305 VSS VDD 2734 DFFHQX1TR $T=101800 32200 0 0 $X=101460 $Y=31920
X936 3992 2305 VSS VDD 2736 DFFHQX1TR $T=102200 17800 0 0 $X=101860 $Y=17520
X937 4002 2305 VSS VDD 2740 DFFHQX1TR $T=102200 53800 0 0 $X=101860 $Y=53520
X938 4017 2305 VSS VDD 4065 DFFHQX1TR $T=104600 75400 1 0 $X=104260 $Y=71400
X939 4006 2305 VSS VDD 2727 DFFHQX1TR $T=105000 53800 1 0 $X=104660 $Y=49800
X940 4015 2202 VSS VDD 2749 DFFHQX1TR $T=105000 89800 1 0 $X=104660 $Y=85800
X941 4073 2305 VSS VDD 2797 DFFHQX1TR $T=112600 75400 1 0 $X=112260 $Y=71400
X942 2774 2202 VSS VDD 4168 DFFHQX1TR $T=117000 118600 0 0 $X=116660 $Y=118320
X943 2364 2305 VSS VDD 4196 DFFHQX1TR $T=123400 68200 0 0 $X=123060 $Y=67920
X944 2184 3698 2526 VDD VSS XOR2X1TR $T=48200 32200 1 0 $X=47860 $Y=28200
X945 2206 2583 3808 VDD VSS XOR2X1TR $T=69400 39400 0 180 $X=65860 $Y=35400
X946 2184 2206 3817 VDD VSS XOR2X1TR $T=71000 32200 1 180 $X=67460 $Y=31920
X947 3818 3823 2587 VDD VSS XOR2X1TR $T=69400 89800 1 0 $X=69060 $Y=85800
X948 2587 2582 2258 VDD VSS XOR2X1TR $T=71400 89800 0 0 $X=71060 $Y=89520
X949 2618 3880 3900 VDD VSS XOR2X1TR $T=79400 32200 0 0 $X=79060 $Y=31920
X950 3900 2259 2271 VDD VSS XOR2X1TR $T=83800 32200 1 0 $X=83460 $Y=28200
X951 2641 2635 2653 VDD VSS XOR2X1TR $T=90200 32200 1 0 $X=89860 $Y=28200
X952 2646 2653 2700 VDD VSS XOR2X1TR $T=93400 32200 1 0 $X=93060 $Y=28200
X953 2680 2658 2668 VDD VSS XOR2X1TR $T=97000 82600 1 180 $X=93460 $Y=82320
X954 2668 2677 2720 VDD VSS XOR2X1TR $T=99000 82600 0 0 $X=98660 $Y=82320
X955 2722 4027 2730 VDD VSS XOR2X1TR $T=107000 118600 0 0 $X=106660 $Y=118320
X956 2732 2712 2750 VDD VSS XOR2X1TR $T=109400 125800 0 0 $X=109060 $Y=125520
X957 2742 4061 2752 VDD VSS XOR2X1TR $T=113000 61000 0 180 $X=109460 $Y=57000
X958 2740 4065 4061 VDD VSS XOR2X1TR $T=109800 61000 0 0 $X=109460 $Y=60720
X959 2733 2736 2798 VDD VSS XOR2X1TR $T=110200 25000 1 0 $X=109860 $Y=21000
X960 4088 2758 2753 VDD VSS XOR2X1TR $T=115800 111400 0 180 $X=112260 $Y=107400
X961 4118 2788 2801 VDD VSS XOR2X1TR $T=118200 89800 1 0 $X=117860 $Y=85800
X962 4119 2789 2802 VDD VSS XOR2X1TR $T=118200 97000 0 0 $X=117860 $Y=96720
X963 4155 4157 4140 VDD VSS XOR2X1TR $T=124200 61000 1 180 $X=120660 $Y=60720
X964 2756 2799 4145 VDD VSS XOR2X1TR $T=121400 39400 1 0 $X=121060 $Y=35400
X965 signature<14> 2822 4191 VDD VSS XOR2X1TR $T=131800 133000 1 180 $X=128260 $Y=132720
X966 2856 signature<15> 2836 VDD VSS XOR2X1TR $T=134200 25000 1 180 $X=130660 $Y=24720
X967 signature<15> 2813 4203 VDD VSS XOR2X1TR $T=131400 17800 0 0 $X=131060 $Y=17520
X968 signature<1> 2823 4205 VDD VSS XOR2X1TR $T=133000 10600 1 0 $X=132660 $Y=6600
X969 signature<6> 4208 4206 VDD VSS XOR2X1TR $T=137400 61000 1 180 $X=133860 $Y=60720
X970 signature<5> 4212 2845 VDD VSS XOR2X1TR $T=138600 53800 0 180 $X=135060 $Y=49800
X971 signature<11> 2849 2846 VDD VSS XOR2X1TR $T=138600 111400 1 180 $X=135060 $Y=111120
X972 signature<9> 2847 2851 VDD VSS XOR2X1TR $T=136200 97000 1 0 $X=135860 $Y=93000
X973 signature<9> 2837 2854 VDD VSS XOR2X1TR $T=136600 104200 1 0 $X=136260 $Y=100200
X974 signature<7> 2858 2853 VDD VSS XOR2X1TR $T=140200 75400 1 180 $X=136660 $Y=75120
X975 signature<2> 4218 2856 VDD VSS XOR2X1TR $T=140600 25000 0 180 $X=137060 $Y=21000
X976 signature<4> 2843 2838 VDD VSS XOR2X1TR $T=140600 46600 0 180 $X=137060 $Y=42600
X977 signature<8> 2842 2859 VDD VSS XOR2X1TR $T=140600 82600 1 180 $X=137060 $Y=82320
X978 signature<13> 2855 2872 VDD VSS XOR2X1TR $T=137400 125800 0 0 $X=137060 $Y=125520
X979 signature<12> 2841 2871 VDD VSS XOR2X1TR $T=137800 118600 0 0 $X=137460 $Y=118320
X980 signature<3> 2862 2860 VDD VSS XOR2X1TR $T=141400 32200 1 180 $X=137860 $Y=31920
X981 2875 4221 signature<12> VDD VSS XOR2X1TR $T=141800 111400 1 180 $X=138260 $Y=111120
X982 signature<0> 2369 2865 VDD VSS XOR2X1TR $T=139800 10600 0 0 $X=139460 $Y=10320
X983 2865 signature<15> 2866 VDD VSS XOR2X1TR $T=139800 17800 1 0 $X=139460 $Y=13800
X984 2545 2202 VSS VDD 2565 DFFQX1TR $T=55800 111400 1 180 $X=48660 $Y=111120
X985 2556 2202 VSS VDD 2200 DFFQX1TR $T=56200 118600 0 180 $X=49060 $Y=114600
X986 2571 2202 VSS VDD 2199 DFFQX1TR $T=63400 97000 1 180 $X=56260 $Y=96720
X987 2572 2202 VSS VDD 2564 DFFQX1TR $T=66200 104200 1 180 $X=59060 $Y=103920
X988 2613 2202 VSS VDD 2563 DFFQX1TR $T=67400 118600 0 180 $X=60260 $Y=114600
X989 2624 2202 VSS VDD 2588 DFFQX1TR $T=76200 118600 0 180 $X=69060 $Y=114600
X990 3833 2202 VSS VDD 2623 DFFQX1TR $T=72600 97000 0 0 $X=72260 $Y=96720
X991 2601 2202 VSS VDD 2281 DFFQX1TR $T=77000 125800 0 0 $X=76660 $Y=125520
X992 3862 2202 VSS VDD 2632 DFFQX1TR $T=77400 118600 1 0 $X=77060 $Y=114600
X993 2590 2202 VSS VDD 2633 DFFQX1TR $T=77400 118600 0 0 $X=77060 $Y=118320
X994 3883 2202 VSS VDD 3921 DFFQX1TR $T=81000 111400 0 0 $X=80660 $Y=111120
X995 2267 2202 VSS VDD 3923 DFFQX1TR $T=82600 89800 0 0 $X=82260 $Y=89520
X996 2638 2202 VSS VDD 2317 DFFQX1TR $T=85400 82600 1 0 $X=85060 $Y=78600
X997 3918 2202 VSS VDD 2666 DFFQX1TR $T=88200 118600 1 0 $X=87860 $Y=114600
X998 3921 2202 VSS VDD 2690 DFFQX1TR $T=88600 111400 0 0 $X=88260 $Y=111120
X999 2637 2305 VSS VDD 2719 DFFQX1TR $T=95000 32200 0 0 $X=94660 $Y=31920
X1000 4009 2305 VSS VDD 4055 DFFQX1TR $T=104200 10600 0 0 $X=103860 $Y=10320
X1001 4034 2305 VSS VDD 4079 DFFQX1TR $T=107800 17800 1 0 $X=107460 $Y=13800
X1002 4055 2305 VSS VDD 4113 DFFQX1TR $T=111000 10600 0 0 $X=110660 $Y=10320
X1003 2743 2305 VSS VDD 2795 DFFQX1TR $T=114200 17800 0 0 $X=113860 $Y=17520
X1004 2795 2305 VSS VDD 4129 DFFQX1TR $T=114200 25000 1 0 $X=113860 $Y=21000
X1005 4079 2305 VSS VDD 4137 DFFQX1TR $T=114600 17800 1 0 $X=114260 $Y=13800
X1006 2769 2305 VSS VDD 4162 DFFQX1TR $T=116600 32200 1 0 $X=116260 $Y=28200
X1007 4104 2305 VSS VDD 4155 DFFQX1TR $T=117000 53800 0 0 $X=116660 $Y=53520
X1008 2777 2305 VSS VDD 4157 DFFQX1TR $T=117800 61000 1 0 $X=117460 $Y=57000
X1009 2763 2202 VSS VDD 2806 DFFQX1TR $T=117800 111400 0 0 $X=117460 $Y=111120
X1010 2776 2202 VSS VDD 4163 DFFQX1TR $T=117800 118600 1 0 $X=117460 $Y=114600
X1011 2794 2202 VSS VDD 4179 DFFQX1TR $T=120200 111400 1 0 $X=119860 $Y=107400
X1012 4132 2305 VSS VDD 2372 DFFQX1TR $T=121000 46600 0 0 $X=120660 $Y=46320
X1013 4145 2305 VSS VDD 4186 DFFQX1TR $T=121800 39400 0 0 $X=121460 $Y=39120
X1014 4146 2305 VSS VDD 4187 DFFQX1TR $T=123000 53800 1 0 $X=122660 $Y=49800
X1015 4154 2305 VSS VDD 2816 DFFQX1TR $T=123400 32200 1 0 $X=123060 $Y=28200
X1016 4147 2305 VSS VDD 4194 DFFQX1TR $T=123800 68200 1 0 $X=123460 $Y=64200
X1017 4159 2305 VSS VDD 2823 DFFQX1TR $T=124200 10600 1 0 $X=123860 $Y=6600
X1018 2812 2305 VSS VDD 2364 DFFQX1TR $T=131000 75400 1 180 $X=123860 $Y=75120
X1019 4160 2202 VSS VDD 2820 DFFQX1TR $T=124200 97000 0 0 $X=123860 $Y=96720
X1020 4192 2305 VSS VDD 2369 DFFQX1TR $T=131400 10600 1 180 $X=124260 $Y=10320
X1021 4193 2305 VSS VDD 2813 DFFQX1TR $T=131400 17800 1 180 $X=124260 $Y=17520
X1022 4167 2305 VSS VDD 4197 DFFQX1TR $T=124600 61000 1 0 $X=124260 $Y=57000
X1023 4181 2305 VSS VDD 2826 DFFQX1TR $T=127400 82600 1 0 $X=127060 $Y=78600
X1024 4182 2202 VSS VDD 2832 DFFQX1TR $T=127400 89800 1 0 $X=127060 $Y=85800
X1025 4183 2305 VSS VDD 2833 DFFQX1TR $T=127800 46600 0 0 $X=127460 $Y=46320
X1026 4195 2305 VSS VDD 2862 DFFQX1TR $T=131400 32200 0 0 $X=131060 $Y=31920
X1027 2819 2305 VSS VDD 4218 DFFQX1TR $T=134200 25000 0 0 $X=133860 $Y=24720
X1028 2180 2198 VDD 2534 VSS NOR2BX1TR $T=52200 104200 0 180 $X=49860 $Y=100200
X1029 2593 2197 VDD 2619 VSS NOR2BX1TR $T=81800 97000 1 180 $X=79460 $Y=96720
X1030 2820 2824 VDD 2847 VSS NOR2BX1TR $T=129800 97000 1 0 $X=129460 $Y=93000
X1031 2563 2565 2200 2573 VSS VDD 3811 CMPR32X2TR $T=58600 118600 0 0 $X=58260 $Y=118320
X1032 2528 2564 3807 3806 VSS VDD 2627 CMPR32X2TR $T=59000 111400 1 0 $X=58660 $Y=107400
X1033 3944 2675 2692 2708 VSS VDD 4017 CMPR32X2TR $T=92600 75400 0 0 $X=92260 $Y=75120
X1034 2185 2181 VSS VDD 2562 OR2X2TR $T=59000 75400 1 0 $X=58660 $Y=71400
X1035 3903 3899 VSS VDD 2630 OR2X2TR $T=82200 17800 1 0 $X=81860 $Y=13800
X1036 2718 2734 VSS VDD 2739 OR2X2TR $T=109800 32200 1 0 $X=109460 $Y=28200
X1037 2725 2756 VSS VDD 4082 OR2X2TR $T=112600 39400 1 0 $X=112260 $Y=35400
X1038 2562 VSS VDD 2183 INVX2TR $T=59400 75400 0 0 $X=59060 $Y=75120
X1039 2203 VSS VDD 2593 INVX2TR $T=74200 82600 0 180 $X=72660 $Y=78600
X1040 3880 VSS VDD 3898 INVX2TR $T=80600 39400 1 0 $X=80260 $Y=35400
X1041 2247 VSS VDD 2648 INVX2TR $T=84200 53800 0 0 $X=83860 $Y=53520
X1042 2632 VSS VDD 3918 INVX2TR $T=85800 118600 1 0 $X=85460 $Y=114600
X1043 2633 VSS VDD 3931 INVX2TR $T=89400 125800 0 0 $X=89060 $Y=125520
X1044 2642 VSS VDD 2649 INVX2TR $T=89800 17800 1 0 $X=89460 $Y=13800
X1045 2209 VSS VDD 2263 INVX2TR $T=92600 75400 1 180 $X=91060 $Y=75120
X1046 2647 VSS VDD 2660 INVX2TR $T=92600 17800 1 0 $X=92260 $Y=13800
X1047 2664 VSS VDD 3962 INVX2TR $T=94600 17800 0 0 $X=94260 $Y=17520
X1048 2212 VSS VDD 2711 INVX2TR $T=96600 125800 0 0 $X=96260 $Y=125520
X1049 4039 VSS VDD 4027 INVX2TR $T=105800 118600 0 0 $X=105460 $Y=118320
X1050 4045 VSS VDD 4032 INVX2TR $T=106600 104200 1 0 $X=106260 $Y=100200
X1051 2741 VSS VDD 4070 INVX2TR $T=111800 32200 1 0 $X=111460 $Y=28200
X1052 2330 VSS VDD 2745 INVX2TR $T=111800 97000 0 0 $X=111460 $Y=96720
X1053 2728 VSS VDD 2762 INVX2TR $T=113400 104200 0 0 $X=113060 $Y=103920
X1054 4076 VSS VDD 4090 INVX2TR $T=113800 82600 0 0 $X=113460 $Y=82320
X1055 2725 VSS VDD 2787 INVX2TR $T=116200 39400 1 0 $X=115860 $Y=35400
X1056 2775 VSS VDD 4107 INVX2TR $T=116200 46600 0 0 $X=115860 $Y=46320
X1057 2768 VSS VDD 4103 INVX2TR $T=119000 82600 1 180 $X=117460 $Y=82320
X1058 2797 VSS VDD 2766 INVX2TR $T=119400 89800 1 180 $X=117860 $Y=89520
X1059 2770 VSS VDD 4139 INVX2TR $T=120200 53800 1 0 $X=119860 $Y=49800
X1060 2810 VSS VDD 4200 INVX2TR $T=131400 97000 0 0 $X=131060 $Y=96720
X1061 3775 2175 VDD VSS 2197 DFFHQX2TR $T=59800 53800 1 0 $X=59460 $Y=49800
X1062 2216 2202 VDD VSS 2211 DFFHQX2TR $T=63800 97000 0 0 $X=63460 $Y=96720
X1063 3808 2175 VDD VSS 2592 DFFHQX2TR $T=65000 46600 1 0 $X=64660 $Y=42600
X1064 2591 2175 VDD VSS 2598 DFFHQX2TR $T=73000 25000 1 0 $X=72660 $Y=21000
X1065 3971 2305 VDD VSS 2696 DFFHQX2TR $T=98200 46600 1 180 $X=89060 $Y=46320
X1066 2650 2202 VDD VSS 2330 DFFHQX2TR $T=90600 97000 0 0 $X=90260 $Y=96720
X1067 2659 2305 VDD VSS 2714 DFFHQX2TR $T=95800 75400 1 0 $X=95460 $Y=71400
X1068 2662 2305 VDD VSS 4014 DFFHQX2TR $T=96200 39400 1 0 $X=95860 $Y=35400
X1069 4019 2202 VDD VSS 2786 DFFHQX2TR $T=104600 89800 0 0 $X=104260 $Y=89520
X1070 4040 2202 VDD VSS 4076 DFFHQX2TR $T=105000 82600 0 0 $X=104660 $Y=82320
X1071 2182 3803 2578 2582 VSS VDD 2277 ADDFHX1TR $T=61800 75400 0 0 $X=61460 $Y=75120
X1072 2581 3835 2619 2615 VSS VDD 2613 ADDFHX1TR $T=68600 111400 1 0 $X=68260 $Y=107400
X1073 2266 3964 2705 4002 VSS VDD 4006 ADDFHX1TR $T=92200 53800 0 0 $X=91860 $Y=53520
X1074 2699 4012 2727 2747 VSS VDD 2726 ADDFHX1TR $T=98200 46600 0 0 $X=97860 $Y=46320
X1075 2180 2248 VSS VDD INVX4TR $T=69800 61000 1 0 $X=69460 $Y=57000
X1076 2592 2244 VSS VDD INVX4TR $T=73800 46600 1 0 $X=73460 $Y=42600
X1077 2582 3823 2579 VSS 3833 VDD OAI2BB1X1TR $T=70200 97000 1 0 $X=69860 $Y=93000
X1078 2260 2259 3915 VSS 2637 VDD OAI2BB1X1TR $T=86200 32200 0 0 $X=85860 $Y=31920
X1079 2635 2646 3948 VSS 2662 VDD OAI2BB1X1TR $T=91800 39400 1 0 $X=91460 $Y=35400
X1080 2677 2680 2674 VSS 3980 VDD OAI2BB1X1TR $T=99800 89800 0 180 $X=97060 $Y=85800
X1081 4039 2715 2311 VSS 2755 VDD OAI2BB1X1TR $T=105800 111400 0 0 $X=105460 $Y=111120
X1082 2625 2603 2606 3880 VDD VSS ADDHX1TR $T=74200 32200 0 0 $X=73860 $Y=31920
X1083 2664 2640 2634 3957 VDD VSS ADDHX1TR $T=89800 25000 1 0 $X=89460 $Y=21000
X1084 2707 2673 2282 2675 VDD VSS ADDHX1TR $T=92200 68200 1 0 $X=91860 $Y=64200
X1085 2251 3876 2614 VSS VDD 2607 ADDHXLTR $T=82600 82600 1 180 $X=77460 $Y=82320
X1086 2646 3927 2272 VSS VDD 2672 ADDHXLTR $T=86600 39400 0 0 $X=86260 $Y=39120
X1087 2618 3898 VSS 2260 VDD NAND2BX1TR $T=83000 39400 1 0 $X=82660 $Y=35400
X1088 3898 2618 VSS 3915 VDD NAND2BX1TR $T=83400 32200 0 0 $X=83060 $Y=31920
X1089 2665 2697 VSS 2758 VDD NAND2BX1TR $T=103400 111400 1 0 $X=103060 $Y=107400
X1090 2775 2757 VSS 2777 VDD NAND2BX1TR $T=118200 53800 1 0 $X=117860 $Y=49800
X1091 4200 2812 VSS 2824 VDD NAND2BX1TR $T=131800 97000 1 0 $X=131460 $Y=93000
X1092 2644 2648 VDD VSS 3938 ICV_268 $T=88600 53800 0 0 $X=88260 $Y=53520
X1093 3996 2716 VDD VSS 4009 ICV_268 $T=99800 17800 1 0 $X=99460 $Y=13800
X1094 2730 2759 VDD VSS 2776 ICV_268 $T=110200 118600 0 0 $X=109860 $Y=118320
X1095 2745 2721 VDD VSS 4119 ICV_268 $T=115400 104200 1 0 $X=115060 $Y=100200
X1096 4140 2759 VDD VSS 4147 ICV_268 $T=120200 68200 1 0 $X=119860 $Y=64200
X1097 4150 2716 VDD VSS 4175 ICV_268 $T=123400 17800 1 0 $X=123060 $Y=13800
X1098 4151 2716 VDD VSS 4176 ICV_268 $T=123400 25000 1 0 $X=123060 $Y=21000
X1099 2805 2364 VDD VSS 4182 ICV_268 $T=124200 89800 1 0 $X=123860 $Y=85800
X1100 4168 4196 VDD VSS 2821 ICV_268 $T=125000 118600 0 0 $X=124660 $Y=118320
X1101 2811 2810 VDD VSS 2834 ICV_268 $T=128600 118600 1 0 $X=128260 $Y=114600
X1102 2834 2812 VDD VSS 2849 ICV_268 $T=132200 111400 0 0 $X=131860 $Y=111120
X1103 2835 2812 VDD VSS 2841 ICV_268 $T=132200 118600 0 0 $X=131860 $Y=118320
X1104 2839 2812 VDD VSS 2858 ICV_268 $T=133000 75400 0 0 $X=132660 $Y=75120
X1105 2830 2812 VDD VSS 4208 ICV_268 $T=133400 61000 1 0 $X=133060 $Y=57000
X1106 2651 2633 VSS 2281 2656 VDD OAI21X2TR $T=89800 125800 1 0 $X=89460 $Y=121800
X1107 2786 2768 VSS 2749 2728 VDD OAI21X2TR $T=119000 82600 0 0 $X=118660 $Y=82320
X1108 VSS VDD 2702 2716 4034 ICV_269 $T=103000 17800 1 0 $X=102660 $Y=13800
X1109 VSS VDD 2750 2759 2774 ICV_269 $T=111000 125800 1 0 $X=110660 $Y=121800
X1110 VSS VDD 2312 2759 4098 ICV_269 $T=113400 118600 0 0 $X=113060 $Y=118320
X1111 VSS VDD 4162 2808 4171 ICV_269 $T=122200 32200 0 0 $X=121860 $Y=31920
X1112 VSS VDD 2804 2364 4181 ICV_269 $T=123800 82600 1 0 $X=123460 $Y=78600
X1113 VSS VDD 2365 2812 2822 ICV_269 $T=125400 125800 0 0 $X=125060 $Y=125520
X1114 VSS VDD 4179 4196 4190 ICV_269 $T=127000 111400 1 0 $X=126660 $Y=107400
X1115 VSS VDD 2833 2808 4201 ICV_269 $T=129400 46600 1 0 $X=129060 $Y=42600
X1116 VSS VDD 4201 2812 2843 ICV_269 $T=133000 46600 1 0 $X=132660 $Y=42600
X1117 VSS 4037 2724 4039 VDD NAND2X2TR $T=107000 111400 1 0 $X=106660 $Y=107400
X1118 VSS 4032 2766 2724 VDD NAND2X2TR $T=109800 97000 1 180 $X=107460 $Y=96720
X1119 VSS 2324 2735 4045 VDD NAND2X2TR $T=110600 104200 0 180 $X=108260 $Y=100200
X1120 VSS 4082 2785 2343 VDD NAND2X2TR $T=114200 39400 0 0 $X=113860 $Y=39120
X1121 2760 2761 2796 VDD VSS XNOR2X1TR $T=114600 25000 0 0 $X=114260 $Y=24720
X1122 2778 2766 2800 VDD VSS XNOR2X1TR $T=117800 82600 1 0 $X=117460 $Y=78600
X1123 4187 2372 2809 VDD VSS XNOR2X1TR $T=127800 53800 0 0 $X=127460 $Y=53520
.ENDS
***************************************
.SUBCKT SIGN_MEMFCIO8 VSS WE OE_ GTP
** N=33 EP=4 IP=0 FDC=3
*.CALIBRE ISOLATED NETS: VDD
D0 VSS WE tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1410 $Y=3050 $D=558
D1 VSS GTP tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1410 $Y=4760 $D=558
D2 VSS OE_ tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1410 $Y=8680 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMFCSA8 VSS GTP
** N=29 EP=2 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD
D0 VSS GTP tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1410 $Y=160 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMFCCAP
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD VSS
.ENDS
***************************************
.SUBCKT SIGN_MEMFCR
** N=12 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WLB WLT
.ENDS
***************************************
.SUBCKT SIGN_MEMFCCAP2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD VSS
.ENDS
***************************************
.SUBCKT SIGN_MEMFCUR
** N=12 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCCSTRAPR VSS WL 4
** N=7 EP=3 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD
M0 4 WL VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=90 $Y=1390 $D=103
.ENDS
***************************************
.SUBCKT ICV_42 1 3 4
** N=5 EP=3 IP=8 FDC=2
X0 1 3 5 SIGN_MEMFLCCSTRAPR $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 4 5 SIGN_MEMFLCCSTRAPR $T=0 3400 1 0 $X=-1000 $Y=700
.ENDS
***************************************
.SUBCKT SIGN_MEMFC1T
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS
.ENDS
***************************************
.SUBCKT SIGN_MEMFCBWM16 VSS D Q
** N=12 EP=3 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: VDD BWEN
D0 VSS D tdndsx AREA=1.024e-13 perim=1.28e-06 $X=15450 $Y=140 $D=558
D1 VSS Q tdndsx AREA=1.024e-13 perim=1.28e-06 $X=17840 $Y=140 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMIOX VSS VDD DPU DW DW_ SP Q DPN STUBWEI GTP OE_ D
** N=301 EP=12 IP=0 FDC=73
M0 13 VSS VSS VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=680 $D=103
M1 32 17 VSS VSS lpnfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=5110 $D=103
M2 VSS OE_ 22 VSS lpnfet w=1.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=450 $Y=8170 $D=103
M3 24 19 32 VSS lpnfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=500 $Y=5110 $D=103
M4 16 22 VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=980 $Y=7870 $D=103
M5 23 15 24 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1020 $Y=5110 $D=103
M6 VSS DW 23 VSS lpnfet w=1.6e-07 l=6.6e-07 m=1 par=1 nf=1 ngcon=1 $X=1540 $Y=5110 $D=103
M7 VSS 16 25 VSS lpnfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1800 $Y=8500 $D=103
M8 14 16 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2330 $Y=8170 $D=103
M9 DW 23 VSS VSS lpnfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2600 $Y=5110 $D=103
M10 27 25 14 VSS lpnfet w=2.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=8180 $D=103
M11 VSS 23 DW VSS lpnfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3080 $Y=5110 $D=103
M12 18 25 27 VSS lpnfet w=1.05e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3360 $Y=7400 $D=103
M13 DW_ 26 VSS VSS lpnfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3560 $Y=5110 $D=103
M14 27 25 18 VSS lpnfet w=1.05e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3840 $Y=7400 $D=103
M15 VSS 26 DW_ VSS lpnfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4040 $Y=5110 $D=103
M16 VSS DPU 27 VSS lpnfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4360 $Y=7400 $D=103
M17 26 DW_ VSS VSS lpnfet w=1.6e-07 l=6.6e-07 m=1 par=1 nf=1 ngcon=1 $X=4560 $Y=5110 $D=103
M18 27 DPU VSS VSS lpnfet w=9.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4840 $Y=7400 $D=103
M19 33 20 27 VSS lpnfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5320 $Y=7270 $D=103
M20 28 15 26 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5620 $Y=5110 $D=103
M21 VSS 29 33 VSS lpnfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5640 $Y=7270 $D=103
M22 34 21 28 VSS lpnfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6100 $Y=4880 $D=103
M23 29 27 VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6160 $Y=7770 $D=103
M24 VSS 17 34 VSS lpnfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6420 $Y=4880 $D=103
M25 19 30 VSS VSS lpnfet w=6.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6940 $Y=4880 $D=103
M26 VSS 19 21 VSS lpnfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7620 $Y=6480 $D=103
M27 30 D VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7650 $Y=940 $D=103
M28 VSS 31 17 VSS lpnfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8220 $Y=5680 $D=103
M29 VSS SP 20 VSS lpnfet w=1.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8220 $Y=7600 $D=103
M30 15 GTP VSS VSS lpnfet w=4.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8700 $Y=5680 $D=103
M31 Q 14 VSS VSS lpnfet w=1.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8820 $Y=6950 $D=103
M32 VSS STUBWEI 31 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9260 $Y=4770 $D=103
M33 VSS 14 Q VSS lpnfet w=1.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9300 $Y=6950 $D=103
M34 VDD OE_ 22 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=410 $Y=9560 $D=192
M35 24 19 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=700 $Y=3210 $D=192
M36 16 22 VDD VDD lppfet w=9.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=850 $Y=10520 $D=192
M37 23 GTP 24 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1220 $Y=3590 $D=192
M38 VDD 16 25 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1650 $Y=9560 $D=192
M39 VDD DW 23 VDD lppfet w=1.6e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=4120 $D=192
M40 VDD 17 24 VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1960 $Y=1160 $D=192
M41 18 25 VDD VDD lppfet w=1.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2170 $Y=9560 $D=192
M42 13 VSS VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=680 $D=192
M43 DW 23 VDD VDD lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=2160 $D=192
M44 27 16 18 VDD lppfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2690 $Y=9860 $D=192
M45 VDD VSS 13 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3000 $Y=680 $D=192
M46 VDD 23 DW VDD lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3000 $Y=2160 $D=192
M47 14 16 27 VDD lppfet w=1.32e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3210 $Y=9860 $D=192
M48 DW_ 26 VDD VDD lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3480 $Y=2160 $D=192
M49 27 16 14 VDD lppfet w=1.32e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3690 $Y=9860 $D=192
M50 VDD 26 DW_ VDD lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3960 $Y=2160 $D=192
M51 VDD DPN 27 VDD lppfet w=1.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4170 $Y=9860 $D=192
M52 26 DW_ VDD VDD lppfet w=1.6e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=4520 $Y=4060 $D=192
M53 27 DPN VDD VDD lppfet w=1.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4650 $Y=9860 $D=192
M54 VDD GTP 15 VDD lppfet w=5.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4930 $Y=2070 $D=192
M55 28 GTP 26 VDD lppfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5100 $Y=3360 $D=192
M56 VDD DPN 27 VDD lppfet w=1.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5130 $Y=9860 $D=192
M57 27 DPN VDD VDD lppfet w=1.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5610 $Y=9860 $D=192
M58 VDD 21 28 VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5620 $Y=2810 $D=192
M59 28 17 VDD VDD lppfet w=1.24e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6100 $Y=2810 $D=192
M60 35 SP 27 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6140 $Y=9330 $D=192
M61 VDD 29 35 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6460 $Y=9330 $D=192
M62 29 27 VDD VDD lppfet w=1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6980 $Y=9330 $D=192
M63 VDD 30 19 VDD lppfet w=1.26e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7040 $Y=3020 $D=192
M64 VDD SP 20 VDD lppfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7340 $Y=10640 $D=192
M65 21 19 VDD VDD lppfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7560 $Y=3400 $D=192
M66 30 D VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7640 $Y=1800 $D=192
M67 Q 18 VDD VDD lppfet w=1.79e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7860 $Y=9770 $D=192
M68 VDD 18 Q VDD lppfet w=1.79e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8340 $Y=9770 $D=192
M69 VDD 31 17 VDD lppfet w=1.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8500 $Y=3090 $D=192
M70 Q 18 VDD VDD lppfet w=1.79e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8820 $Y=9770 $D=192
M71 31 STUBWEI VDD VDD lppfet w=4.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9020 $Y=3500 $D=192
M72 VDD 18 Q VDD lppfet w=1.63e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9300 $Y=9770 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMFLIO VSS WE GTP OE_
** N=36 EP=4 IP=0 FDC=3
*.CALIBRE ISOLATED NETS: VDD
D0 VSS WE tdndsx AREA=1.024e-13 perim=1.28e-06 $X=4640 $Y=1840 $D=558
D1 VSS GTP tdndsx AREA=1.024e-13 perim=1.28e-06 $X=4640 $Y=3780 $D=558
D2 VSS OE_ tdndsx AREA=1.024e-13 perim=1.28e-06 $X=4640 $Y=7160 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMSA8 VSS VDD DPU SP DR DR_ DPN GTP
** N=263 EP=8 IP=0 FDC=57
*.CALIBRE ISOLATED NETS: DW DW_
M0 17 13 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=220 $Y=4450 $D=103
M1 VSS 17 18 VSS lpnfet w=6.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=5290 $D=103
M2 11 18 VSS VSS lpnfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=980 $Y=3310 $D=103
M3 VSS 15 DPU VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=6240 $D=103
M4 VSS 18 11 VSS lpnfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1460 $Y=3310 $D=103
M5 22 16 VSS VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1920 $Y=5320 $D=103
M6 23 11 VSS VSS lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1980 $Y=3310 $D=103
M7 20 13 22 VSS lpnfet w=1.66e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2320 $Y=5180 $D=103
M8 19 13 23 VSS lpnfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2380 $Y=3610 $D=103
M9 20 12 VDD VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3260 $Y=6690 $D=103
M10 15 14 20 VSS lpnfet w=2.31e-06 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=3780 $Y=3620 $D=103
M11 14 15 20 VSS lpnfet w=9.7e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=3780 $Y=6690 $D=103
M12 20 14 15 VSS lpnfet w=2.31e-06 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=4400 $Y=3620 $D=103
M13 20 15 14 VSS lpnfet w=9.7e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=4400 $Y=6690 $D=103
M14 VSS GTP 13 VSS lpnfet w=7.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4720 $Y=1650 $D=103
M15 14 15 20 VSS lpnfet w=2.31e-06 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=5020 $Y=3620 $D=103
M16 15 14 20 VSS lpnfet w=9.7e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=5020 $Y=6690 $D=103
M17 20 15 14 VSS lpnfet w=2.31e-06 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=5640 $Y=3620 $D=103
M18 20 14 15 VSS lpnfet w=9.7e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=5640 $Y=6690 $D=103
M19 VDD 12 20 VSS lpnfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6220 $Y=6690 $D=103
M20 VSS 19 SP VSS lpnfet w=1.06e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7100 $Y=3230 $D=103
M21 24 13 20 VSS lpnfet w=1.66e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7160 $Y=5180 $D=103
M22 VSS 16 24 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7560 $Y=5320 $D=103
M23 12 11 VSS VSS lpnfet w=2.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7620 $Y=3230 $D=103
M24 21 14 VSS VSS lpnfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8080 $Y=6240 $D=103
M25 VSS 12 16 VSS lpnfet w=2.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8300 $Y=4350 $D=103
M26 DPN 21 VSS VSS lpnfet w=1.46e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8820 $Y=4350 $D=103
M27 VSS 21 DPN VSS lpnfet w=1.46e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9300 $Y=4350 $D=103
M28 VDD 13 17 VDD lppfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=410 $Y=2020 $D=192
M29 DPU 15 VDD VDD lppfet w=1.64e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=450 $Y=7970 $D=192
M30 18 17 VDD VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=930 $Y=2200 $D=192
M31 DR 11 DR_ VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1390 $Y=8260 $D=192
M32 11 18 VDD VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1870 $Y=1340 $D=192
M33 VDD 11 DR VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1910 $Y=8260 $D=192
M34 VDD 18 11 VDD lppfet w=1.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2350 $Y=1340 $D=192
M35 DR 11 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2390 $Y=8260 $D=192
M36 19 11 VDD VDD lppfet w=7.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2870 $Y=1780 $D=192
M37 14 SP DR VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2910 $Y=8260 $D=192
M38 13 GTP VDD VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2980 $Y=620 $D=192
M39 VDD 13 19 VDD lppfet w=5.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3350 $Y=1780 $D=192
M40 DR SP 14 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3390 $Y=8260 $D=192
M41 VDD GTP 13 VDD lppfet w=5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3460 $Y=620 $D=192
M42 14 15 VDD VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4260 $Y=9190 $D=192
M43 15 16 14 VDD lppfet w=4.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4740 $Y=9190 $D=192
M44 VDD 14 15 VDD lppfet w=8.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5220 $Y=9190 $D=192
M45 15 SP DR_ VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6090 $Y=8260 $D=192
M46 SP 19 VDD VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6540 $Y=1100 $D=192
M47 DR_ SP 15 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6570 $Y=8260 $D=192
M48 VDD 19 SP VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7020 $Y=1100 $D=192
M49 VDD 11 DR_ VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7090 $Y=8260 $D=192
M50 12 11 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7500 $Y=1100 $D=192
M51 DR_ 11 VDD VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=8260 $D=192
M52 DR 11 DR_ VDD lppfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8090 $Y=8260 $D=192
M53 VDD 12 16 VDD lppfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8300 $Y=1960 $D=192
M54 DPN 21 VDD VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8820 $Y=1770 $D=192
M55 VDD 14 21 VDD lppfet w=1.64e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9030 $Y=7970 $D=192
M56 VDD 21 DPN VDD lppfet w=7.7e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9300 $Y=1770 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMFLSA VSS GTP
** N=32 EP=2 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD
D0 VSS GTP tdndsx AREA=1.024e-13 perim=1.28e-06 $X=4640 $Y=840 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMCD2 VSS VDD BL0 BL0_ BL1_ BL1 A0_ A0 GTP DR_ DR DW DW_ G0 G1
** N=409 EP=15 IP=0 FDC=60
*.CALIBRE ISOLATED NETS: DRSA DWSA STUBDW STUBDR_ STUBDR STUBDW_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0
M0 38 40 VSS VSS lpnfet w=1.75e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=25100 $D=103
M1 41 G0 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=200 $Y=23530 $D=103
M2 42 A0_ VSS VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=16020 $D=103
M3 BL0_ 30 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=920 $D=103
M4 30 32 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=4060 $D=103
M5 31 32 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=10940 $D=103
M6 BL0 31 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=12000 $D=103
M7 33 G1 41 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=520 $Y=23530 $D=103
M8 32 38 42 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=16020 $D=103
M9 VSS 40 38 VSS lpnfet w=1.75e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=25100 $D=103
M10 VSS 30 BL0_ VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=920 $D=103
M11 VSS 32 30 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=4060 $D=103
M12 VSS 32 31 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=10940 $D=103
M13 VSS 31 BL0 VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=12000 $D=103
M14 VSS 33 36 VSS lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=940 $Y=24300 $D=103
M15 BL1_ 34 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=920 $D=103
M16 34 39 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=4060 $D=103
M17 35 39 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=10940 $D=103
M18 BL1 35 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=12000 $D=103
M19 37 33 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1580 $Y=24300 $D=103
M20 43 38 39 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=16020 $D=103
M21 VSS 34 BL1_ VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=920 $D=103
M22 VSS 39 34 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=4060 $D=103
M23 VSS 39 35 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=10940 $D=103
M24 VSS 35 BL1 VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=12000 $D=103
M25 VSS A0 43 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1940 $Y=16020 $D=103
M26 GTP 36 37 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=23840 $D=103
M27 VSS 37 40 VSS lpnfet w=1.34e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=25280 $D=103
M28 BL1 38 VDD VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=28670 $D=192
M29 BL0 38 VDD VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=33850 $D=192
M30 32 A0_ VDD VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=19190 $D=192
M31 33 G0 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=22510 $D=192
M32 30 32 DW VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=5390 $D=192
M33 BL0_ 32 DR_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=6180 $D=192
M34 BL0 32 DR VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=8060 $D=192
M35 31 32 DW_ VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=9320 $D=192
M36 BL1_ 38 BL1 VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=28670 $D=192
M37 BL0_ 38 BL0 VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=33850 $D=192
M38 VDD 38 32 VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=820 $Y=19190 $D=192
M39 VDD G1 33 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=820 $Y=22510 $D=192
M40 DW 32 30 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=5390 $D=192
M41 DR_ 32 BL0_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=6180 $D=192
M42 DR 32 BL0 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=8060 $D=192
M43 DW_ 32 31 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=9320 $D=192
M44 VDD 38 BL1_ VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=28670 $D=192
M45 VDD 38 BL0_ VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=33850 $D=192
M46 34 39 DW VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=5390 $D=192
M47 BL1_ 39 DR_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=6180 $D=192
M48 BL1 39 DR VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=8060 $D=192
M49 35 39 DW_ VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=9320 $D=192
M50 39 38 VDD VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1460 $Y=19190 $D=192
M51 38 40 VDD VDD lppfet w=5.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1680 $Y=32970 $D=192
M52 40 37 VDD VDD lppfet w=2.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1780 $Y=28670 $D=192
M53 DW 39 34 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=5390 $D=192
M54 DR_ 39 BL1_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=6180 $D=192
M55 DR 39 BL1 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=8060 $D=192
M56 DW_ 39 35 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=9320 $D=192
M57 VDD A0 39 VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1940 $Y=19190 $D=192
M58 VDD 33 36 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=21720 $D=192
M59 GTP 33 37 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=22290 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMCD VSS VDD BL0 BL0_ BL1_ BL1 A0_ A0 GTP DR_ DR DW DW_ G0 G1
** N=409 EP=15 IP=0 FDC=60
*.CALIBRE ISOLATED NETS: DRSA DWSA STUBDW STUBDR_ STUBDR STUBDW_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0
M0 38 40 VSS VSS lpnfet w=1.75e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=25100 $D=103
M1 41 G0 VSS VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=200 $Y=23530 $D=103
M2 42 A0_ VSS VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=16020 $D=103
M3 BL0_ 30 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=920 $D=103
M4 30 32 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=4060 $D=103
M5 31 32 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=10940 $D=103
M6 BL0 31 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=12000 $D=103
M7 33 G1 41 VSS lpnfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=520 $Y=23530 $D=103
M8 32 38 42 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=16020 $D=103
M9 VSS 40 38 VSS lpnfet w=1.75e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=25100 $D=103
M10 VSS 30 BL0_ VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=920 $D=103
M11 VSS 32 30 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=4060 $D=103
M12 VSS 32 31 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=10940 $D=103
M13 VSS 31 BL0 VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=12000 $D=103
M14 VSS 33 36 VSS lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=940 $Y=24300 $D=103
M15 BL1_ 34 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=920 $D=103
M16 34 39 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=4060 $D=103
M17 35 39 VSS VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=10940 $D=103
M18 BL1 35 VSS VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=12000 $D=103
M19 37 33 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1580 $Y=24300 $D=103
M20 43 38 39 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=16020 $D=103
M21 VSS 34 BL1_ VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=920 $D=103
M22 VSS 39 34 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=4060 $D=103
M23 VSS 39 35 VSS lpnfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=10940 $D=103
M24 VSS 35 BL1 VSS lpnfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=12000 $D=103
M25 VSS A0 43 VSS lpnfet w=1.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1940 $Y=16020 $D=103
M26 GTP 36 37 VSS lpnfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=23840 $D=103
M27 VSS 37 40 VSS lpnfet w=1.34e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=25280 $D=103
M28 BL1 38 VDD VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=28670 $D=192
M29 BL0 38 VDD VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=33850 $D=192
M30 32 A0_ VDD VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=19190 $D=192
M31 33 G0 VDD VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=340 $Y=22510 $D=192
M32 30 32 DW VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=5390 $D=192
M33 BL0_ 32 DR_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=6180 $D=192
M34 BL0 32 DR VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=8060 $D=192
M35 31 32 DW_ VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=420 $Y=9320 $D=192
M36 BL1_ 38 BL1 VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=28670 $D=192
M37 BL0_ 38 BL0 VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=33850 $D=192
M38 VDD 38 32 VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=820 $Y=19190 $D=192
M39 VDD G1 33 VDD lppfet w=3.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=820 $Y=22510 $D=192
M40 DW 32 30 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=5390 $D=192
M41 DR_ 32 BL0_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=6180 $D=192
M42 DR 32 BL0 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=8060 $D=192
M43 DW_ 32 31 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=900 $Y=9320 $D=192
M44 VDD 38 BL1_ VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=28670 $D=192
M45 VDD 38 BL0_ VDD lppfet w=5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=33850 $D=192
M46 34 39 DW VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=5390 $D=192
M47 BL1_ 39 DR_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=6180 $D=192
M48 BL1 39 DR VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=8060 $D=192
M49 35 39 DW_ VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1380 $Y=9320 $D=192
M50 39 38 VDD VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1460 $Y=19190 $D=192
M51 38 40 VDD VDD lppfet w=5.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1680 $Y=32970 $D=192
M52 40 37 VDD VDD lppfet w=2.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1780 $Y=28670 $D=192
M53 DW 39 34 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=5390 $D=192
M54 DR_ 39 BL1_ VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=6180 $D=192
M55 DR 39 BL1 VDD lppfet w=1.08e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=8060 $D=192
M56 DW_ 39 35 VDD lppfet w=6.1e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1860 $Y=9320 $D=192
M57 VDD A0 39 VDD lppfet w=1.48e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1940 $Y=19190 $D=192
M58 VDD 33 36 VDD lppfet w=3.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=21720 $D=192
M59 GTP 33 37 VDD lppfet w=7.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2100 $Y=22290 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMMUX_CD_ODD VSS VDD STUBDW_0 STUBDR_0 STUBDR__0 STUBDW__0 YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 A0_ A0 GTP BL0_0 BL0__0 BL1_0
+ BL1__0 BL0_2 BL0__2 BL1_2 BL1__2 BL0_4 BL0__4 BL1_4 BL1__4 BL0_6 BL0__6 BL1_6 BL1__6 BL0_1 BL0__1 BL1_1 BL1__1 BL0_3 BL0__3 BL1_3
+ BL1__3 BL0_5 BL0__5 BL1_5 BL1__5 BL0_7 BL0__7 BL1_7 BL1__7
** N=65 EP=49 IP=232 FDC=480
*.CALIBRE ISOLATED NETS: DRSA_0 DWSA_0 DRSA_2 DWSA_2 DRSA_4 DWSA_4 DRSA_1 DWSA_1 DRSA_3 DWSA_3 DRSA_5 DWSA_5 STUBDW_1 STUBDR__1 STUBDR_1 STUBDW__1
X0 VSS VDD BL0_0 BL0__0 BL1__0 BL1_0 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 VDD YP1_3 SIGN_MEMCD2 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS VDD BL0_2 BL0__2 BL1__2 BL1_2 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 VDD YP1_1 SIGN_MEMCD2 $T=4800 0 0 0 $X=3800 $Y=-1000
X2 VSS VDD BL0_4 BL0__4 BL1__4 BL1_4 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 YP0_3 VDD SIGN_MEMCD2 $T=9600 0 0 0 $X=8600 $Y=-1000
X3 VSS VDD BL0_6 BL0__6 BL1__6 BL1_6 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 YP0_1 VDD SIGN_MEMCD2 $T=14400 0 0 0 $X=13400 $Y=-1000
X4 VSS VDD BL0_1 BL0__1 BL1__1 BL1_1 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 VDD YP1_2 SIGN_MEMCD $T=4800 0 1 180 $X=1400 $Y=-1000
X5 VSS VDD BL0_3 BL0__3 BL1__3 BL1_3 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 VDD YP1_0 SIGN_MEMCD $T=9600 0 1 180 $X=6200 $Y=-1000
X6 VSS VDD BL0_5 BL0__5 BL1__5 BL1_5 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 YP0_2 VDD SIGN_MEMCD $T=14400 0 1 180 $X=11000 $Y=-1000
X7 VSS VDD BL0_7 BL0__7 BL1__7 BL1_7 A0_ A0 GTP STUBDR__0 STUBDR_0 STUBDW_0 STUBDW__0 YP0_0 VDD SIGN_MEMCD $T=19200 0 1 180 $X=15800 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_62 1 2 3 4 5 6 7 8 9 10 11 12 13 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=62 EP=55 IP=100 FDC=616
X0 1 3 4 SIGN_MEMFCBWM16 $T=0 0 0 270 $X=-1000 $Y=-20200
X1 1 2 60 5 6 61 4 62 9 10 11 3 SIGN_MEMIOX $T=1200 -9600 0 270 $X=200 $Y=-20200
X2 1 9 10 11 SIGN_MEMFLIO $T=1200 0 0 270 $X=200 $Y=-10600
X3 1 2 60 61 7 8 62 12 SIGN_MEMSA8 $T=12470 -9600 0 270 $X=11470 $Y=-20200
X4 1 12 SIGN_MEMFLSA $T=12470 0 0 270 $X=11470 $Y=-10600
X5 1 2 5 7 8 6 19 20 21 22 23 24 25 26 13 18 27 28 29 30
+ 31 36 37 38 39 44 45 46 47 52 53 54 55 35 34 33 32 43 42 41
+ 40 51 50 49 48 59 58 57 56
+ SIGN_MEMMUX_CD_ODD $T=22810 0 0 270 $X=21810 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_136 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53
** N=53 EP=53 IP=59 FDC=616
X0 4 1 3 2 18 21 20 19 6 5 7 5 9 8 10 11 12 13 14 15
+ 16 17 5 53 52 51 50 49 48 47 46 45 44 43 42 41 40 39 38 37
+ 36 35 34 33 32 31 30 29 28 27 26 25 24 23 22
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPEG
** N=5 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL BL_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPOP
** N=5 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD BL VSS BL_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPEP
** N=5 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD BL BL_ VSS
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPOG
** N=5 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL BL_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAP_ROW16
** N=34 EP=0 IP=64 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL_0 BL__0 BL_4 BL__4 BL_8 BL__8 BL_12 BL__12 BL_1 BL__1 BL_5 BL__5 BL_9 BL__9 BL_13 BL__13 BL_2 BL__2
*+ BL_6 BL__6 BL_10 BL__10 BL_14 BL__14 BL_3 BL__3 BL_7 BL__7 BL_11 BL__11 BL_15 BL__15
.ENDS
***************************************
.SUBCKT ICV_60
** N=34 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_135
** N=34 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT A8FCELLE_D_LP 2 4 8 9
** N=17 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 4 9 8 4 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=380 $Y=850 $D=103
M1 9 8 4 4 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=850 $D=103
M2 2 9 8 2 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=370 $Y=260 $D=192
M3 9 8 2 2 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=260 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMCCEG VSS VDD 9 10
** N=10 EP=4 IP=9 FDC=4
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL BL_ WP
X0 VDD VSS 9 10 A8FCELLE_D_LP $T=0 0 0 0 $X=-220 $Y=-470
.ENDS
***************************************
.SUBCKT A8FCELLO_D_LP 2 4 8 9
** N=17 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 2 9 8 2 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=380 $Y=850 $D=103
M1 9 8 2 2 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=850 $D=103
M2 4 9 8 4 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=370 $Y=260 $D=192
M3 9 8 4 4 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=260 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMCCOP VDD VSS 9 10
** N=10 EP=4 IP=9 FDC=4
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL BL_ WP
X0 VSS VDD 9 10 A8FCELLO_D_LP $T=0 0 0 0 $X=-220 $Y=-470
.ENDS
***************************************
.SUBCKT SIGN_MEMCCEP VDD VSS 9 10
** N=10 EP=4 IP=9 FDC=4
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL BL_ WP
X0 VDD VSS 9 10 A8FCELLE_D_LP $T=0 0 0 0 $X=-220 $Y=-470
.ENDS
***************************************
.SUBCKT SIGN_MEMCCOG VSS VDD 9 10
** N=10 EP=4 IP=9 FDC=4
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL BL_ WP
X0 VSS VDD 9 10 A8FCELLO_D_LP $T=0 0 0 0 $X=-220 $Y=-470
.ENDS
***************************************
.SUBCKT SIGN_MEMBIT_MUX_0 VSS VDD 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100
** N=100 EP=34 IP=160 FDC=64
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL_0 BL__0 BL_4 BL__4 BL_8 BL__8 BL_12 BL__12 BL_1 BL__1 BL_5 BL__5 BL_9 BL__9 BL_13 BL__13 BL_2 BL__2 BL_6
*+ BL__6 BL_10 BL__10 BL_14 BL__14 BL_3 BL__3 BL_7 BL__7 BL_11 BL__11 BL_15 BL__15 WP
X0 VSS VDD 69 70 SIGN_MEMCCEG $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS VDD 71 72 SIGN_MEMCCEG $T=4800 0 0 0 $X=3800 $Y=-1000
X2 VSS VDD 73 74 SIGN_MEMCCEG $T=9600 0 0 0 $X=8600 $Y=-1000
X3 VSS VDD 75 76 SIGN_MEMCCEG $T=14400 0 0 0 $X=13400 $Y=-1000
X4 VDD VSS 77 78 SIGN_MEMCCOP $T=2400 0 1 180 $X=200 $Y=-1000
X5 VDD VSS 79 80 SIGN_MEMCCOP $T=7200 0 1 180 $X=5000 $Y=-1000
X6 VDD VSS 81 82 SIGN_MEMCCOP $T=12000 0 1 180 $X=9800 $Y=-1000
X7 VDD VSS 83 84 SIGN_MEMCCOP $T=16800 0 1 180 $X=14600 $Y=-1000
X8 VDD VSS 85 86 SIGN_MEMCCEP $T=2400 0 0 0 $X=1400 $Y=-1000
X9 VDD VSS 87 88 SIGN_MEMCCEP $T=7200 0 0 0 $X=6200 $Y=-1000
X10 VDD VSS 89 90 SIGN_MEMCCEP $T=12000 0 0 0 $X=11000 $Y=-1000
X11 VDD VSS 91 92 SIGN_MEMCCEP $T=16800 0 0 0 $X=15800 $Y=-1000
X12 VSS VDD 93 94 SIGN_MEMCCOG $T=4800 0 1 180 $X=2600 $Y=-1000
X13 VSS VDD 95 96 SIGN_MEMCCOG $T=9600 0 1 180 $X=7400 $Y=-1000
X14 VSS VDD 97 98 SIGN_MEMCCOG $T=14400 0 1 180 $X=12200 $Y=-1000
X15 VSS VDD 99 100 SIGN_MEMCCOG $T=19200 0 1 180 $X=17000 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMBIT_MUX_1 VSS VDD 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100
** N=100 EP=34 IP=160 FDC=64
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL_0 BL__0 BL_4 BL__4 BL_8 BL__8 BL_12 BL__12 BL_1 BL__1 BL_5 BL__5 BL_9 BL__9 BL_13 BL__13 BL_2 BL__2 BL_6
*+ BL__6 BL_10 BL__10 BL_14 BL__14 BL_3 BL__3 BL_7 BL__7 BL_11 BL__11 BL_15 BL__15 WP
X0 VSS VDD 69 70 SIGN_MEMCCEG $T=1200 1700 0 180 $X=-1000 $Y=-1000
X1 VSS VDD 71 72 SIGN_MEMCCEG $T=6000 1700 0 180 $X=3800 $Y=-1000
X2 VSS VDD 73 74 SIGN_MEMCCEG $T=10800 1700 0 180 $X=8600 $Y=-1000
X3 VSS VDD 75 76 SIGN_MEMCCEG $T=15600 1700 0 180 $X=13400 $Y=-1000
X4 VDD VSS 77 78 SIGN_MEMCCOP $T=1200 1700 1 0 $X=200 $Y=-1000
X5 VDD VSS 79 80 SIGN_MEMCCOP $T=6000 1700 1 0 $X=5000 $Y=-1000
X6 VDD VSS 81 82 SIGN_MEMCCOP $T=10800 1700 1 0 $X=9800 $Y=-1000
X7 VDD VSS 83 84 SIGN_MEMCCOP $T=15600 1700 1 0 $X=14600 $Y=-1000
X8 VDD VSS 85 86 SIGN_MEMCCEP $T=3600 1700 0 180 $X=1400 $Y=-1000
X9 VDD VSS 87 88 SIGN_MEMCCEP $T=8400 1700 0 180 $X=6200 $Y=-1000
X10 VDD VSS 89 90 SIGN_MEMCCEP $T=13200 1700 0 180 $X=11000 $Y=-1000
X11 VDD VSS 91 92 SIGN_MEMCCEP $T=18000 1700 0 180 $X=15800 $Y=-1000
X12 VSS VDD 93 94 SIGN_MEMCCOG $T=3600 1700 1 0 $X=2600 $Y=-1000
X13 VSS VDD 95 96 SIGN_MEMCCOG $T=8400 1700 1 0 $X=7400 $Y=-1000
X14 VSS VDD 97 98 SIGN_MEMCCOG $T=13200 1700 1 0 $X=12200 $Y=-1000
X15 VSS VDD 99 100 SIGN_MEMCCOG $T=18000 1700 1 0 $X=17000 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMBIT_MUX_2 VSS VDD 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100
** N=100 EP=34 IP=160 FDC=64
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL_0 BL__0 BL_4 BL__4 BL_8 BL__8 BL_12 BL__12 BL_1 BL__1 BL_5 BL__5 BL_9 BL__9 BL_13 BL__13 BL_2 BL__2 BL_6
*+ BL__6 BL_10 BL__10 BL_14 BL__14 BL_3 BL__3 BL_7 BL__7 BL_11 BL__11 BL_15 BL__15 WP
X0 VSS VDD 69 70 SIGN_MEMCCEG $T=1200 0 1 180 $X=-1000 $Y=-1000
X1 VSS VDD 71 72 SIGN_MEMCCEG $T=6000 0 1 180 $X=3800 $Y=-1000
X2 VSS VDD 73 74 SIGN_MEMCCEG $T=10800 0 1 180 $X=8600 $Y=-1000
X3 VSS VDD 75 76 SIGN_MEMCCEG $T=15600 0 1 180 $X=13400 $Y=-1000
X4 VDD VSS 77 78 SIGN_MEMCCOP $T=1200 0 0 0 $X=200 $Y=-1000
X5 VDD VSS 79 80 SIGN_MEMCCOP $T=6000 0 0 0 $X=5000 $Y=-1000
X6 VDD VSS 81 82 SIGN_MEMCCOP $T=10800 0 0 0 $X=9800 $Y=-1000
X7 VDD VSS 83 84 SIGN_MEMCCOP $T=15600 0 0 0 $X=14600 $Y=-1000
X8 VDD VSS 85 86 SIGN_MEMCCEP $T=3600 0 1 180 $X=1400 $Y=-1000
X9 VDD VSS 87 88 SIGN_MEMCCEP $T=8400 0 1 180 $X=6200 $Y=-1000
X10 VDD VSS 89 90 SIGN_MEMCCEP $T=13200 0 1 180 $X=11000 $Y=-1000
X11 VDD VSS 91 92 SIGN_MEMCCEP $T=18000 0 1 180 $X=15800 $Y=-1000
X12 VSS VDD 93 94 SIGN_MEMCCOG $T=3600 0 0 0 $X=2600 $Y=-1000
X13 VSS VDD 95 96 SIGN_MEMCCOG $T=8400 0 0 0 $X=7400 $Y=-1000
X14 VSS VDD 97 98 SIGN_MEMCCOG $T=13200 0 0 0 $X=12200 $Y=-1000
X15 VSS VDD 99 100 SIGN_MEMCCOG $T=18000 0 0 0 $X=17000 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMBIT_MUX_3 VSS VDD 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100
** N=100 EP=34 IP=160 FDC=64
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL BL_0 BL__0 BL_4 BL__4 BL_8 BL__8 BL_12 BL__12 BL_1 BL__1 BL_5 BL__5 BL_9 BL__9 BL_13 BL__13 BL_2 BL__2 BL_6
*+ BL__6 BL_10 BL__10 BL_14 BL__14 BL_3 BL__3 BL_7 BL__7 BL_11 BL__11 BL_15 BL__15 WP
X0 VSS VDD 69 70 SIGN_MEMCCEG $T=0 1700 1 0 $X=-1000 $Y=-1000
X1 VSS VDD 71 72 SIGN_MEMCCEG $T=4800 1700 1 0 $X=3800 $Y=-1000
X2 VSS VDD 73 74 SIGN_MEMCCEG $T=9600 1700 1 0 $X=8600 $Y=-1000
X3 VSS VDD 75 76 SIGN_MEMCCEG $T=14400 1700 1 0 $X=13400 $Y=-1000
X4 VDD VSS 77 78 SIGN_MEMCCOP $T=2400 1700 0 180 $X=200 $Y=-1000
X5 VDD VSS 79 80 SIGN_MEMCCOP $T=7200 1700 0 180 $X=5000 $Y=-1000
X6 VDD VSS 81 82 SIGN_MEMCCOP $T=12000 1700 0 180 $X=9800 $Y=-1000
X7 VDD VSS 83 84 SIGN_MEMCCOP $T=16800 1700 0 180 $X=14600 $Y=-1000
X8 VDD VSS 85 86 SIGN_MEMCCEP $T=2400 1700 1 0 $X=1400 $Y=-1000
X9 VDD VSS 87 88 SIGN_MEMCCEP $T=7200 1700 1 0 $X=6200 $Y=-1000
X10 VDD VSS 89 90 SIGN_MEMCCEP $T=12000 1700 1 0 $X=11000 $Y=-1000
X11 VDD VSS 91 92 SIGN_MEMCCEP $T=16800 1700 1 0 $X=15800 $Y=-1000
X12 VSS VDD 93 94 SIGN_MEMCCOG $T=4800 1700 0 180 $X=2600 $Y=-1000
X13 VSS VDD 95 96 SIGN_MEMCCOG $T=9600 1700 0 180 $X=7400 $Y=-1000
X14 VSS VDD 97 98 SIGN_MEMCCOG $T=14400 1700 0 180 $X=12200 $Y=-1000
X15 VSS VDD 99 100 SIGN_MEMCCOG $T=19200 1700 0 180 $X=17000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_43 1 2 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25
+ 26 27 28 29 30 31 32 33 34 35 36 37 39 40 41 42 107 108 109 110
+ 111 112 113 114
** N=234 EP=44 IP=400 FDC=376
*.SEEDPROM
M0 8 39 115 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1390 $D=103
M1 145 40 8 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1880 $D=103
M2 8 41 175 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=4790 $D=103
M3 205 42 8 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=5280 $D=103
M4 9 39 123 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=1290 $Y=1390 $D=103
M5 152 40 9 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=1290 $Y=1880 $D=103
M6 9 41 182 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=1290 $Y=4790 $D=103
M7 213 42 9 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=1290 $Y=5280 $D=103
M8 10 39 122 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2150 $Y=1390 $D=103
M9 153 40 10 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2150 $Y=1880 $D=103
M10 10 41 183 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2150 $Y=4790 $D=103
M11 212 42 10 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2150 $Y=5280 $D=103
M12 11 39 130 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2490 $Y=1390 $D=103
M13 161 40 11 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2490 $Y=1880 $D=103
M14 11 41 191 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2490 $Y=4790 $D=103
M15 220 42 11 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=2490 $Y=5280 $D=103
M16 12 39 131 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3350 $Y=1390 $D=103
M17 160 40 12 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3350 $Y=1880 $D=103
M18 12 41 190 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3350 $Y=4790 $D=103
M19 221 42 12 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3350 $Y=5280 $D=103
M20 13 39 139 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3690 $Y=1390 $D=103
M21 168 40 13 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3690 $Y=1880 $D=103
M22 13 41 198 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3690 $Y=4790 $D=103
M23 229 42 13 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=3690 $Y=5280 $D=103
M24 14 39 138 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4550 $Y=1390 $D=103
M25 169 40 14 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4550 $Y=1880 $D=103
M26 14 41 199 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4550 $Y=4790 $D=103
M27 228 42 14 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4550 $Y=5280 $D=103
M28 15 39 116 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4890 $Y=1390 $D=103
M29 147 40 15 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4890 $Y=1880 $D=103
M30 15 41 177 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4890 $Y=4790 $D=103
M31 206 42 15 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=4890 $Y=5280 $D=103
M32 16 39 117 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=5750 $Y=1390 $D=103
M33 146 40 16 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=5750 $Y=1880 $D=103
M34 16 41 176 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=5750 $Y=4790 $D=103
M35 207 42 16 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=5750 $Y=5280 $D=103
M36 17 39 125 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6090 $Y=1390 $D=103
M37 154 40 17 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6090 $Y=1880 $D=103
M38 17 41 184 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6090 $Y=4790 $D=103
M39 215 42 17 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6090 $Y=5280 $D=103
M40 18 39 124 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6950 $Y=1390 $D=103
M41 155 40 18 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6950 $Y=1880 $D=103
M42 18 41 185 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6950 $Y=4790 $D=103
M43 214 42 18 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=6950 $Y=5280 $D=103
M44 19 39 132 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=7290 $Y=1390 $D=103
M45 163 40 19 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=7290 $Y=1880 $D=103
M46 19 41 193 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=7290 $Y=4790 $D=103
M47 222 42 19 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=7290 $Y=5280 $D=103
M48 20 39 133 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8150 $Y=1390 $D=103
M49 162 40 20 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8150 $Y=1880 $D=103
M50 20 41 192 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8150 $Y=4790 $D=103
M51 223 42 20 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8150 $Y=5280 $D=103
M52 21 39 141 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8490 $Y=1390 $D=103
M53 170 40 21 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8490 $Y=1880 $D=103
M54 21 41 200 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8490 $Y=4790 $D=103
M55 231 42 21 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=8490 $Y=5280 $D=103
M56 22 39 140 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9350 $Y=1390 $D=103
M57 171 40 22 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9350 $Y=1880 $D=103
M58 22 41 201 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9350 $Y=4790 $D=103
M59 230 42 22 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9350 $Y=5280 $D=103
M60 23 39 118 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9690 $Y=1390 $D=103
M61 149 40 23 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9690 $Y=1880 $D=103
M62 23 41 179 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9690 $Y=4790 $D=103
M63 208 42 23 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=9690 $Y=5280 $D=103
M64 24 39 119 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10550 $Y=1390 $D=103
M65 148 40 24 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10550 $Y=1880 $D=103
M66 24 41 178 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10550 $Y=4790 $D=103
M67 209 42 24 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10550 $Y=5280 $D=103
M68 25 39 127 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10890 $Y=1390 $D=103
M69 156 40 25 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10890 $Y=1880 $D=103
M70 25 41 186 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10890 $Y=4790 $D=103
M71 217 42 25 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=10890 $Y=5280 $D=103
M72 26 39 126 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=11750 $Y=1390 $D=103
M73 157 40 26 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=11750 $Y=1880 $D=103
M74 26 41 187 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=11750 $Y=4790 $D=103
M75 216 42 26 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=11750 $Y=5280 $D=103
M76 27 39 134 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12090 $Y=1390 $D=103
M77 165 40 27 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12090 $Y=1880 $D=103
M78 27 41 195 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12090 $Y=4790 $D=103
M79 224 42 27 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12090 $Y=5280 $D=103
M80 28 39 135 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12950 $Y=1390 $D=103
M81 164 40 28 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12950 $Y=1880 $D=103
M82 28 41 194 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12950 $Y=4790 $D=103
M83 225 42 28 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12950 $Y=5280 $D=103
M84 29 39 143 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13290 $Y=1390 $D=103
M85 172 40 29 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13290 $Y=1880 $D=103
M86 29 41 202 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13290 $Y=4790 $D=103
M87 233 42 29 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13290 $Y=5280 $D=103
M88 30 39 142 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14150 $Y=1390 $D=103
M89 173 40 30 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14150 $Y=1880 $D=103
M90 30 41 203 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14150 $Y=4790 $D=103
M91 232 42 30 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14150 $Y=5280 $D=103
M92 31 39 120 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14490 $Y=1390 $D=103
M93 151 40 31 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14490 $Y=1880 $D=103
M94 31 41 181 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14490 $Y=4790 $D=103
M95 210 42 31 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14490 $Y=5280 $D=103
M96 32 39 121 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15350 $Y=1390 $D=103
M97 150 40 32 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15350 $Y=1880 $D=103
M98 32 41 180 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15350 $Y=4790 $D=103
M99 211 42 32 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15350 $Y=5280 $D=103
M100 33 39 129 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15690 $Y=1390 $D=103
M101 158 40 33 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15690 $Y=1880 $D=103
M102 33 41 188 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15690 $Y=4790 $D=103
M103 219 42 33 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15690 $Y=5280 $D=103
M104 34 39 128 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16550 $Y=1390 $D=103
M105 159 40 34 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16550 $Y=1880 $D=103
M106 34 41 189 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16550 $Y=4790 $D=103
M107 218 42 34 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16550 $Y=5280 $D=103
M108 35 39 136 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16890 $Y=1390 $D=103
M109 167 40 35 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16890 $Y=1880 $D=103
M110 35 41 197 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16890 $Y=4790 $D=103
M111 226 42 35 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16890 $Y=5280 $D=103
M112 36 39 137 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17750 $Y=1390 $D=103
M113 166 40 36 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17750 $Y=1880 $D=103
M114 36 41 196 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17750 $Y=4790 $D=103
M115 227 42 36 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17750 $Y=5280 $D=103
M116 37 39 144 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18090 $Y=1390 $D=103
M117 174 40 37 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18090 $Y=1880 $D=103
M118 37 41 204 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18090 $Y=4790 $D=103
M119 234 42 37 1 lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18090 $Y=5280 $D=103
X120 1 2 107 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131
+ 132 133 134 135 136 137 138 139 140 141 142 143 108 144
+ SIGN_MEMBIT_MUX_0 $T=0 0 0 0 $X=-1000 $Y=-1000
X121 1 2 145 109 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 110
+ SIGN_MEMBIT_MUX_1 $T=0 1700 0 0 $X=-1000 $Y=700
X122 1 2 175 111 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191
+ 192 193 194 195 196 197 198 199 200 201 202 203 204 112
+ SIGN_MEMBIT_MUX_2 $T=0 3400 0 0 $X=-1000 $Y=2400
X123 1 2 113 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 114 234
+ SIGN_MEMBIT_MUX_3 $T=0 5100 0 0 $X=-1000 $Y=4100
.ENDS
***************************************
.SUBCKT ICV_44 1 2 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 40 41 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
** N=66 EP=56 IP=100 FDC=752
*.SEEDPROM
X0 1 2 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 40 41 43 44 45 46 51 52 53 54
+ 55 56 57 58
+ ICV_43 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 2 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 40 41 47 48 49 50 59 60 61 62
+ 63 64 65 66
+ ICV_43 $T=0 6800 0 0 $X=-1000 $Y=5800
.ENDS
***************************************
.SUBCKT ICV_45 1 2 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 51 52 53 54 55 56 57 58
+ 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78
+ 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98
** N=98 EP=80 IP=132 FDC=1504
*.SEEDPROM
X0 1 2 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 51 52 53 54 55 56 57 58
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ ICV_44 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 2 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 59 60 61 62 63 64 65 66
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98
+ ICV_44 $T=0 13600 0 0 $X=-1000 $Y=12600
.ENDS
***************************************
.SUBCKT ICV_46 1 2 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 67 68 69 70 71 72 73 74
+ 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94
+ 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114
+ 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134
+ 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154
+ 155 156 157 158 159 160 161 162
** N=162 EP=128 IP=196 FDC=3008
*.SEEDPROM
X0 1 2 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 67 68 69 70 71 72 73 74
+ 75 76 77 78 79 80 81 82 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ ICV_45 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 2 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ ICV_45 $T=0 27200 0 0 $X=-1000 $Y=26200
.ENDS
***************************************
.SUBCKT SIGN_MEMBIT_COL VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_0 WP_1 WP_2 WP_3 WP_4 WP_5 WP_6 WP_7
+ WP_8 WP_9 WP_10 WP_11 WP_12 WP_13 WP_14 WP_15 WP_16 WP_17 WP_18 WP_19 WP_20 WP_21 WP_22 WP_23 WP_24 WP_25 WP_26 WP_27
+ WP_28 WP_29 WP_30 WP_31 WP_32 WP_33 WP_34 WP_35 WP_36 WP_37 WP_38 WP_39 WP_40 WP_41 WP_42 WP_43 WP_44 WP_45 WP_46 WP_47
+ WP_48 WP_49 WP_50 WP_51 WP_52 WP_53 WP_54 WP_55 WP_56 WP_57 WP_58 WP_59 WP_60 WP_61 WP_62 WP_63 WP_64 WP_65 WP_66 WP_67
+ WP_68 WP_69 WP_70 WP_71 WP_72 WP_73 WP_74 WP_75 WP_76 WP_77 WP_78 WP_79 WP_80 WP_81 WP_82 WP_83 WP_84 WP_85 WP_86 WP_87
+ WP_88 WP_89 WP_90 WP_91 WP_92 WP_93 WP_94 WP_95 WP_96 WP_97 WP_98 WP_99 WP_100 WP_101 WP_102 WP_103 WP_104 WP_105 WP_106 WP_107
+ WP_108 WP_109 WP_110 WP_111 WP_112 WP_113 WP_114 WP_115 WP_116 WP_117 WP_118 WP_119 WP_120 WP_121 WP_122 WP_123 WP_124 WP_125 WP_126 WP_127
+ WP_128 WP_129 WP_130 WP_131 WP_132 WP_133 WP_134 WP_135 WP_136 WP_137 WP_138 WP_139 WP_140 WP_141 WP_142 WP_143 WP_144 WP_145 WP_146 WP_147
+ WP_148 WP_149 WP_150 WP_151 WP_152 WP_153 WP_154 WP_155 WP_156 WP_157 WP_158 WP_159 WP_160 WP_161 WP_162 WP_163 WP_164 WP_165 WP_166 WP_167
+ WP_168 WP_169 WP_170 WP_171 WP_172 WP_173 WP_174 WP_175 WP_176 WP_177 WP_178 WP_179 WP_180 WP_181 WP_182 WP_183 WP_184 WP_185 WP_186 WP_187
+ WP_188 WP_189 WP_190 WP_191 WP_192 WP_193 WP_194 WP_195 WP_196 WP_197 WP_198 WP_199 WP_200 WP_201 WP_202 WP_203 WP_204 WP_205 WP_206 WP_207
+ WP_208 WP_209 WP_210 WP_211 WP_212 WP_213 WP_214 WP_215 WP_216 WP_217 WP_218 WP_219 WP_220 WP_221 WP_222 WP_223 WP_224 WP_225 WP_226 WP_227
+ WP_228 WP_229 WP_230 WP_231 WP_232 WP_233 WP_234 WP_235 WP_236 WP_237 WP_238 WP_239 WP_240 WP_241 WP_242 WP_243 WP_244 WP_245 WP_246 WP_247
+ WP_248 WP_249 WP_250 WP_251 WP_252 WP_253 WP_254 WP_255 547 548 549 550 551 552 553 554 555 556 557 558
+ 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578
+ 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598
+ 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618
+ 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658
+ 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678
+ 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
+ 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718
+ 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738
+ 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758
+ 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778
+ 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798
+ 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878
+ 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898
+ 899 900 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918
+ 919 920 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938
+ 939 940 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958
+ 959 960 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978
+ 979 980 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998
+ 999 1000 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018
+ 1019 1020 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038
+ 1039 1040 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058
** N=1058 EP=800 IP=1296 FDC=24064
*.SEEDPROM
*.CALIBRE ISOLATED NETS: WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19
*+ WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39
*+ WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 WL_59
*+ WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79
*+ WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98 WL_99
*+ WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 WL_119
*+ WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138 WL_139
*+ WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158 WL_159
*+ WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178 WL_179
*+ WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198 WL_199
*+ WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218 WL_219
*+ WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238 WL_239
*+ WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255 BL_0 BL_15
X0 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_0 WP_1 WP_2 WP_3 WP_4 WP_5 WP_6 WP_7
+ WP_8 WP_9 WP_10 WP_11 WP_12 WP_13 WP_14 WP_15 WP_16 WP_17 WP_18 WP_19 WP_20 WP_21 WP_22 WP_23 WP_24 WP_25 WP_26 WP_27
+ WP_28 WP_29 WP_30 WP_31 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610
+ ICV_46 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_32 WP_33 WP_34 WP_35 WP_36 WP_37 WP_38 WP_39
+ WP_40 WP_41 WP_42 WP_43 WP_44 WP_45 WP_46 WP_47 WP_48 WP_49 WP_50 WP_51 WP_52 WP_53 WP_54 WP_55 WP_56 WP_57 WP_58 WP_59
+ WP_60 WP_61 WP_62 WP_63 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626
+ 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646
+ 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666
+ 667 668 669 670 671 672 673 674
+ ICV_46 $T=0 54400 0 0 $X=-1000 $Y=53400
X2 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_64 WP_65 WP_66 WP_67 WP_68 WP_69 WP_70 WP_71
+ WP_72 WP_73 WP_74 WP_75 WP_76 WP_77 WP_78 WP_79 WP_80 WP_81 WP_82 WP_83 WP_84 WP_85 WP_86 WP_87 WP_88 WP_89 WP_90 WP_91
+ WP_92 WP_93 WP_94 WP_95 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738
+ ICV_46 $T=0 108800 0 0 $X=-1000 $Y=107800
X3 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_96 WP_97 WP_98 WP_99 WP_100 WP_101 WP_102 WP_103
+ WP_104 WP_105 WP_106 WP_107 WP_108 WP_109 WP_110 WP_111 WP_112 WP_113 WP_114 WP_115 WP_116 WP_117 WP_118 WP_119 WP_120 WP_121 WP_122 WP_123
+ WP_124 WP_125 WP_126 WP_127 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754
+ 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774
+ 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794
+ 795 796 797 798 799 800 801 802
+ ICV_46 $T=0 163200 0 0 $X=-1000 $Y=162200
X4 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_128 WP_129 WP_130 WP_131 WP_132 WP_133 WP_134 WP_135
+ WP_136 WP_137 WP_138 WP_139 WP_140 WP_141 WP_142 WP_143 WP_144 WP_145 WP_146 WP_147 WP_148 WP_149 WP_150 WP_151 WP_152 WP_153 WP_154 WP_155
+ WP_156 WP_157 WP_158 WP_159 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866
+ ICV_46 $T=0 217600 0 0 $X=-1000 $Y=216600
X5 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_160 WP_161 WP_162 WP_163 WP_164 WP_165 WP_166 WP_167
+ WP_168 WP_169 WP_170 WP_171 WP_172 WP_173 WP_174 WP_175 WP_176 WP_177 WP_178 WP_179 WP_180 WP_181 WP_182 WP_183 WP_184 WP_185 WP_186 WP_187
+ WP_188 WP_189 WP_190 WP_191 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882
+ 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902
+ 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922
+ 923 924 925 926 927 928 929 930
+ ICV_46 $T=0 272000 0 0 $X=-1000 $Y=271000
X6 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_192 WP_193 WP_194 WP_195 WP_196 WP_197 WP_198 WP_199
+ WP_200 WP_201 WP_202 WP_203 WP_204 WP_205 WP_206 WP_207 WP_208 WP_209 WP_210 WP_211 WP_212 WP_213 WP_214 WP_215 WP_216 WP_217 WP_218 WP_219
+ WP_220 WP_221 WP_222 WP_223 931 932 933 934 935 936 937 938 939 940 941 942 943 944 945 946
+ 947 948 949 950 951 952 953 954 955 956 957 958 959 960 961 962 963 964 965 966
+ 967 968 969 970 971 972 973 974 975 976 977 978 979 980 981 982 983 984 985 986
+ 987 988 989 990 991 992 993 994
+ ICV_46 $T=0 326400 0 0 $X=-1000 $Y=325400
X7 VSS VDD BL__0 BL__1 BL_1 BL_2 BL__2 BL__3 BL_3 BL_4 BL__4 BL__5 BL_5 BL_6 BL__6 BL__7 BL_7 BL_8 BL__8 BL__9
+ BL_9 BL_10 BL__10 BL__11 BL_11 BL_12 BL__12 BL__13 BL_13 BL_14 BL__14 BL__15 WP_224 WP_225 WP_226 WP_227 WP_228 WP_229 WP_230 WP_231
+ WP_232 WP_233 WP_234 WP_235 WP_236 WP_237 WP_238 WP_239 WP_240 WP_241 WP_242 WP_243 WP_244 WP_245 WP_246 WP_247 WP_248 WP_249 WP_250 WP_251
+ WP_252 WP_253 WP_254 WP_255 995 996 997 998 999 1000 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010
+ 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030
+ 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050
+ 1051 1052 1053 1054 1055 1056 1057 1058
+ ICV_46 $T=0 380800 0 0 $X=-1000 $Y=379800
.ENDS
***************************************
.SUBCKT ICV_56 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=1058 FDC=24064
*.SEEDPROM
X0 1 2 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277
+ 278 279 280 281 282 283 284 285 286 287 288 289 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150
+ 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210
+ 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230
+ 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250
+ 251 252 253 254 255 256 257 258 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ SIGN_MEMBIT_COL $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_133 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPEG2
** N=7 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL BLT BL_ BLT_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPOP2
** N=7 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD BL BLT VSS BL_ BLT_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPEP2
** N=7 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD BL BLT BL_ BLT_ VSS
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAPOG2
** N=7 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL BLT BL_ BLT_
.ENDS
***************************************
.SUBCKT SIGN_MEMPCAP_ROWX16
** N=66 EP=0 IP=96 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL_0 BLT_0 BL__0 BLT__0 BL_4 BLT_4 BL__4 BLT__4 BL_8 BLT_8 BL__8 BLT__8 BL_12 BLT_12 BL__12 BLT__12 BL_1 BLT_1
*+ BL__1 BLT__1 BL_5 BLT_5 BL__5 BLT__5 BL_9 BLT_9 BL__9 BLT__9 BL_13 BLT_13 BL__13 BLT__13 BL_2 BLT_2 BL__2 BLT__2 BL_6 BLT_6
*+ BL__6 BLT__6 BL_10 BLT_10 BL__10 BLT__10 BL_14 BLT_14 BL__14 BLT__14 BL_3 BLT_3 BL__3 BLT__3 BL_7 BLT_7 BL__7 BLT__7 BL_11 BLT_11
*+ BL__11 BLT__11 BL_15 BLT_15 BL__15 BLT__15
.ENDS
***************************************
.SUBCKT ICV_58
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_134
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_137 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 310 341 406
+ 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426
+ 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446
+ 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466
+ 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486
+ 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506
+ 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526
+ 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546
+ 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566
+ 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586
+ 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606
+ 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626
+ 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646
+ 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666
+ 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686
+ 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706
+ 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726
+ 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746
+ 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766
+ 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786
+ 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806
+ 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826
+ 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846
+ 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866
+ 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886
+ 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906
+ 907 908 909 910 911 912 913 914 915 916 917
** N=917 EP=791 IP=955 FDC=24680
*.SEEDPROM
X0 2 1 3 4 5 262 263 268 269 270 271 272 273 274 275 276 277 264 265 266
+ 267 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328
+ 329 330 331 332 333 334 335 336 337 338 339 340 341
+ ICV_136 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 311 312
+ 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 406 407 408 409 410 411 412 413 414 415 416 417
+ 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437
+ 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457
+ 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477
+ 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497
+ 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517
+ 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537
+ 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557
+ 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577
+ 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597
+ 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617
+ 618 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637
+ 638 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657
+ 658 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677
+ 678 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697
+ 698 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717
+ 718 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737
+ 738 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757
+ 758 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777
+ 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797
+ 798 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817
+ 818 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837
+ 838 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857
+ 858 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877
+ 878 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897
+ 898 899 900 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917
+ ICV_133 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT SIGN_MEMMUX_CD_EVEN VSS VDD DWSA_5 DRSA_5 DRSA_6 DWSA_6 YP0_0 YP0_1 YP0_2 YP0_3 YP1_0 YP1_1 YP1_2 YP1_3 A0_ A0 GTP BL0_1 BL0__1 BL1_1
+ BL1__1 BL0_3 BL0__3 BL1_3 BL1__3 BL0_5 BL0__5 BL1_5 BL1__5 BL0_7 BL0__7 BL1_7 BL1__7 BL0_0 BL0__0 BL1_0 BL1__0 BL0_2 BL0__2 BL1_2
+ BL1__2 BL0_4 BL0__4 BL1_4 BL1__4 BL0_6 BL0__6 BL1_6 BL1__6
** N=65 EP=49 IP=232 FDC=480
*.CALIBRE ISOLATED NETS: DRSA_1 DWSA_1 DRSA_3 DWSA_3 DRSA_7 DWSA_7 DRSA_0 DWSA_0 DRSA_2 DWSA_2 DRSA_4 DWSA_4 STUBDW STUBDR_ STUBDR STUBDW_
X0 VSS VDD BL0_1 BL0__1 BL1__1 BL1_1 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 YP0_1 VDD SIGN_MEMCD2 $T=4800 0 1 180 $X=1400 $Y=-1000
X1 VSS VDD BL0_3 BL0__3 BL1__3 BL1_3 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 YP0_3 VDD SIGN_MEMCD2 $T=9600 0 1 180 $X=6200 $Y=-1000
X2 VSS VDD BL0_5 BL0__5 BL1__5 BL1_5 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 VDD YP1_1 SIGN_MEMCD2 $T=14400 0 1 180 $X=11000 $Y=-1000
X3 VSS VDD BL0_7 BL0__7 BL1__7 BL1_7 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 VDD YP1_3 SIGN_MEMCD2 $T=19200 0 1 180 $X=15800 $Y=-1000
X4 VSS VDD BL0_0 BL0__0 BL1__0 BL1_0 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 YP0_0 VDD SIGN_MEMCD $T=0 0 0 0 $X=-1000 $Y=-1000
X5 VSS VDD BL0_2 BL0__2 BL1__2 BL1_2 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 YP0_2 VDD SIGN_MEMCD $T=4800 0 0 0 $X=3800 $Y=-1000
X6 VSS VDD BL0_4 BL0__4 BL1__4 BL1_4 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 VDD YP1_0 SIGN_MEMCD $T=9600 0 0 0 $X=8600 $Y=-1000
X7 VSS VDD BL0_6 BL0__6 BL1__6 BL1_6 A0_ A0 GTP DRSA_6 DRSA_5 DWSA_5 DWSA_6 VDD YP1_2 SIGN_MEMCD $T=14400 0 0 0 $X=13400 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_53 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55
** N=62 EP=55 IP=100 FDC=616
X0 1 3 4 SIGN_MEMFCBWM16 $T=0 0 0 270 $X=-1000 $Y=-20200
X1 1 2 60 5 6 61 4 62 9 10 11 3 SIGN_MEMIOX $T=1200 -9600 0 270 $X=200 $Y=-20200
X2 1 9 10 11 SIGN_MEMFLIO $T=1200 0 0 270 $X=200 $Y=-10600
X3 1 2 60 61 7 8 62 12 SIGN_MEMSA8 $T=12470 -9600 0 270 $X=11470 $Y=-20200
X4 1 12 SIGN_MEMFLSA $T=12470 0 0 270 $X=11470 $Y=-10600
X5 1 2 5 7 8 6 22 21 20 19 18 17 16 15 13 14 23 31 30 29
+ 28 39 38 37 36 47 46 45 44 55 54 53 52 24 25 26 27 32 33 34
+ 35 40 41 42 43 48 49 50 51
+ SIGN_MEMMUX_CD_EVEN $T=22810 0 0 270 $X=21810 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_131 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=57 EP=53 IP=59 FDC=616
X0 1 3 4 2 8 11 10 9 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_51
** N=34 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_130
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=1058 FDC=24064
*.SEEDPROM
X0 1 2 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277
+ 278 279 280 281 282 283 284 285 286 287 288 289 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150
+ 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210
+ 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230
+ 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250
+ 251 252 253 254 255 256 257 258 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ SIGN_MEMBIT_COL $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_128 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_49
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_129
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_132 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 314 345 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921
** N=921 EP=791 IP=959 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280
+ 281 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345
+ ICV_131 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 344 343
+ 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326 325 324 323
+ 322 321 320 319 318 317 316 315 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601
+ 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661
+ 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681
+ 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701
+ 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721
+ 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741
+ 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761
+ 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781
+ 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801
+ 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821
+ 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841
+ 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861
+ 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881
+ 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901
+ 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921
+ ICV_128 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCCSTRAP VSS WL NDL NDR
** N=8 EP=4 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: VDD
M0 NDL WL VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=90 $Y=1390 $D=103
M1 NDR WL VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1390 $D=103
.ENDS
***************************************
.SUBCKT ICV_92 1 3 4
** N=6 EP=3 IP=10 FDC=4
X0 1 3 5 6 SIGN_MEMFLCCSTRAP $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 4 5 6 SIGN_MEMFLCCSTRAP $T=0 3400 1 0 $X=-1000 $Y=700
.ENDS
***************************************
.SUBCKT ICV_93 1 3 4 5 6
** N=6 EP=5 IP=8 FDC=8
X0 1 3 4 ICV_92 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 5 6 ICV_92 $T=0 3400 0 0 $X=-1000 $Y=2400
.ENDS
***************************************
.SUBCKT ICV_94 1 3 4 5 6 7 8 9 10
** N=10 EP=9 IP=12 FDC=16
X0 1 3 4 5 6 ICV_93 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 7 8 9 10 ICV_93 $T=0 6800 0 0 $X=-1000 $Y=5800
.ENDS
***************************************
.SUBCKT ICV_95 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=17 IP=20 FDC=32
X0 1 3 4 5 6 7 8 9 10 ICV_94 $T=0 0 0 0 $X=-1000 $Y=-1000
X1 1 11 12 13 14 15 16 17 18 ICV_94 $T=0 13600 0 0 $X=-1000 $Y=12600
.ENDS
***************************************
.SUBCKT ICV_142 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -38400 0 270 $X=62320 $Y=-40600
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -38400 0 270 $X=89520 $Y=-40600
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -38400 0 270 $X=116720 $Y=-40600
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -38400 0 270 $X=143920 $Y=-40600
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -38400 0 270 $X=171120 $Y=-40600
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -38400 0 270 $X=198320 $Y=-40600
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -38400 0 270 $X=225520 $Y=-40600
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -38400 0 270 $X=252720 $Y=-40600
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -38400 0 270 $X=279920 $Y=-40600
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -38400 0 270 $X=307120 $Y=-40600
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -38400 0 270 $X=334320 $Y=-40600
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -38400 0 270 $X=361520 $Y=-40600
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -38400 0 270 $X=388720 $Y=-40600
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -38400 0 270 $X=415920 $Y=-40600
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -38400 0 270 $X=443120 $Y=-40600
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -38400 0 270 $X=470320 $Y=-40600
.ENDS
***************************************
.SUBCKT ICV_126 1 2 3 4 5 6 7 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=63 EP=53 IP=59 FDC=616
X0 1 3 4 2 22 25 24 23 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_125
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_123 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_124
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_127 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 265 267 269 271 272 273 274 275 276 277 278 279 280 281 314 345 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921
** N=921 EP=791 IP=959 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 272 273 274 275 276 277 278 279 280 281 265 267 269
+ 271 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345
+ ICV_126 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 315 316
+ 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336
+ 337 338 339 340 341 342 343 344 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601
+ 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661
+ 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681
+ 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701
+ 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721
+ 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741
+ 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761
+ 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781
+ 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801
+ 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821
+ 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841
+ 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861
+ 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881
+ 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901
+ 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921
+ ICV_123 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_121 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=57 EP=53 IP=59 FDC=616
X0 1 3 4 2 8 11 10 9 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_120
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_118 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_119
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_122 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 314 345 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921
** N=921 EP=791 IP=959 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280
+ 281 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345
+ ICV_121 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 344 343
+ 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326 325 324 323
+ 322 321 320 319 318 317 316 315 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601
+ 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661
+ 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681
+ 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701
+ 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721
+ 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741
+ 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761
+ 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781
+ 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801
+ 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821
+ 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841
+ 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861
+ 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881
+ 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901
+ 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921
+ ICV_118 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_141 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -78000 0 270 $X=62320 $Y=-80200
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -78000 0 270 $X=89520 $Y=-80200
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -78000 0 270 $X=116720 $Y=-80200
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -78000 0 270 $X=143920 $Y=-80200
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -78000 0 270 $X=171120 $Y=-80200
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -78000 0 270 $X=198320 $Y=-80200
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -78000 0 270 $X=225520 $Y=-80200
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -78000 0 270 $X=252720 $Y=-80200
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -78000 0 270 $X=279920 $Y=-80200
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -78000 0 270 $X=307120 $Y=-80200
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -78000 0 270 $X=334320 $Y=-80200
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -78000 0 270 $X=361520 $Y=-80200
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -78000 0 270 $X=388720 $Y=-80200
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -78000 0 270 $X=415920 $Y=-80200
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -78000 0 270 $X=443120 $Y=-80200
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -78000 0 270 $X=470320 $Y=-80200
.ENDS
***************************************
.SUBCKT ICV_116 1 2 3 4 5 6 7 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=63 EP=53 IP=59 FDC=616
X0 1 3 4 2 22 25 24 23 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_115
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_113 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_114
** N=67 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_117 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 282 315 346 411
+ 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431
+ 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451
+ 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471
+ 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491
+ 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511
+ 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531
+ 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551
+ 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571
+ 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591
+ 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611
+ 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631
+ 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651
+ 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670 671
+ 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691
+ 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710 711
+ 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730 731
+ 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750 751
+ 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771
+ 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791
+ 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810 811
+ 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830 831
+ 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850 851
+ 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870 871
+ 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890 891
+ 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910 911
+ 912 913 914 915 916 917 918 919 920 921 922
** N=922 EP=791 IP=960 FDC=24680
*.SEEDPROM
X0 4 1 2 3 262 263 264 273 274 275 276 277 278 279 280 281 282 266 268 270
+ 272 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333
+ 334 335 336 337 338 339 340 341 342 343 344 345 346
+ ICV_116 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 316 317
+ 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337
+ 338 339 340 341 342 343 344 345 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822
+ 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842
+ 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862
+ 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882
+ 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902
+ 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922
+ ICV_113 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_111 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=57 EP=53 IP=59 FDC=616
X0 1 3 4 2 8 11 10 9 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_110
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_108 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_109
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_112 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 314 345 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921
** N=921 EP=791 IP=959 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280
+ 281 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345
+ ICV_111 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 344 343
+ 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326 325 324 323
+ 322 321 320 319 318 317 316 315 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601
+ 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661
+ 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681
+ 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701
+ 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721
+ 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741
+ 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761
+ 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781
+ 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801
+ 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821
+ 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841
+ 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861
+ 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881
+ 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901
+ 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921
+ ICV_108 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_140 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -117600 0 270 $X=62320 $Y=-119800
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -117600 0 270 $X=89520 $Y=-119800
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -117600 0 270 $X=116720 $Y=-119800
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -117600 0 270 $X=143920 $Y=-119800
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -117600 0 270 $X=171120 $Y=-119800
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -117600 0 270 $X=198320 $Y=-119800
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -117600 0 270 $X=225520 $Y=-119800
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -117600 0 270 $X=252720 $Y=-119800
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -117600 0 270 $X=279920 $Y=-119800
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -117600 0 270 $X=307120 $Y=-119800
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -117600 0 270 $X=334320 $Y=-119800
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -117600 0 270 $X=361520 $Y=-119800
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -117600 0 270 $X=388720 $Y=-119800
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -117600 0 270 $X=415920 $Y=-119800
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -117600 0 270 $X=443120 $Y=-119800
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -117600 0 270 $X=470320 $Y=-119800
.ENDS
***************************************
.SUBCKT ICV_106 1 2 3 4 5 6 7 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57
** N=63 EP=53 IP=59 FDC=616
X0 1 3 4 2 22 25 24 23 5 6 7 6 13 12 14 15 16 17 18 19
+ 20 21 6 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43 42 41
+ 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_105
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_103 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_104
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_107 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 265 267 269 271 272 273 274 275 276 277 278 279 280 281 314 345 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921
** N=921 EP=791 IP=959 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 272 273 274 275 276 277 278 279 280 281 265 267 269
+ 271 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345
+ ICV_106 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 315 316
+ 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336
+ 337 338 339 340 341 342 343 344 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601
+ 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641
+ 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661
+ 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681
+ 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701
+ 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721
+ 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741
+ 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761
+ 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781
+ 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801
+ 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821
+ 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841
+ 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861
+ 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881
+ 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901
+ 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921
+ ICV_103 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_139 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53
** N=68 EP=53 IP=95 FDC=617
D0 1 1 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=140 $Y=-146660 $D=558
D1 1 3 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=140 $Y=-141760 $D=558
D2 1 4 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=140 $Y=-139360 $D=558
X3 1 2 58 5 6 59 4 60 20 19 21 3 SIGN_MEMIOX $T=1200 -147600 1 90 $X=200 $Y=-148600
X4 1 20 19 21 SIGN_MEMFLIO $T=1200 -157200 1 90 $X=200 $Y=-158200
X5 1 2 58 59 7 8 60 19 SIGN_MEMSA8 $T=12470 -147600 1 90 $X=11470 $Y=-148600
X6 1 19 SIGN_MEMFLSA $T=12470 -157200 1 90 $X=11470 $Y=-158200
X7 1 2 5 7 8 6 18 17 16 15 14 13 12 11 10 9 19 29 28 27
+ 26 37 36 35 34 45 44 43 42 53 52 51 50 22 23 24 25 30 31 32
+ 33 38 39 40 41 46 47 48 49
+ SIGN_MEMMUX_CD_EVEN $T=22810 -157200 1 90 $X=21810 $Y=-158200
.ENDS
***************************************
.SUBCKT ICV_138 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 387 388 389 390 391 392 393 394 395 396 397 398
+ 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418
+ 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438
+ 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458
+ 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478
+ 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498
+ 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518
+ 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538
+ 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558
+ 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578
+ 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598
+ 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618
+ 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658
+ 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678
+ 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
+ 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718
+ 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738
+ 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758
+ 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778
+ 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798
+ 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878
+ 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898
** N=898 EP=800 IP=1158 FDC=24064
*.SEEDPROM
X1 1 2 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277
+ 278 279 280 281 282 283 284 285 286 287 288 289 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150
+ 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210
+ 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230
+ 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250
+ 251 252 253 254 255 256 257 258 387 388 389 390 391 392 393 394 395 396 397 398
+ 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418
+ 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438
+ 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458
+ 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478
+ 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498
+ 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518
+ 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538
+ 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558
+ 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578
+ 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598
+ 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618
+ 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658
+ 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678
+ 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
+ 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718
+ 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738
+ 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758
+ 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778
+ 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798
+ 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878
+ 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898
+ SIGN_MEMBIT_COL $T=63320 -157200 1 90 $X=62320 $Y=-158200
.ENDS
***************************************
.SUBCKT SIGN_MEMWING_8_LEFT VDD VSS D_0 Q_0 D_1 Q_1 D_2 Q_2 D_3 Q_3 D_4 Q_4 D_5 Q_5 D_6 Q_6 D_7 Q_7 GTP_0 WL_0
+ WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 WL_20
+ WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40
+ WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 WL_59 WL_60
+ WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80
+ WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98 WL_99 WL_100
+ WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 WL_119 WL_120
+ WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138 WL_139 WL_140
+ WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158 WL_159 WL_160
+ WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178 WL_179 WL_180
+ WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198 WL_199 WL_200
+ WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218 WL_219 WL_220
+ WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238 WL_239 WL_240
+ WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255 WE OE_ A0 A0_ YP1_3
+ YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 577 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680
+ 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700
+ 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740
+ 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760
+ 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780
+ 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800
+ 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820
+ 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840
+ 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860
+ 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880
+ 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900
+ 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920
+ 921 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 938 939 940
+ 941 942 943 944 945 946 947 948 949 950 951 952 953 954 955 956 957 958 959 960
+ 961 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980
+ 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 1000
+ 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020
+ 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040
+ 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060
+ 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080
+ 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
+ 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120
+ 1121
** N=4718 EP=801 IP=7451 FDC=202561
*.SEEDPROM
*.CALIBRE ISOLATED NETS: BLT__0 BLT_0 BLT__1 BLT_1 BLT__2 BLT_2 BLT__3 BLT_3 BLT__4 BLT_4 BLT__5 BLT_5 BLT__6 BLT_6 BLT__7 BLT_7 BLT__8 BLT_8 BLT__9 BLT_9
*+ BLT__10 BLT_10 BLT__11 BLT_11 BLT__12 BLT_12 BLT__13 BLT_13 BLT__14 BLT_14 BLT__15 BLT_15 BLT_31 BLT__31 BLT_30 BLT__30 BLT_29 BLT__29 BLT_28 BLT__28
*+ BLT_27 BLT__27 BLT_26 BLT__26 BLT_25 BLT__25 BLT_24 BLT__24 BLT_23 BLT__23 BLT_22 BLT__22 BLT_21 BLT__21 BLT_20 BLT__20 BLT_19 BLT__19 BLT_18 BLT__18
*+ BLT_17 BLT__17 BLT_16 BLT__16 BLT__32 BLT_32 BLT__33 BLT_33 BLT__34 BLT_34 BLT__35 BLT_35 BLT__36 BLT_36 BLT__37 BLT_37 BLT__38 BLT_38 BLT__39 BLT_39
*+ BLT__40 BLT_40 BLT__41 BLT_41 BLT__42 BLT_42 BLT__43 BLT_43 BLT__44 BLT_44 BLT__45 BLT_45 BLT__46 BLT_46 BLT__47 BLT_47 BLT_63 BLT__63 BLT_62 BLT__62
*+ BLT_61 BLT__61 BLT_60 BLT__60 BLT_59 BLT__59 BLT_58 BLT__58 BLT_57 BLT__57 BLT_56 BLT__56 BLT_55 BLT__55 BLT_54 BLT__54 BLT_53 BLT__53 BLT_52 BLT__52
*+ BLT_51 BLT__51 BLT_50 BLT__50 BLT_49 BLT__49 BLT_48 BLT__48 BLT__64 BLT_64 BLT__65 BLT_65 BLT__66 BLT_66 BLT__67 BLT_67 BLT__68 BLT_68 BLT__69 BLT_69
*+ BLT__70 BLT_70 BLT__71 BLT_71 BLT__72 BLT_72 BLT__73 BLT_73 BLT__74 BLT_74 BLT__75 BLT_75 BLT__76 BLT_76 BLT__77 BLT_77 BLT__78 BLT_78 BLT__79 BLT_79
*+ BLT_95 BLT__95 BLT_94 BLT__94 BLT_93 BLT__93 BLT_92 BLT__92 BLT_91 BLT__91 BLT_90 BLT__90 BLT_89 BLT__89 BLT_88 BLT__88 BLT_87 BLT__87 BLT_86 BLT__86
*+ BLT_85 BLT__85 BLT_84 BLT__84 BLT_83 BLT__83 BLT_82 BLT__82 BLT_81 BLT__81 BLT_80 BLT__80 BLT__96 BLT_96 BLT__97 BLT_97 BLT__98 BLT_98 BLT__99 BLT_99
*+ BLT__100 BLT_100 BLT__101 BLT_101 BLT__102 BLT_102 BLT__103 BLT_103 BLT__104 BLT_104 BLT__105 BLT_105 BLT__106 BLT_106 BLT__107 BLT_107 BLT__108 BLT_108 BLT__109 BLT_109
*+ BLT__110 BLT_110 BLT__111 BLT_111 BLT_127 BLT__127 BLT_126 BLT__126 BLT_125 BLT__125 BLT_124 BLT__124 BLT_123 BLT__123 BLT_122 BLT__122 BLT_121 BLT__121 BLT_120 BLT__120
*+ BLT_119 BLT__119 BLT_118 BLT__118 BLT_117 BLT__117 BLT_116 BLT__116 BLT_115 BLT__115 BLT_114 BLT__114 BLT_113 BLT__113 BLT_112 BLT__112
M0 1122 WL_0 1123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=64710 $D=103
M1 1124 WL_1 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=65200 $D=103
M2 1122 WL_2 1125 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=68110 $D=103
M3 1126 WL_3 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=68600 $D=103
M4 1122 WL_4 1127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=71510 $D=103
M5 1128 WL_5 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=72000 $D=103
M6 1122 WL_6 1129 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=74910 $D=103
M7 1130 WL_7 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=75400 $D=103
M8 1122 WL_8 1131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=78310 $D=103
M9 1132 WL_9 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=78800 $D=103
M10 1122 WL_10 1133 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=81710 $D=103
M11 1134 WL_11 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=82200 $D=103
M12 1122 WL_12 1135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=85110 $D=103
M13 1136 WL_13 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=85600 $D=103
M14 1122 WL_14 1137 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=88510 $D=103
M15 1138 WL_15 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=89000 $D=103
M16 1122 WL_16 1139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=91910 $D=103
M17 1140 WL_17 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=92400 $D=103
M18 1122 WL_18 1141 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=95310 $D=103
M19 1142 WL_19 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=95800 $D=103
M20 1122 WL_20 1143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=98710 $D=103
M21 1144 WL_21 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=99200 $D=103
M22 1122 WL_22 1145 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=102110 $D=103
M23 1146 WL_23 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=102600 $D=103
M24 1122 WL_24 1147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=105510 $D=103
M25 1148 WL_25 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=106000 $D=103
M26 1122 WL_26 1149 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=108910 $D=103
M27 1150 WL_27 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=109400 $D=103
M28 1122 WL_28 1151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=112310 $D=103
M29 1152 WL_29 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=112800 $D=103
M30 1122 WL_30 1153 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=115710 $D=103
M31 1154 WL_31 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=116200 $D=103
M32 1122 WL_32 1155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=119110 $D=103
M33 1156 WL_33 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=119600 $D=103
M34 1122 WL_34 1157 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=122510 $D=103
M35 1158 WL_35 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=123000 $D=103
M36 1122 WL_36 1159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=125910 $D=103
M37 1160 WL_37 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=126400 $D=103
M38 1122 WL_38 1161 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=129310 $D=103
M39 1162 WL_39 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=129800 $D=103
M40 1122 WL_40 1163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=132710 $D=103
M41 1164 WL_41 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=133200 $D=103
M42 1122 WL_42 1165 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=136110 $D=103
M43 1166 WL_43 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=136600 $D=103
M44 1122 WL_44 1167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=139510 $D=103
M45 1168 WL_45 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=140000 $D=103
M46 1122 WL_46 1169 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=142910 $D=103
M47 1170 WL_47 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=143400 $D=103
M48 1122 WL_48 1171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=146310 $D=103
M49 1172 WL_49 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=146800 $D=103
M50 1122 WL_50 1173 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=149710 $D=103
M51 1174 WL_51 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=150200 $D=103
M52 1122 WL_52 1175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=153110 $D=103
M53 1176 WL_53 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=153600 $D=103
M54 1122 WL_54 1177 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=156510 $D=103
M55 1178 WL_55 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=157000 $D=103
M56 1122 WL_56 1179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=159910 $D=103
M57 1180 WL_57 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=160400 $D=103
M58 1122 WL_58 1181 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=163310 $D=103
M59 1182 WL_59 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=163800 $D=103
M60 1122 WL_60 1183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=166710 $D=103
M61 1184 WL_61 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=167200 $D=103
M62 1122 WL_62 1185 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=170110 $D=103
M63 1186 WL_63 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=170600 $D=103
M64 1122 WL_64 1187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=173510 $D=103
M65 1188 WL_65 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=174000 $D=103
M66 1122 WL_66 1189 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=176910 $D=103
M67 1190 WL_67 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=177400 $D=103
M68 1122 WL_68 1191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=180310 $D=103
M69 1192 WL_69 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=180800 $D=103
M70 1122 WL_70 1193 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=183710 $D=103
M71 1194 WL_71 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=184200 $D=103
M72 1122 WL_72 1195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=187110 $D=103
M73 1196 WL_73 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=187600 $D=103
M74 1122 WL_74 1197 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=190510 $D=103
M75 1198 WL_75 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=191000 $D=103
M76 1122 WL_76 1199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=193910 $D=103
M77 1200 WL_77 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=194400 $D=103
M78 1122 WL_78 1201 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=197310 $D=103
M79 1202 WL_79 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=197800 $D=103
M80 1122 WL_80 1203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=200710 $D=103
M81 1204 WL_81 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=201200 $D=103
M82 1122 WL_82 1205 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=204110 $D=103
M83 1206 WL_83 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=204600 $D=103
M84 1122 WL_84 1207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=207510 $D=103
M85 1208 WL_85 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=208000 $D=103
M86 1122 WL_86 1209 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=210910 $D=103
M87 1210 WL_87 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=211400 $D=103
M88 1122 WL_88 1211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=214310 $D=103
M89 1212 WL_89 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=214800 $D=103
M90 1122 WL_90 1213 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=217710 $D=103
M91 1214 WL_91 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=218200 $D=103
M92 1122 WL_92 1215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=221110 $D=103
M93 1216 WL_93 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=221600 $D=103
M94 1122 WL_94 1217 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=224510 $D=103
M95 1218 WL_95 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=225000 $D=103
M96 1122 WL_96 1219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=227910 $D=103
M97 1220 WL_97 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=228400 $D=103
M98 1122 WL_98 1221 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=231310 $D=103
M99 1222 WL_99 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=231800 $D=103
M100 1122 WL_100 1223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=234710 $D=103
M101 1224 WL_101 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=235200 $D=103
M102 1122 WL_102 1225 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=238110 $D=103
M103 1226 WL_103 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=238600 $D=103
M104 1122 WL_104 1227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=241510 $D=103
M105 1228 WL_105 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=242000 $D=103
M106 1122 WL_106 1229 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=244910 $D=103
M107 1230 WL_107 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=245400 $D=103
M108 1122 WL_108 1231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=248310 $D=103
M109 1232 WL_109 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=248800 $D=103
M110 1122 WL_110 1233 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=251710 $D=103
M111 1234 WL_111 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=252200 $D=103
M112 1122 WL_112 1235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=255110 $D=103
M113 1236 WL_113 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=255600 $D=103
M114 1122 WL_114 1237 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=258510 $D=103
M115 1238 WL_115 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=259000 $D=103
M116 1122 WL_116 1239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=261910 $D=103
M117 1240 WL_117 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=262400 $D=103
M118 1122 WL_118 1241 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=265310 $D=103
M119 1242 WL_119 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=265800 $D=103
M120 1122 WL_120 1243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=268710 $D=103
M121 1244 WL_121 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=269200 $D=103
M122 1122 WL_122 1245 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=272110 $D=103
M123 1246 WL_123 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=272600 $D=103
M124 1122 WL_124 1247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=275510 $D=103
M125 1248 WL_125 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=276000 $D=103
M126 1122 WL_126 1249 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=278910 $D=103
M127 1250 WL_127 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=279400 $D=103
M128 1122 WL_128 1251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=282310 $D=103
M129 1252 WL_129 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=282800 $D=103
M130 1122 WL_130 1253 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=285710 $D=103
M131 1254 WL_131 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=286200 $D=103
M132 1122 WL_132 1255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=289110 $D=103
M133 1256 WL_133 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=289600 $D=103
M134 1122 WL_134 1257 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=292510 $D=103
M135 1258 WL_135 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=293000 $D=103
M136 1122 WL_136 1259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=295910 $D=103
M137 1260 WL_137 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=296400 $D=103
M138 1122 WL_138 1261 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=299310 $D=103
M139 1262 WL_139 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=299800 $D=103
M140 1122 WL_140 1263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=302710 $D=103
M141 1264 WL_141 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=303200 $D=103
M142 1122 WL_142 1265 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=306110 $D=103
M143 1266 WL_143 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=306600 $D=103
M144 1122 WL_144 1267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=309510 $D=103
M145 1268 WL_145 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=310000 $D=103
M146 1122 WL_146 1269 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=312910 $D=103
M147 1270 WL_147 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=313400 $D=103
M148 1122 WL_148 1271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=316310 $D=103
M149 1272 WL_149 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=316800 $D=103
M150 1122 WL_150 1273 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=319710 $D=103
M151 1274 WL_151 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=320200 $D=103
M152 1122 WL_152 1275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=323110 $D=103
M153 1276 WL_153 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=323600 $D=103
M154 1122 WL_154 1277 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=326510 $D=103
M155 1278 WL_155 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=327000 $D=103
M156 1122 WL_156 1279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=329910 $D=103
M157 1280 WL_157 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=330400 $D=103
M158 1122 WL_158 1281 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=333310 $D=103
M159 1282 WL_159 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=333800 $D=103
M160 1122 WL_160 1283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=336710 $D=103
M161 1284 WL_161 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=337200 $D=103
M162 1122 WL_162 1285 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=340110 $D=103
M163 1286 WL_163 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=340600 $D=103
M164 1122 WL_164 1287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=343510 $D=103
M165 1288 WL_165 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=344000 $D=103
M166 1122 WL_166 1289 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=346910 $D=103
M167 1290 WL_167 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=347400 $D=103
M168 1122 WL_168 1291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=350310 $D=103
M169 1292 WL_169 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=350800 $D=103
M170 1122 WL_170 1293 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=353710 $D=103
M171 1294 WL_171 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=354200 $D=103
M172 1122 WL_172 1295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=357110 $D=103
M173 1296 WL_173 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=357600 $D=103
M174 1122 WL_174 1297 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=360510 $D=103
M175 1298 WL_175 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=361000 $D=103
M176 1122 WL_176 1299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=363910 $D=103
M177 1300 WL_177 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=364400 $D=103
M178 1122 WL_178 1301 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=367310 $D=103
M179 1302 WL_179 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=367800 $D=103
M180 1122 WL_180 1303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=370710 $D=103
M181 1304 WL_181 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=371200 $D=103
M182 1122 WL_182 1305 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=374110 $D=103
M183 1306 WL_183 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=374600 $D=103
M184 1122 WL_184 1307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=377510 $D=103
M185 1308 WL_185 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=378000 $D=103
M186 1122 WL_186 1309 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=380910 $D=103
M187 1310 WL_187 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=381400 $D=103
M188 1122 WL_188 1311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=384310 $D=103
M189 1312 WL_189 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=384800 $D=103
M190 1122 WL_190 1313 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=387710 $D=103
M191 1314 WL_191 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=388200 $D=103
M192 1122 WL_192 1315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=391110 $D=103
M193 1316 WL_193 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=391600 $D=103
M194 1122 WL_194 1317 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=394510 $D=103
M195 1318 WL_195 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=395000 $D=103
M196 1122 WL_196 1319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=397910 $D=103
M197 1320 WL_197 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=398400 $D=103
M198 1122 WL_198 1321 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=401310 $D=103
M199 1322 WL_199 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=401800 $D=103
M200 1122 WL_200 1323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=404710 $D=103
M201 1324 WL_201 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=405200 $D=103
M202 1122 WL_202 1325 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=408110 $D=103
M203 1326 WL_203 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=408600 $D=103
M204 1122 WL_204 1327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=411510 $D=103
M205 1328 WL_205 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=412000 $D=103
M206 1122 WL_206 1329 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=414910 $D=103
M207 1330 WL_207 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=415400 $D=103
M208 1122 WL_208 1331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=418310 $D=103
M209 1332 WL_209 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=418800 $D=103
M210 1122 WL_210 1333 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=421710 $D=103
M211 1334 WL_211 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=422200 $D=103
M212 1122 WL_212 1335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=425110 $D=103
M213 1336 WL_213 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=425600 $D=103
M214 1122 WL_214 1337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=428510 $D=103
M215 1338 WL_215 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=429000 $D=103
M216 1122 WL_216 1339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=431910 $D=103
M217 1340 WL_217 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=432400 $D=103
M218 1122 WL_218 1341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=435310 $D=103
M219 1342 WL_219 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=435800 $D=103
M220 1122 WL_220 1343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=438710 $D=103
M221 1344 WL_221 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=439200 $D=103
M222 1122 WL_222 1345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=442110 $D=103
M223 1346 WL_223 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=442600 $D=103
M224 1122 WL_224 1347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=445510 $D=103
M225 1348 WL_225 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=446000 $D=103
M226 1122 WL_226 1349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=448910 $D=103
M227 1350 WL_227 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=449400 $D=103
M228 1122 WL_228 1351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=452310 $D=103
M229 1352 WL_229 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=452800 $D=103
M230 1122 WL_230 1353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=455710 $D=103
M231 1354 WL_231 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=456200 $D=103
M232 1122 WL_232 1355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=459110 $D=103
M233 1356 WL_233 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=459600 $D=103
M234 1122 WL_234 1357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=462510 $D=103
M235 1358 WL_235 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=463000 $D=103
M236 1122 WL_236 1359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=465910 $D=103
M237 1360 WL_237 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=466400 $D=103
M238 1122 WL_238 1361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=469310 $D=103
M239 1362 WL_239 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=469800 $D=103
M240 1122 WL_240 1363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=472710 $D=103
M241 1364 WL_241 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=473200 $D=103
M242 1122 WL_242 1365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=476110 $D=103
M243 1366 WL_243 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=476600 $D=103
M244 1122 WL_244 1367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=479510 $D=103
M245 1368 WL_245 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=480000 $D=103
M246 1122 WL_246 1369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=482910 $D=103
M247 1370 WL_247 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=483400 $D=103
M248 1122 WL_248 1371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=486310 $D=103
M249 1372 WL_249 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=486800 $D=103
M250 1122 WL_250 1373 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=489710 $D=103
M251 1374 WL_251 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=490200 $D=103
M252 1122 WL_252 1375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=493110 $D=103
M253 1376 WL_253 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=493600 $D=103
M254 1122 WL_254 1377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=496510 $D=103
M255 1378 WL_255 1122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=497000 $D=103
M256 1379 WL_0 1382 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=64710 $D=103
M257 1384 WL_1 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=65200 $D=103
M258 1379 WL_2 1386 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=68110 $D=103
M259 1388 WL_3 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=68600 $D=103
M260 1379 WL_4 1390 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=71510 $D=103
M261 1392 WL_5 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=72000 $D=103
M262 1379 WL_6 1394 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=74910 $D=103
M263 1396 WL_7 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=75400 $D=103
M264 1379 WL_8 1398 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=78310 $D=103
M265 1400 WL_9 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=78800 $D=103
M266 1379 WL_10 1402 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=81710 $D=103
M267 1404 WL_11 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=82200 $D=103
M268 1379 WL_12 1406 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=85110 $D=103
M269 1408 WL_13 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=85600 $D=103
M270 1379 WL_14 1410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=88510 $D=103
M271 1412 WL_15 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=89000 $D=103
M272 1379 WL_16 1414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=91910 $D=103
M273 1416 WL_17 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=92400 $D=103
M274 1379 WL_18 1418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=95310 $D=103
M275 1420 WL_19 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=95800 $D=103
M276 1379 WL_20 1422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=98710 $D=103
M277 1424 WL_21 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=99200 $D=103
M278 1379 WL_22 1426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=102110 $D=103
M279 1428 WL_23 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=102600 $D=103
M280 1379 WL_24 1430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=105510 $D=103
M281 1432 WL_25 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=106000 $D=103
M282 1379 WL_26 1434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=108910 $D=103
M283 1436 WL_27 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=109400 $D=103
M284 1379 WL_28 1438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=112310 $D=103
M285 1440 WL_29 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=112800 $D=103
M286 1379 WL_30 1442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=115710 $D=103
M287 1444 WL_31 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=116200 $D=103
M288 1379 WL_32 1446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=119110 $D=103
M289 1448 WL_33 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=119600 $D=103
M290 1379 WL_34 1450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=122510 $D=103
M291 1452 WL_35 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=123000 $D=103
M292 1379 WL_36 1454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=125910 $D=103
M293 1456 WL_37 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=126400 $D=103
M294 1379 WL_38 1458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=129310 $D=103
M295 1460 WL_39 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=129800 $D=103
M296 1379 WL_40 1462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=132710 $D=103
M297 1464 WL_41 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=133200 $D=103
M298 1379 WL_42 1466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=136110 $D=103
M299 1468 WL_43 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=136600 $D=103
M300 1379 WL_44 1470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=139510 $D=103
M301 1472 WL_45 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=140000 $D=103
M302 1379 WL_46 1474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=142910 $D=103
M303 1476 WL_47 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=143400 $D=103
M304 1379 WL_48 1478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=146310 $D=103
M305 1480 WL_49 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=146800 $D=103
M306 1379 WL_50 1482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=149710 $D=103
M307 1484 WL_51 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=150200 $D=103
M308 1379 WL_52 1486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=153110 $D=103
M309 1488 WL_53 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=153600 $D=103
M310 1379 WL_54 1490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=156510 $D=103
M311 1492 WL_55 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=157000 $D=103
M312 1379 WL_56 1494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=159910 $D=103
M313 1496 WL_57 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=160400 $D=103
M314 1379 WL_58 1498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=163310 $D=103
M315 1500 WL_59 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=163800 $D=103
M316 1379 WL_60 1502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=166710 $D=103
M317 1504 WL_61 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=167200 $D=103
M318 1379 WL_62 1506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=170110 $D=103
M319 1508 WL_63 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=170600 $D=103
M320 1379 WL_64 1510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=173510 $D=103
M321 1512 WL_65 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=174000 $D=103
M322 1379 WL_66 1514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=176910 $D=103
M323 1516 WL_67 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=177400 $D=103
M324 1379 WL_68 1518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=180310 $D=103
M325 1520 WL_69 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=180800 $D=103
M326 1379 WL_70 1522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=183710 $D=103
M327 1524 WL_71 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=184200 $D=103
M328 1379 WL_72 1526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=187110 $D=103
M329 1528 WL_73 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=187600 $D=103
M330 1379 WL_74 1530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=190510 $D=103
M331 1532 WL_75 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=191000 $D=103
M332 1379 WL_76 1534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=193910 $D=103
M333 1536 WL_77 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=194400 $D=103
M334 1379 WL_78 1538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=197310 $D=103
M335 1540 WL_79 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=197800 $D=103
M336 1379 WL_80 1542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=200710 $D=103
M337 1544 WL_81 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=201200 $D=103
M338 1379 WL_82 1546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=204110 $D=103
M339 1548 WL_83 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=204600 $D=103
M340 1379 WL_84 1550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=207510 $D=103
M341 1552 WL_85 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=208000 $D=103
M342 1379 WL_86 1554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=210910 $D=103
M343 1556 WL_87 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=211400 $D=103
M344 1379 WL_88 1558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=214310 $D=103
M345 1560 WL_89 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=214800 $D=103
M346 1379 WL_90 1562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=217710 $D=103
M347 1564 WL_91 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=218200 $D=103
M348 1379 WL_92 1566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=221110 $D=103
M349 1568 WL_93 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=221600 $D=103
M350 1379 WL_94 1570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=224510 $D=103
M351 1572 WL_95 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=225000 $D=103
M352 1379 WL_96 1574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=227910 $D=103
M353 1576 WL_97 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=228400 $D=103
M354 1379 WL_98 1578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=231310 $D=103
M355 1580 WL_99 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=231800 $D=103
M356 1379 WL_100 1582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=234710 $D=103
M357 1584 WL_101 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=235200 $D=103
M358 1379 WL_102 1586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=238110 $D=103
M359 1588 WL_103 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=238600 $D=103
M360 1379 WL_104 1590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=241510 $D=103
M361 1592 WL_105 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=242000 $D=103
M362 1379 WL_106 1594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=244910 $D=103
M363 1596 WL_107 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=245400 $D=103
M364 1379 WL_108 1598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=248310 $D=103
M365 1600 WL_109 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=248800 $D=103
M366 1379 WL_110 1602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=251710 $D=103
M367 1604 WL_111 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=252200 $D=103
M368 1379 WL_112 1606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=255110 $D=103
M369 1608 WL_113 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=255600 $D=103
M370 1379 WL_114 1610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=258510 $D=103
M371 1612 WL_115 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=259000 $D=103
M372 1379 WL_116 1614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=261910 $D=103
M373 1616 WL_117 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=262400 $D=103
M374 1379 WL_118 1618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=265310 $D=103
M375 1620 WL_119 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=265800 $D=103
M376 1379 WL_120 1622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=268710 $D=103
M377 1624 WL_121 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=269200 $D=103
M378 1379 WL_122 1626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=272110 $D=103
M379 1628 WL_123 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=272600 $D=103
M380 1379 WL_124 1630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=275510 $D=103
M381 1632 WL_125 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=276000 $D=103
M382 1379 WL_126 1634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=278910 $D=103
M383 1636 WL_127 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=279400 $D=103
M384 1379 WL_128 1638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=282310 $D=103
M385 1640 WL_129 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=282800 $D=103
M386 1379 WL_130 1642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=285710 $D=103
M387 1644 WL_131 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=286200 $D=103
M388 1379 WL_132 1646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=289110 $D=103
M389 1648 WL_133 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=289600 $D=103
M390 1379 WL_134 1650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=292510 $D=103
M391 1652 WL_135 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=293000 $D=103
M392 1379 WL_136 1654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=295910 $D=103
M393 1656 WL_137 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=296400 $D=103
M394 1379 WL_138 1658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=299310 $D=103
M395 1660 WL_139 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=299800 $D=103
M396 1379 WL_140 1662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=302710 $D=103
M397 1664 WL_141 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=303200 $D=103
M398 1379 WL_142 1666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=306110 $D=103
M399 1668 WL_143 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=306600 $D=103
M400 1379 WL_144 1670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=309510 $D=103
M401 1672 WL_145 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=310000 $D=103
M402 1379 WL_146 1674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=312910 $D=103
M403 1676 WL_147 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=313400 $D=103
M404 1379 WL_148 1678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=316310 $D=103
M405 1680 WL_149 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=316800 $D=103
M406 1379 WL_150 1682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=319710 $D=103
M407 1684 WL_151 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=320200 $D=103
M408 1379 WL_152 1686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=323110 $D=103
M409 1688 WL_153 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=323600 $D=103
M410 1379 WL_154 1690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=326510 $D=103
M411 1692 WL_155 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=327000 $D=103
M412 1379 WL_156 1694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=329910 $D=103
M413 1696 WL_157 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=330400 $D=103
M414 1379 WL_158 1698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=333310 $D=103
M415 1700 WL_159 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=333800 $D=103
M416 1379 WL_160 1702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=336710 $D=103
M417 1704 WL_161 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=337200 $D=103
M418 1379 WL_162 1706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=340110 $D=103
M419 1708 WL_163 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=340600 $D=103
M420 1379 WL_164 1710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=343510 $D=103
M421 1712 WL_165 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=344000 $D=103
M422 1379 WL_166 1714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=346910 $D=103
M423 1716 WL_167 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=347400 $D=103
M424 1379 WL_168 1718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=350310 $D=103
M425 1720 WL_169 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=350800 $D=103
M426 1379 WL_170 1722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=353710 $D=103
M427 1724 WL_171 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=354200 $D=103
M428 1379 WL_172 1726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=357110 $D=103
M429 1728 WL_173 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=357600 $D=103
M430 1379 WL_174 1730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=360510 $D=103
M431 1732 WL_175 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=361000 $D=103
M432 1379 WL_176 1734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=363910 $D=103
M433 1736 WL_177 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=364400 $D=103
M434 1379 WL_178 1738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=367310 $D=103
M435 1740 WL_179 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=367800 $D=103
M436 1379 WL_180 1742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=370710 $D=103
M437 1744 WL_181 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=371200 $D=103
M438 1379 WL_182 1746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=374110 $D=103
M439 1748 WL_183 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=374600 $D=103
M440 1379 WL_184 1750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=377510 $D=103
M441 1752 WL_185 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=378000 $D=103
M442 1379 WL_186 1754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=380910 $D=103
M443 1756 WL_187 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=381400 $D=103
M444 1379 WL_188 1758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=384310 $D=103
M445 1760 WL_189 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=384800 $D=103
M446 1379 WL_190 1762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=387710 $D=103
M447 1764 WL_191 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=388200 $D=103
M448 1379 WL_192 1766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=391110 $D=103
M449 1768 WL_193 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=391600 $D=103
M450 1379 WL_194 1770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=394510 $D=103
M451 1772 WL_195 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=395000 $D=103
M452 1379 WL_196 1774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=397910 $D=103
M453 1776 WL_197 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=398400 $D=103
M454 1379 WL_198 1778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=401310 $D=103
M455 1780 WL_199 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=401800 $D=103
M456 1379 WL_200 1782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=404710 $D=103
M457 1784 WL_201 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=405200 $D=103
M458 1379 WL_202 1786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=408110 $D=103
M459 1788 WL_203 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=408600 $D=103
M460 1379 WL_204 1790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=411510 $D=103
M461 1792 WL_205 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=412000 $D=103
M462 1379 WL_206 1794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=414910 $D=103
M463 1796 WL_207 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=415400 $D=103
M464 1379 WL_208 1798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=418310 $D=103
M465 1800 WL_209 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=418800 $D=103
M466 1379 WL_210 1802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=421710 $D=103
M467 1804 WL_211 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=422200 $D=103
M468 1379 WL_212 1806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=425110 $D=103
M469 1808 WL_213 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=425600 $D=103
M470 1379 WL_214 1810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=428510 $D=103
M471 1812 WL_215 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=429000 $D=103
M472 1379 WL_216 1814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=431910 $D=103
M473 1816 WL_217 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=432400 $D=103
M474 1379 WL_218 1818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=435310 $D=103
M475 1820 WL_219 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=435800 $D=103
M476 1379 WL_220 1822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=438710 $D=103
M477 1824 WL_221 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=439200 $D=103
M478 1379 WL_222 1826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=442110 $D=103
M479 1828 WL_223 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=442600 $D=103
M480 1379 WL_224 1830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=445510 $D=103
M481 1832 WL_225 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=446000 $D=103
M482 1379 WL_226 1834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=448910 $D=103
M483 1836 WL_227 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=449400 $D=103
M484 1379 WL_228 1838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=452310 $D=103
M485 1840 WL_229 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=452800 $D=103
M486 1379 WL_230 1842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=455710 $D=103
M487 1844 WL_231 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=456200 $D=103
M488 1379 WL_232 1846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=459110 $D=103
M489 1848 WL_233 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=459600 $D=103
M490 1379 WL_234 1850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=462510 $D=103
M491 1852 WL_235 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=463000 $D=103
M492 1379 WL_236 1854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=465910 $D=103
M493 1856 WL_237 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=466400 $D=103
M494 1379 WL_238 1858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=469310 $D=103
M495 1860 WL_239 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=469800 $D=103
M496 1379 WL_240 1862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=472710 $D=103
M497 1864 WL_241 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=473200 $D=103
M498 1379 WL_242 1866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=476110 $D=103
M499 1868 WL_243 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=476600 $D=103
M500 1379 WL_244 1870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=479510 $D=103
M501 1872 WL_245 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=480000 $D=103
M502 1379 WL_246 1874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=482910 $D=103
M503 1876 WL_247 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=483400 $D=103
M504 1379 WL_248 1878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=486310 $D=103
M505 1880 WL_249 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=486800 $D=103
M506 1379 WL_250 1882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=489710 $D=103
M507 1884 WL_251 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=490200 $D=103
M508 1379 WL_252 1886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=493110 $D=103
M509 1888 WL_253 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=493600 $D=103
M510 1379 WL_254 1890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=496510 $D=103
M511 1892 WL_255 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=497000 $D=103
M512 1380 WL_0 1381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=64710 $D=103
M513 1383 WL_1 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=65200 $D=103
M514 1380 WL_2 1385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=68110 $D=103
M515 1387 WL_3 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=68600 $D=103
M516 1380 WL_4 1389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=71510 $D=103
M517 1391 WL_5 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=72000 $D=103
M518 1380 WL_6 1393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=74910 $D=103
M519 1395 WL_7 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=75400 $D=103
M520 1380 WL_8 1397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=78310 $D=103
M521 1399 WL_9 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=78800 $D=103
M522 1380 WL_10 1401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=81710 $D=103
M523 1403 WL_11 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=82200 $D=103
M524 1380 WL_12 1405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=85110 $D=103
M525 1407 WL_13 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=85600 $D=103
M526 1380 WL_14 1409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=88510 $D=103
M527 1411 WL_15 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=89000 $D=103
M528 1380 WL_16 1413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=91910 $D=103
M529 1415 WL_17 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=92400 $D=103
M530 1380 WL_18 1417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=95310 $D=103
M531 1419 WL_19 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=95800 $D=103
M532 1380 WL_20 1421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=98710 $D=103
M533 1423 WL_21 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=99200 $D=103
M534 1380 WL_22 1425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=102110 $D=103
M535 1427 WL_23 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=102600 $D=103
M536 1380 WL_24 1429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=105510 $D=103
M537 1431 WL_25 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=106000 $D=103
M538 1380 WL_26 1433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=108910 $D=103
M539 1435 WL_27 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=109400 $D=103
M540 1380 WL_28 1437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=112310 $D=103
M541 1439 WL_29 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=112800 $D=103
M542 1380 WL_30 1441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=115710 $D=103
M543 1443 WL_31 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=116200 $D=103
M544 1380 WL_32 1445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=119110 $D=103
M545 1447 WL_33 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=119600 $D=103
M546 1380 WL_34 1449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=122510 $D=103
M547 1451 WL_35 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=123000 $D=103
M548 1380 WL_36 1453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=125910 $D=103
M549 1455 WL_37 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=126400 $D=103
M550 1380 WL_38 1457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=129310 $D=103
M551 1459 WL_39 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=129800 $D=103
M552 1380 WL_40 1461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=132710 $D=103
M553 1463 WL_41 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=133200 $D=103
M554 1380 WL_42 1465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=136110 $D=103
M555 1467 WL_43 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=136600 $D=103
M556 1380 WL_44 1469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=139510 $D=103
M557 1471 WL_45 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=140000 $D=103
M558 1380 WL_46 1473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=142910 $D=103
M559 1475 WL_47 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=143400 $D=103
M560 1380 WL_48 1477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=146310 $D=103
M561 1479 WL_49 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=146800 $D=103
M562 1380 WL_50 1481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=149710 $D=103
M563 1483 WL_51 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=150200 $D=103
M564 1380 WL_52 1485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=153110 $D=103
M565 1487 WL_53 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=153600 $D=103
M566 1380 WL_54 1489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=156510 $D=103
M567 1491 WL_55 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=157000 $D=103
M568 1380 WL_56 1493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=159910 $D=103
M569 1495 WL_57 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=160400 $D=103
M570 1380 WL_58 1497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=163310 $D=103
M571 1499 WL_59 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=163800 $D=103
M572 1380 WL_60 1501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=166710 $D=103
M573 1503 WL_61 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=167200 $D=103
M574 1380 WL_62 1505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=170110 $D=103
M575 1507 WL_63 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=170600 $D=103
M576 1380 WL_64 1509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=173510 $D=103
M577 1511 WL_65 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=174000 $D=103
M578 1380 WL_66 1513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=176910 $D=103
M579 1515 WL_67 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=177400 $D=103
M580 1380 WL_68 1517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=180310 $D=103
M581 1519 WL_69 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=180800 $D=103
M582 1380 WL_70 1521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=183710 $D=103
M583 1523 WL_71 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=184200 $D=103
M584 1380 WL_72 1525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=187110 $D=103
M585 1527 WL_73 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=187600 $D=103
M586 1380 WL_74 1529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=190510 $D=103
M587 1531 WL_75 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=191000 $D=103
M588 1380 WL_76 1533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=193910 $D=103
M589 1535 WL_77 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=194400 $D=103
M590 1380 WL_78 1537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=197310 $D=103
M591 1539 WL_79 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=197800 $D=103
M592 1380 WL_80 1541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=200710 $D=103
M593 1543 WL_81 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=201200 $D=103
M594 1380 WL_82 1545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=204110 $D=103
M595 1547 WL_83 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=204600 $D=103
M596 1380 WL_84 1549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=207510 $D=103
M597 1551 WL_85 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=208000 $D=103
M598 1380 WL_86 1553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=210910 $D=103
M599 1555 WL_87 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=211400 $D=103
M600 1380 WL_88 1557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=214310 $D=103
M601 1559 WL_89 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=214800 $D=103
M602 1380 WL_90 1561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=217710 $D=103
M603 1563 WL_91 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=218200 $D=103
M604 1380 WL_92 1565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=221110 $D=103
M605 1567 WL_93 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=221600 $D=103
M606 1380 WL_94 1569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=224510 $D=103
M607 1571 WL_95 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=225000 $D=103
M608 1380 WL_96 1573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=227910 $D=103
M609 1575 WL_97 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=228400 $D=103
M610 1380 WL_98 1577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=231310 $D=103
M611 1579 WL_99 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=231800 $D=103
M612 1380 WL_100 1581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=234710 $D=103
M613 1583 WL_101 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=235200 $D=103
M614 1380 WL_102 1585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=238110 $D=103
M615 1587 WL_103 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=238600 $D=103
M616 1380 WL_104 1589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=241510 $D=103
M617 1591 WL_105 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=242000 $D=103
M618 1380 WL_106 1593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=244910 $D=103
M619 1595 WL_107 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=245400 $D=103
M620 1380 WL_108 1597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=248310 $D=103
M621 1599 WL_109 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=248800 $D=103
M622 1380 WL_110 1601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=251710 $D=103
M623 1603 WL_111 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=252200 $D=103
M624 1380 WL_112 1605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=255110 $D=103
M625 1607 WL_113 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=255600 $D=103
M626 1380 WL_114 1609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=258510 $D=103
M627 1611 WL_115 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=259000 $D=103
M628 1380 WL_116 1613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=261910 $D=103
M629 1615 WL_117 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=262400 $D=103
M630 1380 WL_118 1617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=265310 $D=103
M631 1619 WL_119 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=265800 $D=103
M632 1380 WL_120 1621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=268710 $D=103
M633 1623 WL_121 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=269200 $D=103
M634 1380 WL_122 1625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=272110 $D=103
M635 1627 WL_123 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=272600 $D=103
M636 1380 WL_124 1629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=275510 $D=103
M637 1631 WL_125 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=276000 $D=103
M638 1380 WL_126 1633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=278910 $D=103
M639 1635 WL_127 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=279400 $D=103
M640 1380 WL_128 1637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=282310 $D=103
M641 1639 WL_129 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=282800 $D=103
M642 1380 WL_130 1641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=285710 $D=103
M643 1643 WL_131 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=286200 $D=103
M644 1380 WL_132 1645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=289110 $D=103
M645 1647 WL_133 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=289600 $D=103
M646 1380 WL_134 1649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=292510 $D=103
M647 1651 WL_135 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=293000 $D=103
M648 1380 WL_136 1653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=295910 $D=103
M649 1655 WL_137 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=296400 $D=103
M650 1380 WL_138 1657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=299310 $D=103
M651 1659 WL_139 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=299800 $D=103
M652 1380 WL_140 1661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=302710 $D=103
M653 1663 WL_141 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=303200 $D=103
M654 1380 WL_142 1665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=306110 $D=103
M655 1667 WL_143 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=306600 $D=103
M656 1380 WL_144 1669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=309510 $D=103
M657 1671 WL_145 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=310000 $D=103
M658 1380 WL_146 1673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=312910 $D=103
M659 1675 WL_147 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=313400 $D=103
M660 1380 WL_148 1677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=316310 $D=103
M661 1679 WL_149 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=316800 $D=103
M662 1380 WL_150 1681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=319710 $D=103
M663 1683 WL_151 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=320200 $D=103
M664 1380 WL_152 1685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=323110 $D=103
M665 1687 WL_153 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=323600 $D=103
M666 1380 WL_154 1689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=326510 $D=103
M667 1691 WL_155 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=327000 $D=103
M668 1380 WL_156 1693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=329910 $D=103
M669 1695 WL_157 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=330400 $D=103
M670 1380 WL_158 1697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=333310 $D=103
M671 1699 WL_159 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=333800 $D=103
M672 1380 WL_160 1701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=336710 $D=103
M673 1703 WL_161 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=337200 $D=103
M674 1380 WL_162 1705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=340110 $D=103
M675 1707 WL_163 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=340600 $D=103
M676 1380 WL_164 1709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=343510 $D=103
M677 1711 WL_165 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=344000 $D=103
M678 1380 WL_166 1713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=346910 $D=103
M679 1715 WL_167 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=347400 $D=103
M680 1380 WL_168 1717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=350310 $D=103
M681 1719 WL_169 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=350800 $D=103
M682 1380 WL_170 1721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=353710 $D=103
M683 1723 WL_171 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=354200 $D=103
M684 1380 WL_172 1725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=357110 $D=103
M685 1727 WL_173 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=357600 $D=103
M686 1380 WL_174 1729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=360510 $D=103
M687 1731 WL_175 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=361000 $D=103
M688 1380 WL_176 1733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=363910 $D=103
M689 1735 WL_177 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=364400 $D=103
M690 1380 WL_178 1737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=367310 $D=103
M691 1739 WL_179 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=367800 $D=103
M692 1380 WL_180 1741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=370710 $D=103
M693 1743 WL_181 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=371200 $D=103
M694 1380 WL_182 1745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=374110 $D=103
M695 1747 WL_183 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=374600 $D=103
M696 1380 WL_184 1749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=377510 $D=103
M697 1751 WL_185 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=378000 $D=103
M698 1380 WL_186 1753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=380910 $D=103
M699 1755 WL_187 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=381400 $D=103
M700 1380 WL_188 1757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=384310 $D=103
M701 1759 WL_189 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=384800 $D=103
M702 1380 WL_190 1761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=387710 $D=103
M703 1763 WL_191 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=388200 $D=103
M704 1380 WL_192 1765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=391110 $D=103
M705 1767 WL_193 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=391600 $D=103
M706 1380 WL_194 1769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=394510 $D=103
M707 1771 WL_195 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=395000 $D=103
M708 1380 WL_196 1773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=397910 $D=103
M709 1775 WL_197 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=398400 $D=103
M710 1380 WL_198 1777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=401310 $D=103
M711 1779 WL_199 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=401800 $D=103
M712 1380 WL_200 1781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=404710 $D=103
M713 1783 WL_201 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=405200 $D=103
M714 1380 WL_202 1785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=408110 $D=103
M715 1787 WL_203 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=408600 $D=103
M716 1380 WL_204 1789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=411510 $D=103
M717 1791 WL_205 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=412000 $D=103
M718 1380 WL_206 1793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=414910 $D=103
M719 1795 WL_207 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=415400 $D=103
M720 1380 WL_208 1797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=418310 $D=103
M721 1799 WL_209 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=418800 $D=103
M722 1380 WL_210 1801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=421710 $D=103
M723 1803 WL_211 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=422200 $D=103
M724 1380 WL_212 1805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=425110 $D=103
M725 1807 WL_213 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=425600 $D=103
M726 1380 WL_214 1809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=428510 $D=103
M727 1811 WL_215 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=429000 $D=103
M728 1380 WL_216 1813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=431910 $D=103
M729 1815 WL_217 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=432400 $D=103
M730 1380 WL_218 1817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=435310 $D=103
M731 1819 WL_219 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=435800 $D=103
M732 1380 WL_220 1821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=438710 $D=103
M733 1823 WL_221 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=439200 $D=103
M734 1380 WL_222 1825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=442110 $D=103
M735 1827 WL_223 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=442600 $D=103
M736 1380 WL_224 1829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=445510 $D=103
M737 1831 WL_225 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=446000 $D=103
M738 1380 WL_226 1833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=448910 $D=103
M739 1835 WL_227 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=449400 $D=103
M740 1380 WL_228 1837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=452310 $D=103
M741 1839 WL_229 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=452800 $D=103
M742 1380 WL_230 1841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=455710 $D=103
M743 1843 WL_231 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=456200 $D=103
M744 1380 WL_232 1845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=459110 $D=103
M745 1847 WL_233 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=459600 $D=103
M746 1380 WL_234 1849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=462510 $D=103
M747 1851 WL_235 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=463000 $D=103
M748 1380 WL_236 1853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=465910 $D=103
M749 1855 WL_237 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=466400 $D=103
M750 1380 WL_238 1857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=469310 $D=103
M751 1859 WL_239 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=469800 $D=103
M752 1380 WL_240 1861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=472710 $D=103
M753 1863 WL_241 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=473200 $D=103
M754 1380 WL_242 1865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=476110 $D=103
M755 1867 WL_243 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=476600 $D=103
M756 1380 WL_244 1869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=479510 $D=103
M757 1871 WL_245 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=480000 $D=103
M758 1380 WL_246 1873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=482910 $D=103
M759 1875 WL_247 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=483400 $D=103
M760 1380 WL_248 1877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=486310 $D=103
M761 1879 WL_249 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=486800 $D=103
M762 1380 WL_250 1881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=489710 $D=103
M763 1883 WL_251 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=490200 $D=103
M764 1380 WL_252 1885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=493110 $D=103
M765 1887 WL_253 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=493600 $D=103
M766 1380 WL_254 1889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=496510 $D=103
M767 1891 WL_255 1380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=497000 $D=103
M768 1894 WL_0 1896 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=64710 $D=103
M769 1898 WL_1 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=65200 $D=103
M770 1894 WL_2 1900 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=68110 $D=103
M771 1902 WL_3 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=68600 $D=103
M772 1894 WL_4 1904 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=71510 $D=103
M773 1906 WL_5 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=72000 $D=103
M774 1894 WL_6 1908 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=74910 $D=103
M775 1910 WL_7 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=75400 $D=103
M776 1894 WL_8 1912 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=78310 $D=103
M777 1914 WL_9 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=78800 $D=103
M778 1894 WL_10 1916 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=81710 $D=103
M779 1918 WL_11 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=82200 $D=103
M780 1894 WL_12 1920 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=85110 $D=103
M781 1922 WL_13 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=85600 $D=103
M782 1894 WL_14 1924 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=88510 $D=103
M783 1926 WL_15 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=89000 $D=103
M784 1894 WL_16 1928 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=91910 $D=103
M785 1930 WL_17 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=92400 $D=103
M786 1894 WL_18 1932 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=95310 $D=103
M787 1934 WL_19 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=95800 $D=103
M788 1894 WL_20 1936 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=98710 $D=103
M789 1938 WL_21 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=99200 $D=103
M790 1894 WL_22 1940 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=102110 $D=103
M791 1942 WL_23 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=102600 $D=103
M792 1894 WL_24 1944 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=105510 $D=103
M793 1946 WL_25 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=106000 $D=103
M794 1894 WL_26 1948 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=108910 $D=103
M795 1950 WL_27 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=109400 $D=103
M796 1894 WL_28 1952 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=112310 $D=103
M797 1954 WL_29 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=112800 $D=103
M798 1894 WL_30 1956 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=115710 $D=103
M799 1958 WL_31 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=116200 $D=103
M800 1894 WL_32 1960 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=119110 $D=103
M801 1962 WL_33 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=119600 $D=103
M802 1894 WL_34 1964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=122510 $D=103
M803 1966 WL_35 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=123000 $D=103
M804 1894 WL_36 1968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=125910 $D=103
M805 1970 WL_37 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=126400 $D=103
M806 1894 WL_38 1972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=129310 $D=103
M807 1974 WL_39 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=129800 $D=103
M808 1894 WL_40 1976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=132710 $D=103
M809 1978 WL_41 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=133200 $D=103
M810 1894 WL_42 1980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=136110 $D=103
M811 1982 WL_43 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=136600 $D=103
M812 1894 WL_44 1984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=139510 $D=103
M813 1986 WL_45 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=140000 $D=103
M814 1894 WL_46 1988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=142910 $D=103
M815 1990 WL_47 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=143400 $D=103
M816 1894 WL_48 1992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=146310 $D=103
M817 1994 WL_49 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=146800 $D=103
M818 1894 WL_50 1996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=149710 $D=103
M819 1998 WL_51 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=150200 $D=103
M820 1894 WL_52 2000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=153110 $D=103
M821 2002 WL_53 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=153600 $D=103
M822 1894 WL_54 2004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=156510 $D=103
M823 2006 WL_55 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=157000 $D=103
M824 1894 WL_56 2008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=159910 $D=103
M825 2010 WL_57 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=160400 $D=103
M826 1894 WL_58 2012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=163310 $D=103
M827 2014 WL_59 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=163800 $D=103
M828 1894 WL_60 2016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=166710 $D=103
M829 2018 WL_61 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=167200 $D=103
M830 1894 WL_62 2020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=170110 $D=103
M831 2022 WL_63 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=170600 $D=103
M832 1894 WL_64 2024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=173510 $D=103
M833 2026 WL_65 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=174000 $D=103
M834 1894 WL_66 2028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=176910 $D=103
M835 2030 WL_67 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=177400 $D=103
M836 1894 WL_68 2032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=180310 $D=103
M837 2034 WL_69 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=180800 $D=103
M838 1894 WL_70 2036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=183710 $D=103
M839 2038 WL_71 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=184200 $D=103
M840 1894 WL_72 2040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=187110 $D=103
M841 2042 WL_73 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=187600 $D=103
M842 1894 WL_74 2044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=190510 $D=103
M843 2046 WL_75 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=191000 $D=103
M844 1894 WL_76 2048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=193910 $D=103
M845 2050 WL_77 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=194400 $D=103
M846 1894 WL_78 2052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=197310 $D=103
M847 2054 WL_79 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=197800 $D=103
M848 1894 WL_80 2056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=200710 $D=103
M849 2058 WL_81 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=201200 $D=103
M850 1894 WL_82 2060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=204110 $D=103
M851 2062 WL_83 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=204600 $D=103
M852 1894 WL_84 2064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=207510 $D=103
M853 2066 WL_85 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=208000 $D=103
M854 1894 WL_86 2068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=210910 $D=103
M855 2070 WL_87 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=211400 $D=103
M856 1894 WL_88 2072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=214310 $D=103
M857 2074 WL_89 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=214800 $D=103
M858 1894 WL_90 2076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=217710 $D=103
M859 2078 WL_91 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=218200 $D=103
M860 1894 WL_92 2080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=221110 $D=103
M861 2082 WL_93 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=221600 $D=103
M862 1894 WL_94 2084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=224510 $D=103
M863 2086 WL_95 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=225000 $D=103
M864 1894 WL_96 2088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=227910 $D=103
M865 2090 WL_97 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=228400 $D=103
M866 1894 WL_98 2092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=231310 $D=103
M867 2094 WL_99 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=231800 $D=103
M868 1894 WL_100 2096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=234710 $D=103
M869 2098 WL_101 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=235200 $D=103
M870 1894 WL_102 2100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=238110 $D=103
M871 2102 WL_103 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=238600 $D=103
M872 1894 WL_104 2104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=241510 $D=103
M873 2106 WL_105 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=242000 $D=103
M874 1894 WL_106 2108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=244910 $D=103
M875 2110 WL_107 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=245400 $D=103
M876 1894 WL_108 2112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=248310 $D=103
M877 2114 WL_109 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=248800 $D=103
M878 1894 WL_110 2116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=251710 $D=103
M879 2118 WL_111 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=252200 $D=103
M880 1894 WL_112 2120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=255110 $D=103
M881 2122 WL_113 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=255600 $D=103
M882 1894 WL_114 2124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=258510 $D=103
M883 2126 WL_115 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=259000 $D=103
M884 1894 WL_116 2128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=261910 $D=103
M885 2130 WL_117 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=262400 $D=103
M886 1894 WL_118 2132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=265310 $D=103
M887 2134 WL_119 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=265800 $D=103
M888 1894 WL_120 2136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=268710 $D=103
M889 2138 WL_121 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=269200 $D=103
M890 1894 WL_122 2140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=272110 $D=103
M891 2142 WL_123 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=272600 $D=103
M892 1894 WL_124 2144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=275510 $D=103
M893 2146 WL_125 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=276000 $D=103
M894 1894 WL_126 2148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=278910 $D=103
M895 2150 WL_127 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=279400 $D=103
M896 1894 WL_128 2152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=282310 $D=103
M897 2154 WL_129 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=282800 $D=103
M898 1894 WL_130 2156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=285710 $D=103
M899 2158 WL_131 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=286200 $D=103
M900 1894 WL_132 2160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=289110 $D=103
M901 2162 WL_133 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=289600 $D=103
M902 1894 WL_134 2164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=292510 $D=103
M903 2166 WL_135 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=293000 $D=103
M904 1894 WL_136 2168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=295910 $D=103
M905 2170 WL_137 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=296400 $D=103
M906 1894 WL_138 2172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=299310 $D=103
M907 2174 WL_139 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=299800 $D=103
M908 1894 WL_140 2176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=302710 $D=103
M909 2178 WL_141 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=303200 $D=103
M910 1894 WL_142 2180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=306110 $D=103
M911 2182 WL_143 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=306600 $D=103
M912 1894 WL_144 2184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=309510 $D=103
M913 2186 WL_145 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=310000 $D=103
M914 1894 WL_146 2188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=312910 $D=103
M915 2190 WL_147 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=313400 $D=103
M916 1894 WL_148 2192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=316310 $D=103
M917 2194 WL_149 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=316800 $D=103
M918 1894 WL_150 2196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=319710 $D=103
M919 2198 WL_151 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=320200 $D=103
M920 1894 WL_152 2200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=323110 $D=103
M921 2202 WL_153 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=323600 $D=103
M922 1894 WL_154 2204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=326510 $D=103
M923 2206 WL_155 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=327000 $D=103
M924 1894 WL_156 2208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=329910 $D=103
M925 2210 WL_157 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=330400 $D=103
M926 1894 WL_158 2212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=333310 $D=103
M927 2214 WL_159 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=333800 $D=103
M928 1894 WL_160 2216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=336710 $D=103
M929 2218 WL_161 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=337200 $D=103
M930 1894 WL_162 2220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=340110 $D=103
M931 2222 WL_163 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=340600 $D=103
M932 1894 WL_164 2224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=343510 $D=103
M933 2226 WL_165 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=344000 $D=103
M934 1894 WL_166 2228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=346910 $D=103
M935 2230 WL_167 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=347400 $D=103
M936 1894 WL_168 2232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=350310 $D=103
M937 2234 WL_169 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=350800 $D=103
M938 1894 WL_170 2236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=353710 $D=103
M939 2238 WL_171 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=354200 $D=103
M940 1894 WL_172 2240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=357110 $D=103
M941 2242 WL_173 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=357600 $D=103
M942 1894 WL_174 2244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=360510 $D=103
M943 2246 WL_175 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=361000 $D=103
M944 1894 WL_176 2248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=363910 $D=103
M945 2250 WL_177 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=364400 $D=103
M946 1894 WL_178 2252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=367310 $D=103
M947 2254 WL_179 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=367800 $D=103
M948 1894 WL_180 2256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=370710 $D=103
M949 2258 WL_181 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=371200 $D=103
M950 1894 WL_182 2260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=374110 $D=103
M951 2262 WL_183 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=374600 $D=103
M952 1894 WL_184 2264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=377510 $D=103
M953 2266 WL_185 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=378000 $D=103
M954 1894 WL_186 2268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=380910 $D=103
M955 2270 WL_187 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=381400 $D=103
M956 1894 WL_188 2272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=384310 $D=103
M957 2274 WL_189 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=384800 $D=103
M958 1894 WL_190 2276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=387710 $D=103
M959 2278 WL_191 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=388200 $D=103
M960 1894 WL_192 2280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=391110 $D=103
M961 2282 WL_193 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=391600 $D=103
M962 1894 WL_194 2284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=394510 $D=103
M963 2286 WL_195 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=395000 $D=103
M964 1894 WL_196 2288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=397910 $D=103
M965 2290 WL_197 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=398400 $D=103
M966 1894 WL_198 2292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=401310 $D=103
M967 2294 WL_199 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=401800 $D=103
M968 1894 WL_200 2296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=404710 $D=103
M969 2298 WL_201 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=405200 $D=103
M970 1894 WL_202 2300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=408110 $D=103
M971 2302 WL_203 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=408600 $D=103
M972 1894 WL_204 2304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=411510 $D=103
M973 2306 WL_205 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=412000 $D=103
M974 1894 WL_206 2308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=414910 $D=103
M975 2310 WL_207 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=415400 $D=103
M976 1894 WL_208 2312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=418310 $D=103
M977 2314 WL_209 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=418800 $D=103
M978 1894 WL_210 2316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=421710 $D=103
M979 2318 WL_211 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=422200 $D=103
M980 1894 WL_212 2320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=425110 $D=103
M981 2322 WL_213 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=425600 $D=103
M982 1894 WL_214 2324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=428510 $D=103
M983 2326 WL_215 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=429000 $D=103
M984 1894 WL_216 2328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=431910 $D=103
M985 2330 WL_217 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=432400 $D=103
M986 1894 WL_218 2332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=435310 $D=103
M987 2334 WL_219 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=435800 $D=103
M988 1894 WL_220 2336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=438710 $D=103
M989 2338 WL_221 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=439200 $D=103
M990 1894 WL_222 2340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=442110 $D=103
M991 2342 WL_223 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=442600 $D=103
M992 1894 WL_224 2344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=445510 $D=103
M993 2346 WL_225 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=446000 $D=103
M994 1894 WL_226 2348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=448910 $D=103
M995 2350 WL_227 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=449400 $D=103
M996 1894 WL_228 2352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=452310 $D=103
M997 2354 WL_229 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=452800 $D=103
M998 1894 WL_230 2356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=455710 $D=103
M999 2358 WL_231 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=456200 $D=103
M1000 1894 WL_232 2360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=459110 $D=103
M1001 2362 WL_233 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=459600 $D=103
M1002 1894 WL_234 2364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=462510 $D=103
M1003 2366 WL_235 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=463000 $D=103
M1004 1894 WL_236 2368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=465910 $D=103
M1005 2370 WL_237 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=466400 $D=103
M1006 1894 WL_238 2372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=469310 $D=103
M1007 2374 WL_239 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=469800 $D=103
M1008 1894 WL_240 2376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=472710 $D=103
M1009 2378 WL_241 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=473200 $D=103
M1010 1894 WL_242 2380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=476110 $D=103
M1011 2382 WL_243 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=476600 $D=103
M1012 1894 WL_244 2384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=479510 $D=103
M1013 2386 WL_245 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=480000 $D=103
M1014 1894 WL_246 2388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=482910 $D=103
M1015 2390 WL_247 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=483400 $D=103
M1016 1894 WL_248 2392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=486310 $D=103
M1017 2394 WL_249 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=486800 $D=103
M1018 1894 WL_250 2396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=489710 $D=103
M1019 2398 WL_251 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=490200 $D=103
M1020 1894 WL_252 2400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=493110 $D=103
M1021 2402 WL_253 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=493600 $D=103
M1022 1894 WL_254 2404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=496510 $D=103
M1023 2406 WL_255 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=497000 $D=103
M1024 1893 WL_0 1895 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=64710 $D=103
M1025 1897 WL_1 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=65200 $D=103
M1026 1893 WL_2 1899 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=68110 $D=103
M1027 1901 WL_3 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=68600 $D=103
M1028 1893 WL_4 1903 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=71510 $D=103
M1029 1905 WL_5 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=72000 $D=103
M1030 1893 WL_6 1907 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=74910 $D=103
M1031 1909 WL_7 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=75400 $D=103
M1032 1893 WL_8 1911 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=78310 $D=103
M1033 1913 WL_9 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=78800 $D=103
M1034 1893 WL_10 1915 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=81710 $D=103
M1035 1917 WL_11 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=82200 $D=103
M1036 1893 WL_12 1919 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=85110 $D=103
M1037 1921 WL_13 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=85600 $D=103
M1038 1893 WL_14 1923 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=88510 $D=103
M1039 1925 WL_15 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=89000 $D=103
M1040 1893 WL_16 1927 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=91910 $D=103
M1041 1929 WL_17 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=92400 $D=103
M1042 1893 WL_18 1931 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=95310 $D=103
M1043 1933 WL_19 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=95800 $D=103
M1044 1893 WL_20 1935 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=98710 $D=103
M1045 1937 WL_21 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=99200 $D=103
M1046 1893 WL_22 1939 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=102110 $D=103
M1047 1941 WL_23 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=102600 $D=103
M1048 1893 WL_24 1943 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=105510 $D=103
M1049 1945 WL_25 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=106000 $D=103
M1050 1893 WL_26 1947 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=108910 $D=103
M1051 1949 WL_27 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=109400 $D=103
M1052 1893 WL_28 1951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=112310 $D=103
M1053 1953 WL_29 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=112800 $D=103
M1054 1893 WL_30 1955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=115710 $D=103
M1055 1957 WL_31 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=116200 $D=103
M1056 1893 WL_32 1959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=119110 $D=103
M1057 1961 WL_33 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=119600 $D=103
M1058 1893 WL_34 1963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=122510 $D=103
M1059 1965 WL_35 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=123000 $D=103
M1060 1893 WL_36 1967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=125910 $D=103
M1061 1969 WL_37 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=126400 $D=103
M1062 1893 WL_38 1971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=129310 $D=103
M1063 1973 WL_39 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=129800 $D=103
M1064 1893 WL_40 1975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=132710 $D=103
M1065 1977 WL_41 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=133200 $D=103
M1066 1893 WL_42 1979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=136110 $D=103
M1067 1981 WL_43 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=136600 $D=103
M1068 1893 WL_44 1983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=139510 $D=103
M1069 1985 WL_45 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=140000 $D=103
M1070 1893 WL_46 1987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=142910 $D=103
M1071 1989 WL_47 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=143400 $D=103
M1072 1893 WL_48 1991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=146310 $D=103
M1073 1993 WL_49 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=146800 $D=103
M1074 1893 WL_50 1995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=149710 $D=103
M1075 1997 WL_51 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=150200 $D=103
M1076 1893 WL_52 1999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=153110 $D=103
M1077 2001 WL_53 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=153600 $D=103
M1078 1893 WL_54 2003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=156510 $D=103
M1079 2005 WL_55 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=157000 $D=103
M1080 1893 WL_56 2007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=159910 $D=103
M1081 2009 WL_57 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=160400 $D=103
M1082 1893 WL_58 2011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=163310 $D=103
M1083 2013 WL_59 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=163800 $D=103
M1084 1893 WL_60 2015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=166710 $D=103
M1085 2017 WL_61 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=167200 $D=103
M1086 1893 WL_62 2019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=170110 $D=103
M1087 2021 WL_63 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=170600 $D=103
M1088 1893 WL_64 2023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=173510 $D=103
M1089 2025 WL_65 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=174000 $D=103
M1090 1893 WL_66 2027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=176910 $D=103
M1091 2029 WL_67 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=177400 $D=103
M1092 1893 WL_68 2031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=180310 $D=103
M1093 2033 WL_69 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=180800 $D=103
M1094 1893 WL_70 2035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=183710 $D=103
M1095 2037 WL_71 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=184200 $D=103
M1096 1893 WL_72 2039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=187110 $D=103
M1097 2041 WL_73 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=187600 $D=103
M1098 1893 WL_74 2043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=190510 $D=103
M1099 2045 WL_75 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=191000 $D=103
M1100 1893 WL_76 2047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=193910 $D=103
M1101 2049 WL_77 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=194400 $D=103
M1102 1893 WL_78 2051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=197310 $D=103
M1103 2053 WL_79 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=197800 $D=103
M1104 1893 WL_80 2055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=200710 $D=103
M1105 2057 WL_81 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=201200 $D=103
M1106 1893 WL_82 2059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=204110 $D=103
M1107 2061 WL_83 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=204600 $D=103
M1108 1893 WL_84 2063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=207510 $D=103
M1109 2065 WL_85 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=208000 $D=103
M1110 1893 WL_86 2067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=210910 $D=103
M1111 2069 WL_87 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=211400 $D=103
M1112 1893 WL_88 2071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=214310 $D=103
M1113 2073 WL_89 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=214800 $D=103
M1114 1893 WL_90 2075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=217710 $D=103
M1115 2077 WL_91 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=218200 $D=103
M1116 1893 WL_92 2079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=221110 $D=103
M1117 2081 WL_93 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=221600 $D=103
M1118 1893 WL_94 2083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=224510 $D=103
M1119 2085 WL_95 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=225000 $D=103
M1120 1893 WL_96 2087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=227910 $D=103
M1121 2089 WL_97 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=228400 $D=103
M1122 1893 WL_98 2091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=231310 $D=103
M1123 2093 WL_99 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=231800 $D=103
M1124 1893 WL_100 2095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=234710 $D=103
M1125 2097 WL_101 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=235200 $D=103
M1126 1893 WL_102 2099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=238110 $D=103
M1127 2101 WL_103 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=238600 $D=103
M1128 1893 WL_104 2103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=241510 $D=103
M1129 2105 WL_105 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=242000 $D=103
M1130 1893 WL_106 2107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=244910 $D=103
M1131 2109 WL_107 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=245400 $D=103
M1132 1893 WL_108 2111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=248310 $D=103
M1133 2113 WL_109 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=248800 $D=103
M1134 1893 WL_110 2115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=251710 $D=103
M1135 2117 WL_111 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=252200 $D=103
M1136 1893 WL_112 2119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=255110 $D=103
M1137 2121 WL_113 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=255600 $D=103
M1138 1893 WL_114 2123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=258510 $D=103
M1139 2125 WL_115 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=259000 $D=103
M1140 1893 WL_116 2127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=261910 $D=103
M1141 2129 WL_117 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=262400 $D=103
M1142 1893 WL_118 2131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=265310 $D=103
M1143 2133 WL_119 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=265800 $D=103
M1144 1893 WL_120 2135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=268710 $D=103
M1145 2137 WL_121 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=269200 $D=103
M1146 1893 WL_122 2139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=272110 $D=103
M1147 2141 WL_123 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=272600 $D=103
M1148 1893 WL_124 2143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=275510 $D=103
M1149 2145 WL_125 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=276000 $D=103
M1150 1893 WL_126 2147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=278910 $D=103
M1151 2149 WL_127 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=279400 $D=103
M1152 1893 WL_128 2151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=282310 $D=103
M1153 2153 WL_129 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=282800 $D=103
M1154 1893 WL_130 2155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=285710 $D=103
M1155 2157 WL_131 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=286200 $D=103
M1156 1893 WL_132 2159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=289110 $D=103
M1157 2161 WL_133 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=289600 $D=103
M1158 1893 WL_134 2163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=292510 $D=103
M1159 2165 WL_135 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=293000 $D=103
M1160 1893 WL_136 2167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=295910 $D=103
M1161 2169 WL_137 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=296400 $D=103
M1162 1893 WL_138 2171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=299310 $D=103
M1163 2173 WL_139 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=299800 $D=103
M1164 1893 WL_140 2175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=302710 $D=103
M1165 2177 WL_141 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=303200 $D=103
M1166 1893 WL_142 2179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=306110 $D=103
M1167 2181 WL_143 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=306600 $D=103
M1168 1893 WL_144 2183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=309510 $D=103
M1169 2185 WL_145 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=310000 $D=103
M1170 1893 WL_146 2187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=312910 $D=103
M1171 2189 WL_147 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=313400 $D=103
M1172 1893 WL_148 2191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=316310 $D=103
M1173 2193 WL_149 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=316800 $D=103
M1174 1893 WL_150 2195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=319710 $D=103
M1175 2197 WL_151 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=320200 $D=103
M1176 1893 WL_152 2199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=323110 $D=103
M1177 2201 WL_153 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=323600 $D=103
M1178 1893 WL_154 2203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=326510 $D=103
M1179 2205 WL_155 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=327000 $D=103
M1180 1893 WL_156 2207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=329910 $D=103
M1181 2209 WL_157 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=330400 $D=103
M1182 1893 WL_158 2211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=333310 $D=103
M1183 2213 WL_159 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=333800 $D=103
M1184 1893 WL_160 2215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=336710 $D=103
M1185 2217 WL_161 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=337200 $D=103
M1186 1893 WL_162 2219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=340110 $D=103
M1187 2221 WL_163 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=340600 $D=103
M1188 1893 WL_164 2223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=343510 $D=103
M1189 2225 WL_165 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=344000 $D=103
M1190 1893 WL_166 2227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=346910 $D=103
M1191 2229 WL_167 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=347400 $D=103
M1192 1893 WL_168 2231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=350310 $D=103
M1193 2233 WL_169 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=350800 $D=103
M1194 1893 WL_170 2235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=353710 $D=103
M1195 2237 WL_171 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=354200 $D=103
M1196 1893 WL_172 2239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=357110 $D=103
M1197 2241 WL_173 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=357600 $D=103
M1198 1893 WL_174 2243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=360510 $D=103
M1199 2245 WL_175 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=361000 $D=103
M1200 1893 WL_176 2247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=363910 $D=103
M1201 2249 WL_177 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=364400 $D=103
M1202 1893 WL_178 2251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=367310 $D=103
M1203 2253 WL_179 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=367800 $D=103
M1204 1893 WL_180 2255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=370710 $D=103
M1205 2257 WL_181 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=371200 $D=103
M1206 1893 WL_182 2259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=374110 $D=103
M1207 2261 WL_183 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=374600 $D=103
M1208 1893 WL_184 2263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=377510 $D=103
M1209 2265 WL_185 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=378000 $D=103
M1210 1893 WL_186 2267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=380910 $D=103
M1211 2269 WL_187 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=381400 $D=103
M1212 1893 WL_188 2271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=384310 $D=103
M1213 2273 WL_189 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=384800 $D=103
M1214 1893 WL_190 2275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=387710 $D=103
M1215 2277 WL_191 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=388200 $D=103
M1216 1893 WL_192 2279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=391110 $D=103
M1217 2281 WL_193 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=391600 $D=103
M1218 1893 WL_194 2283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=394510 $D=103
M1219 2285 WL_195 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=395000 $D=103
M1220 1893 WL_196 2287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=397910 $D=103
M1221 2289 WL_197 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=398400 $D=103
M1222 1893 WL_198 2291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=401310 $D=103
M1223 2293 WL_199 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=401800 $D=103
M1224 1893 WL_200 2295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=404710 $D=103
M1225 2297 WL_201 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=405200 $D=103
M1226 1893 WL_202 2299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=408110 $D=103
M1227 2301 WL_203 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=408600 $D=103
M1228 1893 WL_204 2303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=411510 $D=103
M1229 2305 WL_205 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=412000 $D=103
M1230 1893 WL_206 2307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=414910 $D=103
M1231 2309 WL_207 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=415400 $D=103
M1232 1893 WL_208 2311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=418310 $D=103
M1233 2313 WL_209 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=418800 $D=103
M1234 1893 WL_210 2315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=421710 $D=103
M1235 2317 WL_211 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=422200 $D=103
M1236 1893 WL_212 2319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=425110 $D=103
M1237 2321 WL_213 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=425600 $D=103
M1238 1893 WL_214 2323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=428510 $D=103
M1239 2325 WL_215 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=429000 $D=103
M1240 1893 WL_216 2327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=431910 $D=103
M1241 2329 WL_217 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=432400 $D=103
M1242 1893 WL_218 2331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=435310 $D=103
M1243 2333 WL_219 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=435800 $D=103
M1244 1893 WL_220 2335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=438710 $D=103
M1245 2337 WL_221 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=439200 $D=103
M1246 1893 WL_222 2339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=442110 $D=103
M1247 2341 WL_223 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=442600 $D=103
M1248 1893 WL_224 2343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=445510 $D=103
M1249 2345 WL_225 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=446000 $D=103
M1250 1893 WL_226 2347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=448910 $D=103
M1251 2349 WL_227 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=449400 $D=103
M1252 1893 WL_228 2351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=452310 $D=103
M1253 2353 WL_229 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=452800 $D=103
M1254 1893 WL_230 2355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=455710 $D=103
M1255 2357 WL_231 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=456200 $D=103
M1256 1893 WL_232 2359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=459110 $D=103
M1257 2361 WL_233 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=459600 $D=103
M1258 1893 WL_234 2363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=462510 $D=103
M1259 2365 WL_235 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=463000 $D=103
M1260 1893 WL_236 2367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=465910 $D=103
M1261 2369 WL_237 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=466400 $D=103
M1262 1893 WL_238 2371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=469310 $D=103
M1263 2373 WL_239 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=469800 $D=103
M1264 1893 WL_240 2375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=472710 $D=103
M1265 2377 WL_241 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=473200 $D=103
M1266 1893 WL_242 2379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=476110 $D=103
M1267 2381 WL_243 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=476600 $D=103
M1268 1893 WL_244 2383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=479510 $D=103
M1269 2385 WL_245 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=480000 $D=103
M1270 1893 WL_246 2387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=482910 $D=103
M1271 2389 WL_247 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=483400 $D=103
M1272 1893 WL_248 2391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=486310 $D=103
M1273 2393 WL_249 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=486800 $D=103
M1274 1893 WL_250 2395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=489710 $D=103
M1275 2397 WL_251 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=490200 $D=103
M1276 1893 WL_252 2399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=493110 $D=103
M1277 2401 WL_253 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=493600 $D=103
M1278 1893 WL_254 2403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=496510 $D=103
M1279 2405 WL_255 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=497000 $D=103
M1280 2407 WL_0 2410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=64710 $D=103
M1281 2412 WL_1 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=65200 $D=103
M1282 2407 WL_2 2414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=68110 $D=103
M1283 2416 WL_3 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=68600 $D=103
M1284 2407 WL_4 2418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=71510 $D=103
M1285 2420 WL_5 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=72000 $D=103
M1286 2407 WL_6 2422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=74910 $D=103
M1287 2424 WL_7 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=75400 $D=103
M1288 2407 WL_8 2426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=78310 $D=103
M1289 2428 WL_9 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=78800 $D=103
M1290 2407 WL_10 2430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=81710 $D=103
M1291 2432 WL_11 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=82200 $D=103
M1292 2407 WL_12 2434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=85110 $D=103
M1293 2436 WL_13 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=85600 $D=103
M1294 2407 WL_14 2438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=88510 $D=103
M1295 2440 WL_15 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=89000 $D=103
M1296 2407 WL_16 2442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=91910 $D=103
M1297 2444 WL_17 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=92400 $D=103
M1298 2407 WL_18 2446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=95310 $D=103
M1299 2448 WL_19 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=95800 $D=103
M1300 2407 WL_20 2450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=98710 $D=103
M1301 2452 WL_21 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=99200 $D=103
M1302 2407 WL_22 2454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=102110 $D=103
M1303 2456 WL_23 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=102600 $D=103
M1304 2407 WL_24 2458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=105510 $D=103
M1305 2460 WL_25 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=106000 $D=103
M1306 2407 WL_26 2462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=108910 $D=103
M1307 2464 WL_27 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=109400 $D=103
M1308 2407 WL_28 2466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=112310 $D=103
M1309 2468 WL_29 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=112800 $D=103
M1310 2407 WL_30 2470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=115710 $D=103
M1311 2472 WL_31 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=116200 $D=103
M1312 2407 WL_32 2474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=119110 $D=103
M1313 2476 WL_33 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=119600 $D=103
M1314 2407 WL_34 2478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=122510 $D=103
M1315 2480 WL_35 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=123000 $D=103
M1316 2407 WL_36 2482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=125910 $D=103
M1317 2484 WL_37 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=126400 $D=103
M1318 2407 WL_38 2486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=129310 $D=103
M1319 2488 WL_39 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=129800 $D=103
M1320 2407 WL_40 2490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=132710 $D=103
M1321 2492 WL_41 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=133200 $D=103
M1322 2407 WL_42 2494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=136110 $D=103
M1323 2496 WL_43 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=136600 $D=103
M1324 2407 WL_44 2498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=139510 $D=103
M1325 2500 WL_45 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=140000 $D=103
M1326 2407 WL_46 2502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=142910 $D=103
M1327 2504 WL_47 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=143400 $D=103
M1328 2407 WL_48 2506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=146310 $D=103
M1329 2508 WL_49 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=146800 $D=103
M1330 2407 WL_50 2510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=149710 $D=103
M1331 2512 WL_51 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=150200 $D=103
M1332 2407 WL_52 2514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=153110 $D=103
M1333 2516 WL_53 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=153600 $D=103
M1334 2407 WL_54 2518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=156510 $D=103
M1335 2520 WL_55 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=157000 $D=103
M1336 2407 WL_56 2522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=159910 $D=103
M1337 2524 WL_57 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=160400 $D=103
M1338 2407 WL_58 2526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=163310 $D=103
M1339 2528 WL_59 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=163800 $D=103
M1340 2407 WL_60 2530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=166710 $D=103
M1341 2532 WL_61 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=167200 $D=103
M1342 2407 WL_62 2534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=170110 $D=103
M1343 2536 WL_63 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=170600 $D=103
M1344 2407 WL_64 2538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=173510 $D=103
M1345 2540 WL_65 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=174000 $D=103
M1346 2407 WL_66 2542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=176910 $D=103
M1347 2544 WL_67 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=177400 $D=103
M1348 2407 WL_68 2546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=180310 $D=103
M1349 2548 WL_69 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=180800 $D=103
M1350 2407 WL_70 2550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=183710 $D=103
M1351 2552 WL_71 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=184200 $D=103
M1352 2407 WL_72 2554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=187110 $D=103
M1353 2556 WL_73 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=187600 $D=103
M1354 2407 WL_74 2558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=190510 $D=103
M1355 2560 WL_75 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=191000 $D=103
M1356 2407 WL_76 2562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=193910 $D=103
M1357 2564 WL_77 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=194400 $D=103
M1358 2407 WL_78 2566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=197310 $D=103
M1359 2568 WL_79 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=197800 $D=103
M1360 2407 WL_80 2570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=200710 $D=103
M1361 2572 WL_81 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=201200 $D=103
M1362 2407 WL_82 2574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=204110 $D=103
M1363 2576 WL_83 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=204600 $D=103
M1364 2407 WL_84 2578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=207510 $D=103
M1365 2580 WL_85 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=208000 $D=103
M1366 2407 WL_86 2582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=210910 $D=103
M1367 2584 WL_87 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=211400 $D=103
M1368 2407 WL_88 2586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=214310 $D=103
M1369 2588 WL_89 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=214800 $D=103
M1370 2407 WL_90 2590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=217710 $D=103
M1371 2592 WL_91 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=218200 $D=103
M1372 2407 WL_92 2594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=221110 $D=103
M1373 2596 WL_93 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=221600 $D=103
M1374 2407 WL_94 2598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=224510 $D=103
M1375 2600 WL_95 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=225000 $D=103
M1376 2407 WL_96 2602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=227910 $D=103
M1377 2604 WL_97 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=228400 $D=103
M1378 2407 WL_98 2606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=231310 $D=103
M1379 2608 WL_99 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=231800 $D=103
M1380 2407 WL_100 2610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=234710 $D=103
M1381 2612 WL_101 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=235200 $D=103
M1382 2407 WL_102 2614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=238110 $D=103
M1383 2616 WL_103 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=238600 $D=103
M1384 2407 WL_104 2618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=241510 $D=103
M1385 2620 WL_105 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=242000 $D=103
M1386 2407 WL_106 2622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=244910 $D=103
M1387 2624 WL_107 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=245400 $D=103
M1388 2407 WL_108 2626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=248310 $D=103
M1389 2628 WL_109 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=248800 $D=103
M1390 2407 WL_110 2630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=251710 $D=103
M1391 2632 WL_111 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=252200 $D=103
M1392 2407 WL_112 2634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=255110 $D=103
M1393 2636 WL_113 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=255600 $D=103
M1394 2407 WL_114 2638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=258510 $D=103
M1395 2640 WL_115 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=259000 $D=103
M1396 2407 WL_116 2642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=261910 $D=103
M1397 2644 WL_117 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=262400 $D=103
M1398 2407 WL_118 2646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=265310 $D=103
M1399 2648 WL_119 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=265800 $D=103
M1400 2407 WL_120 2650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=268710 $D=103
M1401 2652 WL_121 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=269200 $D=103
M1402 2407 WL_122 2654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=272110 $D=103
M1403 2656 WL_123 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=272600 $D=103
M1404 2407 WL_124 2658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=275510 $D=103
M1405 2660 WL_125 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=276000 $D=103
M1406 2407 WL_126 2662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=278910 $D=103
M1407 2664 WL_127 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=279400 $D=103
M1408 2407 WL_128 2666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=282310 $D=103
M1409 2668 WL_129 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=282800 $D=103
M1410 2407 WL_130 2670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=285710 $D=103
M1411 2672 WL_131 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=286200 $D=103
M1412 2407 WL_132 2674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=289110 $D=103
M1413 2676 WL_133 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=289600 $D=103
M1414 2407 WL_134 2678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=292510 $D=103
M1415 2680 WL_135 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=293000 $D=103
M1416 2407 WL_136 2682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=295910 $D=103
M1417 2684 WL_137 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=296400 $D=103
M1418 2407 WL_138 2686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=299310 $D=103
M1419 2688 WL_139 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=299800 $D=103
M1420 2407 WL_140 2690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=302710 $D=103
M1421 2692 WL_141 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=303200 $D=103
M1422 2407 WL_142 2694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=306110 $D=103
M1423 2696 WL_143 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=306600 $D=103
M1424 2407 WL_144 2698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=309510 $D=103
M1425 2700 WL_145 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=310000 $D=103
M1426 2407 WL_146 2702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=312910 $D=103
M1427 2704 WL_147 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=313400 $D=103
M1428 2407 WL_148 2706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=316310 $D=103
M1429 2708 WL_149 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=316800 $D=103
M1430 2407 WL_150 2710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=319710 $D=103
M1431 2712 WL_151 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=320200 $D=103
M1432 2407 WL_152 2714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=323110 $D=103
M1433 2716 WL_153 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=323600 $D=103
M1434 2407 WL_154 2718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=326510 $D=103
M1435 2720 WL_155 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=327000 $D=103
M1436 2407 WL_156 2722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=329910 $D=103
M1437 2724 WL_157 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=330400 $D=103
M1438 2407 WL_158 2726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=333310 $D=103
M1439 2728 WL_159 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=333800 $D=103
M1440 2407 WL_160 2730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=336710 $D=103
M1441 2732 WL_161 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=337200 $D=103
M1442 2407 WL_162 2734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=340110 $D=103
M1443 2736 WL_163 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=340600 $D=103
M1444 2407 WL_164 2738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=343510 $D=103
M1445 2740 WL_165 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=344000 $D=103
M1446 2407 WL_166 2742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=346910 $D=103
M1447 2744 WL_167 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=347400 $D=103
M1448 2407 WL_168 2746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=350310 $D=103
M1449 2748 WL_169 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=350800 $D=103
M1450 2407 WL_170 2750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=353710 $D=103
M1451 2752 WL_171 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=354200 $D=103
M1452 2407 WL_172 2754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=357110 $D=103
M1453 2756 WL_173 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=357600 $D=103
M1454 2407 WL_174 2758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=360510 $D=103
M1455 2760 WL_175 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=361000 $D=103
M1456 2407 WL_176 2762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=363910 $D=103
M1457 2764 WL_177 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=364400 $D=103
M1458 2407 WL_178 2766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=367310 $D=103
M1459 2768 WL_179 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=367800 $D=103
M1460 2407 WL_180 2770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=370710 $D=103
M1461 2772 WL_181 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=371200 $D=103
M1462 2407 WL_182 2774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=374110 $D=103
M1463 2776 WL_183 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=374600 $D=103
M1464 2407 WL_184 2778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=377510 $D=103
M1465 2780 WL_185 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=378000 $D=103
M1466 2407 WL_186 2782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=380910 $D=103
M1467 2784 WL_187 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=381400 $D=103
M1468 2407 WL_188 2786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=384310 $D=103
M1469 2788 WL_189 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=384800 $D=103
M1470 2407 WL_190 2790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=387710 $D=103
M1471 2792 WL_191 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=388200 $D=103
M1472 2407 WL_192 2794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=391110 $D=103
M1473 2796 WL_193 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=391600 $D=103
M1474 2407 WL_194 2798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=394510 $D=103
M1475 2800 WL_195 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=395000 $D=103
M1476 2407 WL_196 2802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=397910 $D=103
M1477 2804 WL_197 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=398400 $D=103
M1478 2407 WL_198 2806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=401310 $D=103
M1479 2808 WL_199 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=401800 $D=103
M1480 2407 WL_200 2810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=404710 $D=103
M1481 2812 WL_201 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=405200 $D=103
M1482 2407 WL_202 2814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=408110 $D=103
M1483 2816 WL_203 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=408600 $D=103
M1484 2407 WL_204 2818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=411510 $D=103
M1485 2820 WL_205 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=412000 $D=103
M1486 2407 WL_206 2822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=414910 $D=103
M1487 2824 WL_207 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=415400 $D=103
M1488 2407 WL_208 2826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=418310 $D=103
M1489 2828 WL_209 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=418800 $D=103
M1490 2407 WL_210 2830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=421710 $D=103
M1491 2832 WL_211 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=422200 $D=103
M1492 2407 WL_212 2834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=425110 $D=103
M1493 2836 WL_213 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=425600 $D=103
M1494 2407 WL_214 2838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=428510 $D=103
M1495 2840 WL_215 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=429000 $D=103
M1496 2407 WL_216 2842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=431910 $D=103
M1497 2844 WL_217 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=432400 $D=103
M1498 2407 WL_218 2846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=435310 $D=103
M1499 2848 WL_219 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=435800 $D=103
M1500 2407 WL_220 2850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=438710 $D=103
M1501 2852 WL_221 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=439200 $D=103
M1502 2407 WL_222 2854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=442110 $D=103
M1503 2856 WL_223 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=442600 $D=103
M1504 2407 WL_224 2858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=445510 $D=103
M1505 2860 WL_225 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=446000 $D=103
M1506 2407 WL_226 2862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=448910 $D=103
M1507 2864 WL_227 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=449400 $D=103
M1508 2407 WL_228 2866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=452310 $D=103
M1509 2868 WL_229 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=452800 $D=103
M1510 2407 WL_230 2870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=455710 $D=103
M1511 2872 WL_231 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=456200 $D=103
M1512 2407 WL_232 2874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=459110 $D=103
M1513 2876 WL_233 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=459600 $D=103
M1514 2407 WL_234 2878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=462510 $D=103
M1515 2880 WL_235 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=463000 $D=103
M1516 2407 WL_236 2882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=465910 $D=103
M1517 2884 WL_237 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=466400 $D=103
M1518 2407 WL_238 2886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=469310 $D=103
M1519 2888 WL_239 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=469800 $D=103
M1520 2407 WL_240 2890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=472710 $D=103
M1521 2892 WL_241 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=473200 $D=103
M1522 2407 WL_242 2894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=476110 $D=103
M1523 2896 WL_243 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=476600 $D=103
M1524 2407 WL_244 2898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=479510 $D=103
M1525 2900 WL_245 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=480000 $D=103
M1526 2407 WL_246 2902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=482910 $D=103
M1527 2904 WL_247 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=483400 $D=103
M1528 2407 WL_248 2906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=486310 $D=103
M1529 2908 WL_249 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=486800 $D=103
M1530 2407 WL_250 2910 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=489710 $D=103
M1531 2912 WL_251 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=490200 $D=103
M1532 2407 WL_252 2914 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=493110 $D=103
M1533 2916 WL_253 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=493600 $D=103
M1534 2407 WL_254 2918 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=496510 $D=103
M1535 2920 WL_255 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=497000 $D=103
M1536 2408 WL_0 2409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=64710 $D=103
M1537 2411 WL_1 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=65200 $D=103
M1538 2408 WL_2 2413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=68110 $D=103
M1539 2415 WL_3 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=68600 $D=103
M1540 2408 WL_4 2417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=71510 $D=103
M1541 2419 WL_5 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=72000 $D=103
M1542 2408 WL_6 2421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=74910 $D=103
M1543 2423 WL_7 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=75400 $D=103
M1544 2408 WL_8 2425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=78310 $D=103
M1545 2427 WL_9 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=78800 $D=103
M1546 2408 WL_10 2429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=81710 $D=103
M1547 2431 WL_11 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=82200 $D=103
M1548 2408 WL_12 2433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=85110 $D=103
M1549 2435 WL_13 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=85600 $D=103
M1550 2408 WL_14 2437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=88510 $D=103
M1551 2439 WL_15 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=89000 $D=103
M1552 2408 WL_16 2441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=91910 $D=103
M1553 2443 WL_17 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=92400 $D=103
M1554 2408 WL_18 2445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=95310 $D=103
M1555 2447 WL_19 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=95800 $D=103
M1556 2408 WL_20 2449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=98710 $D=103
M1557 2451 WL_21 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=99200 $D=103
M1558 2408 WL_22 2453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=102110 $D=103
M1559 2455 WL_23 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=102600 $D=103
M1560 2408 WL_24 2457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=105510 $D=103
M1561 2459 WL_25 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=106000 $D=103
M1562 2408 WL_26 2461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=108910 $D=103
M1563 2463 WL_27 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=109400 $D=103
M1564 2408 WL_28 2465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=112310 $D=103
M1565 2467 WL_29 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=112800 $D=103
M1566 2408 WL_30 2469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=115710 $D=103
M1567 2471 WL_31 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=116200 $D=103
M1568 2408 WL_32 2473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=119110 $D=103
M1569 2475 WL_33 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=119600 $D=103
M1570 2408 WL_34 2477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=122510 $D=103
M1571 2479 WL_35 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=123000 $D=103
M1572 2408 WL_36 2481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=125910 $D=103
M1573 2483 WL_37 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=126400 $D=103
M1574 2408 WL_38 2485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=129310 $D=103
M1575 2487 WL_39 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=129800 $D=103
M1576 2408 WL_40 2489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=132710 $D=103
M1577 2491 WL_41 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=133200 $D=103
M1578 2408 WL_42 2493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=136110 $D=103
M1579 2495 WL_43 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=136600 $D=103
M1580 2408 WL_44 2497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=139510 $D=103
M1581 2499 WL_45 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=140000 $D=103
M1582 2408 WL_46 2501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=142910 $D=103
M1583 2503 WL_47 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=143400 $D=103
M1584 2408 WL_48 2505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=146310 $D=103
M1585 2507 WL_49 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=146800 $D=103
M1586 2408 WL_50 2509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=149710 $D=103
M1587 2511 WL_51 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=150200 $D=103
M1588 2408 WL_52 2513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=153110 $D=103
M1589 2515 WL_53 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=153600 $D=103
M1590 2408 WL_54 2517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=156510 $D=103
M1591 2519 WL_55 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=157000 $D=103
M1592 2408 WL_56 2521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=159910 $D=103
M1593 2523 WL_57 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=160400 $D=103
M1594 2408 WL_58 2525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=163310 $D=103
M1595 2527 WL_59 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=163800 $D=103
M1596 2408 WL_60 2529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=166710 $D=103
M1597 2531 WL_61 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=167200 $D=103
M1598 2408 WL_62 2533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=170110 $D=103
M1599 2535 WL_63 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=170600 $D=103
M1600 2408 WL_64 2537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=173510 $D=103
M1601 2539 WL_65 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=174000 $D=103
M1602 2408 WL_66 2541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=176910 $D=103
M1603 2543 WL_67 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=177400 $D=103
M1604 2408 WL_68 2545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=180310 $D=103
M1605 2547 WL_69 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=180800 $D=103
M1606 2408 WL_70 2549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=183710 $D=103
M1607 2551 WL_71 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=184200 $D=103
M1608 2408 WL_72 2553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=187110 $D=103
M1609 2555 WL_73 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=187600 $D=103
M1610 2408 WL_74 2557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=190510 $D=103
M1611 2559 WL_75 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=191000 $D=103
M1612 2408 WL_76 2561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=193910 $D=103
M1613 2563 WL_77 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=194400 $D=103
M1614 2408 WL_78 2565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=197310 $D=103
M1615 2567 WL_79 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=197800 $D=103
M1616 2408 WL_80 2569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=200710 $D=103
M1617 2571 WL_81 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=201200 $D=103
M1618 2408 WL_82 2573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=204110 $D=103
M1619 2575 WL_83 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=204600 $D=103
M1620 2408 WL_84 2577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=207510 $D=103
M1621 2579 WL_85 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=208000 $D=103
M1622 2408 WL_86 2581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=210910 $D=103
M1623 2583 WL_87 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=211400 $D=103
M1624 2408 WL_88 2585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=214310 $D=103
M1625 2587 WL_89 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=214800 $D=103
M1626 2408 WL_90 2589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=217710 $D=103
M1627 2591 WL_91 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=218200 $D=103
M1628 2408 WL_92 2593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=221110 $D=103
M1629 2595 WL_93 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=221600 $D=103
M1630 2408 WL_94 2597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=224510 $D=103
M1631 2599 WL_95 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=225000 $D=103
M1632 2408 WL_96 2601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=227910 $D=103
M1633 2603 WL_97 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=228400 $D=103
M1634 2408 WL_98 2605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=231310 $D=103
M1635 2607 WL_99 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=231800 $D=103
M1636 2408 WL_100 2609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=234710 $D=103
M1637 2611 WL_101 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=235200 $D=103
M1638 2408 WL_102 2613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=238110 $D=103
M1639 2615 WL_103 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=238600 $D=103
M1640 2408 WL_104 2617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=241510 $D=103
M1641 2619 WL_105 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=242000 $D=103
M1642 2408 WL_106 2621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=244910 $D=103
M1643 2623 WL_107 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=245400 $D=103
M1644 2408 WL_108 2625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=248310 $D=103
M1645 2627 WL_109 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=248800 $D=103
M1646 2408 WL_110 2629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=251710 $D=103
M1647 2631 WL_111 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=252200 $D=103
M1648 2408 WL_112 2633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=255110 $D=103
M1649 2635 WL_113 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=255600 $D=103
M1650 2408 WL_114 2637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=258510 $D=103
M1651 2639 WL_115 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=259000 $D=103
M1652 2408 WL_116 2641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=261910 $D=103
M1653 2643 WL_117 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=262400 $D=103
M1654 2408 WL_118 2645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=265310 $D=103
M1655 2647 WL_119 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=265800 $D=103
M1656 2408 WL_120 2649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=268710 $D=103
M1657 2651 WL_121 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=269200 $D=103
M1658 2408 WL_122 2653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=272110 $D=103
M1659 2655 WL_123 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=272600 $D=103
M1660 2408 WL_124 2657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=275510 $D=103
M1661 2659 WL_125 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=276000 $D=103
M1662 2408 WL_126 2661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=278910 $D=103
M1663 2663 WL_127 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=279400 $D=103
M1664 2408 WL_128 2665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=282310 $D=103
M1665 2667 WL_129 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=282800 $D=103
M1666 2408 WL_130 2669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=285710 $D=103
M1667 2671 WL_131 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=286200 $D=103
M1668 2408 WL_132 2673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=289110 $D=103
M1669 2675 WL_133 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=289600 $D=103
M1670 2408 WL_134 2677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=292510 $D=103
M1671 2679 WL_135 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=293000 $D=103
M1672 2408 WL_136 2681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=295910 $D=103
M1673 2683 WL_137 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=296400 $D=103
M1674 2408 WL_138 2685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=299310 $D=103
M1675 2687 WL_139 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=299800 $D=103
M1676 2408 WL_140 2689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=302710 $D=103
M1677 2691 WL_141 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=303200 $D=103
M1678 2408 WL_142 2693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=306110 $D=103
M1679 2695 WL_143 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=306600 $D=103
M1680 2408 WL_144 2697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=309510 $D=103
M1681 2699 WL_145 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=310000 $D=103
M1682 2408 WL_146 2701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=312910 $D=103
M1683 2703 WL_147 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=313400 $D=103
M1684 2408 WL_148 2705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=316310 $D=103
M1685 2707 WL_149 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=316800 $D=103
M1686 2408 WL_150 2709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=319710 $D=103
M1687 2711 WL_151 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=320200 $D=103
M1688 2408 WL_152 2713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=323110 $D=103
M1689 2715 WL_153 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=323600 $D=103
M1690 2408 WL_154 2717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=326510 $D=103
M1691 2719 WL_155 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=327000 $D=103
M1692 2408 WL_156 2721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=329910 $D=103
M1693 2723 WL_157 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=330400 $D=103
M1694 2408 WL_158 2725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=333310 $D=103
M1695 2727 WL_159 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=333800 $D=103
M1696 2408 WL_160 2729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=336710 $D=103
M1697 2731 WL_161 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=337200 $D=103
M1698 2408 WL_162 2733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=340110 $D=103
M1699 2735 WL_163 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=340600 $D=103
M1700 2408 WL_164 2737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=343510 $D=103
M1701 2739 WL_165 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=344000 $D=103
M1702 2408 WL_166 2741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=346910 $D=103
M1703 2743 WL_167 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=347400 $D=103
M1704 2408 WL_168 2745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=350310 $D=103
M1705 2747 WL_169 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=350800 $D=103
M1706 2408 WL_170 2749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=353710 $D=103
M1707 2751 WL_171 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=354200 $D=103
M1708 2408 WL_172 2753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=357110 $D=103
M1709 2755 WL_173 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=357600 $D=103
M1710 2408 WL_174 2757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=360510 $D=103
M1711 2759 WL_175 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=361000 $D=103
M1712 2408 WL_176 2761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=363910 $D=103
M1713 2763 WL_177 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=364400 $D=103
M1714 2408 WL_178 2765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=367310 $D=103
M1715 2767 WL_179 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=367800 $D=103
M1716 2408 WL_180 2769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=370710 $D=103
M1717 2771 WL_181 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=371200 $D=103
M1718 2408 WL_182 2773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=374110 $D=103
M1719 2775 WL_183 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=374600 $D=103
M1720 2408 WL_184 2777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=377510 $D=103
M1721 2779 WL_185 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=378000 $D=103
M1722 2408 WL_186 2781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=380910 $D=103
M1723 2783 WL_187 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=381400 $D=103
M1724 2408 WL_188 2785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=384310 $D=103
M1725 2787 WL_189 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=384800 $D=103
M1726 2408 WL_190 2789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=387710 $D=103
M1727 2791 WL_191 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=388200 $D=103
M1728 2408 WL_192 2793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=391110 $D=103
M1729 2795 WL_193 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=391600 $D=103
M1730 2408 WL_194 2797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=394510 $D=103
M1731 2799 WL_195 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=395000 $D=103
M1732 2408 WL_196 2801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=397910 $D=103
M1733 2803 WL_197 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=398400 $D=103
M1734 2408 WL_198 2805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=401310 $D=103
M1735 2807 WL_199 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=401800 $D=103
M1736 2408 WL_200 2809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=404710 $D=103
M1737 2811 WL_201 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=405200 $D=103
M1738 2408 WL_202 2813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=408110 $D=103
M1739 2815 WL_203 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=408600 $D=103
M1740 2408 WL_204 2817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=411510 $D=103
M1741 2819 WL_205 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=412000 $D=103
M1742 2408 WL_206 2821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=414910 $D=103
M1743 2823 WL_207 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=415400 $D=103
M1744 2408 WL_208 2825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=418310 $D=103
M1745 2827 WL_209 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=418800 $D=103
M1746 2408 WL_210 2829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=421710 $D=103
M1747 2831 WL_211 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=422200 $D=103
M1748 2408 WL_212 2833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=425110 $D=103
M1749 2835 WL_213 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=425600 $D=103
M1750 2408 WL_214 2837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=428510 $D=103
M1751 2839 WL_215 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=429000 $D=103
M1752 2408 WL_216 2841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=431910 $D=103
M1753 2843 WL_217 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=432400 $D=103
M1754 2408 WL_218 2845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=435310 $D=103
M1755 2847 WL_219 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=435800 $D=103
M1756 2408 WL_220 2849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=438710 $D=103
M1757 2851 WL_221 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=439200 $D=103
M1758 2408 WL_222 2853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=442110 $D=103
M1759 2855 WL_223 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=442600 $D=103
M1760 2408 WL_224 2857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=445510 $D=103
M1761 2859 WL_225 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=446000 $D=103
M1762 2408 WL_226 2861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=448910 $D=103
M1763 2863 WL_227 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=449400 $D=103
M1764 2408 WL_228 2865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=452310 $D=103
M1765 2867 WL_229 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=452800 $D=103
M1766 2408 WL_230 2869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=455710 $D=103
M1767 2871 WL_231 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=456200 $D=103
M1768 2408 WL_232 2873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=459110 $D=103
M1769 2875 WL_233 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=459600 $D=103
M1770 2408 WL_234 2877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=462510 $D=103
M1771 2879 WL_235 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=463000 $D=103
M1772 2408 WL_236 2881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=465910 $D=103
M1773 2883 WL_237 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=466400 $D=103
M1774 2408 WL_238 2885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=469310 $D=103
M1775 2887 WL_239 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=469800 $D=103
M1776 2408 WL_240 2889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=472710 $D=103
M1777 2891 WL_241 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=473200 $D=103
M1778 2408 WL_242 2893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=476110 $D=103
M1779 2895 WL_243 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=476600 $D=103
M1780 2408 WL_244 2897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=479510 $D=103
M1781 2899 WL_245 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=480000 $D=103
M1782 2408 WL_246 2901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=482910 $D=103
M1783 2903 WL_247 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=483400 $D=103
M1784 2408 WL_248 2905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=486310 $D=103
M1785 2907 WL_249 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=486800 $D=103
M1786 2408 WL_250 2909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=489710 $D=103
M1787 2911 WL_251 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=490200 $D=103
M1788 2408 WL_252 2913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=493110 $D=103
M1789 2915 WL_253 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=493600 $D=103
M1790 2408 WL_254 2917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=496510 $D=103
M1791 2919 WL_255 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=497000 $D=103
M1792 2922 WL_0 2924 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=64710 $D=103
M1793 2926 WL_1 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=65200 $D=103
M1794 2922 WL_2 2928 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=68110 $D=103
M1795 2930 WL_3 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=68600 $D=103
M1796 2922 WL_4 2932 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=71510 $D=103
M1797 2934 WL_5 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=72000 $D=103
M1798 2922 WL_6 2936 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=74910 $D=103
M1799 2938 WL_7 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=75400 $D=103
M1800 2922 WL_8 2940 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=78310 $D=103
M1801 2942 WL_9 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=78800 $D=103
M1802 2922 WL_10 2944 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=81710 $D=103
M1803 2946 WL_11 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=82200 $D=103
M1804 2922 WL_12 2948 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=85110 $D=103
M1805 2950 WL_13 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=85600 $D=103
M1806 2922 WL_14 2952 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=88510 $D=103
M1807 2954 WL_15 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=89000 $D=103
M1808 2922 WL_16 2956 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=91910 $D=103
M1809 2958 WL_17 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=92400 $D=103
M1810 2922 WL_18 2960 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=95310 $D=103
M1811 2962 WL_19 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=95800 $D=103
M1812 2922 WL_20 2964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=98710 $D=103
M1813 2966 WL_21 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=99200 $D=103
M1814 2922 WL_22 2968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=102110 $D=103
M1815 2970 WL_23 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=102600 $D=103
M1816 2922 WL_24 2972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=105510 $D=103
M1817 2974 WL_25 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=106000 $D=103
M1818 2922 WL_26 2976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=108910 $D=103
M1819 2978 WL_27 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=109400 $D=103
M1820 2922 WL_28 2980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=112310 $D=103
M1821 2982 WL_29 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=112800 $D=103
M1822 2922 WL_30 2984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=115710 $D=103
M1823 2986 WL_31 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=116200 $D=103
M1824 2922 WL_32 2988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=119110 $D=103
M1825 2990 WL_33 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=119600 $D=103
M1826 2922 WL_34 2992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=122510 $D=103
M1827 2994 WL_35 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=123000 $D=103
M1828 2922 WL_36 2996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=125910 $D=103
M1829 2998 WL_37 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=126400 $D=103
M1830 2922 WL_38 3000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=129310 $D=103
M1831 3002 WL_39 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=129800 $D=103
M1832 2922 WL_40 3004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=132710 $D=103
M1833 3006 WL_41 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=133200 $D=103
M1834 2922 WL_42 3008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=136110 $D=103
M1835 3010 WL_43 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=136600 $D=103
M1836 2922 WL_44 3012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=139510 $D=103
M1837 3014 WL_45 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=140000 $D=103
M1838 2922 WL_46 3016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=142910 $D=103
M1839 3018 WL_47 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=143400 $D=103
M1840 2922 WL_48 3020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=146310 $D=103
M1841 3022 WL_49 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=146800 $D=103
M1842 2922 WL_50 3024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=149710 $D=103
M1843 3026 WL_51 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=150200 $D=103
M1844 2922 WL_52 3028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=153110 $D=103
M1845 3030 WL_53 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=153600 $D=103
M1846 2922 WL_54 3032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=156510 $D=103
M1847 3034 WL_55 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=157000 $D=103
M1848 2922 WL_56 3036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=159910 $D=103
M1849 3038 WL_57 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=160400 $D=103
M1850 2922 WL_58 3040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=163310 $D=103
M1851 3042 WL_59 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=163800 $D=103
M1852 2922 WL_60 3044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=166710 $D=103
M1853 3046 WL_61 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=167200 $D=103
M1854 2922 WL_62 3048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=170110 $D=103
M1855 3050 WL_63 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=170600 $D=103
M1856 2922 WL_64 3052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=173510 $D=103
M1857 3054 WL_65 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=174000 $D=103
M1858 2922 WL_66 3056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=176910 $D=103
M1859 3058 WL_67 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=177400 $D=103
M1860 2922 WL_68 3060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=180310 $D=103
M1861 3062 WL_69 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=180800 $D=103
M1862 2922 WL_70 3064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=183710 $D=103
M1863 3066 WL_71 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=184200 $D=103
M1864 2922 WL_72 3068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=187110 $D=103
M1865 3070 WL_73 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=187600 $D=103
M1866 2922 WL_74 3072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=190510 $D=103
M1867 3074 WL_75 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=191000 $D=103
M1868 2922 WL_76 3076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=193910 $D=103
M1869 3078 WL_77 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=194400 $D=103
M1870 2922 WL_78 3080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=197310 $D=103
M1871 3082 WL_79 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=197800 $D=103
M1872 2922 WL_80 3084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=200710 $D=103
M1873 3086 WL_81 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=201200 $D=103
M1874 2922 WL_82 3088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=204110 $D=103
M1875 3090 WL_83 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=204600 $D=103
M1876 2922 WL_84 3092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=207510 $D=103
M1877 3094 WL_85 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=208000 $D=103
M1878 2922 WL_86 3096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=210910 $D=103
M1879 3098 WL_87 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=211400 $D=103
M1880 2922 WL_88 3100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=214310 $D=103
M1881 3102 WL_89 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=214800 $D=103
M1882 2922 WL_90 3104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=217710 $D=103
M1883 3106 WL_91 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=218200 $D=103
M1884 2922 WL_92 3108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=221110 $D=103
M1885 3110 WL_93 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=221600 $D=103
M1886 2922 WL_94 3112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=224510 $D=103
M1887 3114 WL_95 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=225000 $D=103
M1888 2922 WL_96 3116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=227910 $D=103
M1889 3118 WL_97 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=228400 $D=103
M1890 2922 WL_98 3120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=231310 $D=103
M1891 3122 WL_99 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=231800 $D=103
M1892 2922 WL_100 3124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=234710 $D=103
M1893 3126 WL_101 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=235200 $D=103
M1894 2922 WL_102 3128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=238110 $D=103
M1895 3130 WL_103 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=238600 $D=103
M1896 2922 WL_104 3132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=241510 $D=103
M1897 3134 WL_105 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=242000 $D=103
M1898 2922 WL_106 3136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=244910 $D=103
M1899 3138 WL_107 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=245400 $D=103
M1900 2922 WL_108 3140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=248310 $D=103
M1901 3142 WL_109 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=248800 $D=103
M1902 2922 WL_110 3144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=251710 $D=103
M1903 3146 WL_111 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=252200 $D=103
M1904 2922 WL_112 3148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=255110 $D=103
M1905 3150 WL_113 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=255600 $D=103
M1906 2922 WL_114 3152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=258510 $D=103
M1907 3154 WL_115 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=259000 $D=103
M1908 2922 WL_116 3156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=261910 $D=103
M1909 3158 WL_117 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=262400 $D=103
M1910 2922 WL_118 3160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=265310 $D=103
M1911 3162 WL_119 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=265800 $D=103
M1912 2922 WL_120 3164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=268710 $D=103
M1913 3166 WL_121 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=269200 $D=103
M1914 2922 WL_122 3168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=272110 $D=103
M1915 3170 WL_123 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=272600 $D=103
M1916 2922 WL_124 3172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=275510 $D=103
M1917 3174 WL_125 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=276000 $D=103
M1918 2922 WL_126 3176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=278910 $D=103
M1919 3178 WL_127 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=279400 $D=103
M1920 2922 WL_128 3180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=282310 $D=103
M1921 3182 WL_129 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=282800 $D=103
M1922 2922 WL_130 3184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=285710 $D=103
M1923 3186 WL_131 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=286200 $D=103
M1924 2922 WL_132 3188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=289110 $D=103
M1925 3190 WL_133 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=289600 $D=103
M1926 2922 WL_134 3192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=292510 $D=103
M1927 3194 WL_135 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=293000 $D=103
M1928 2922 WL_136 3196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=295910 $D=103
M1929 3198 WL_137 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=296400 $D=103
M1930 2922 WL_138 3200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=299310 $D=103
M1931 3202 WL_139 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=299800 $D=103
M1932 2922 WL_140 3204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=302710 $D=103
M1933 3206 WL_141 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=303200 $D=103
M1934 2922 WL_142 3208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=306110 $D=103
M1935 3210 WL_143 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=306600 $D=103
M1936 2922 WL_144 3212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=309510 $D=103
M1937 3214 WL_145 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=310000 $D=103
M1938 2922 WL_146 3216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=312910 $D=103
M1939 3218 WL_147 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=313400 $D=103
M1940 2922 WL_148 3220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=316310 $D=103
M1941 3222 WL_149 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=316800 $D=103
M1942 2922 WL_150 3224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=319710 $D=103
M1943 3226 WL_151 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=320200 $D=103
M1944 2922 WL_152 3228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=323110 $D=103
M1945 3230 WL_153 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=323600 $D=103
M1946 2922 WL_154 3232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=326510 $D=103
M1947 3234 WL_155 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=327000 $D=103
M1948 2922 WL_156 3236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=329910 $D=103
M1949 3238 WL_157 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=330400 $D=103
M1950 2922 WL_158 3240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=333310 $D=103
M1951 3242 WL_159 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=333800 $D=103
M1952 2922 WL_160 3244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=336710 $D=103
M1953 3246 WL_161 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=337200 $D=103
M1954 2922 WL_162 3248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=340110 $D=103
M1955 3250 WL_163 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=340600 $D=103
M1956 2922 WL_164 3252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=343510 $D=103
M1957 3254 WL_165 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=344000 $D=103
M1958 2922 WL_166 3256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=346910 $D=103
M1959 3258 WL_167 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=347400 $D=103
M1960 2922 WL_168 3260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=350310 $D=103
M1961 3262 WL_169 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=350800 $D=103
M1962 2922 WL_170 3264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=353710 $D=103
M1963 3266 WL_171 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=354200 $D=103
M1964 2922 WL_172 3268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=357110 $D=103
M1965 3270 WL_173 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=357600 $D=103
M1966 2922 WL_174 3272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=360510 $D=103
M1967 3274 WL_175 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=361000 $D=103
M1968 2922 WL_176 3276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=363910 $D=103
M1969 3278 WL_177 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=364400 $D=103
M1970 2922 WL_178 3280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=367310 $D=103
M1971 3282 WL_179 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=367800 $D=103
M1972 2922 WL_180 3284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=370710 $D=103
M1973 3286 WL_181 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=371200 $D=103
M1974 2922 WL_182 3288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=374110 $D=103
M1975 3290 WL_183 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=374600 $D=103
M1976 2922 WL_184 3292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=377510 $D=103
M1977 3294 WL_185 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=378000 $D=103
M1978 2922 WL_186 3296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=380910 $D=103
M1979 3298 WL_187 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=381400 $D=103
M1980 2922 WL_188 3300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=384310 $D=103
M1981 3302 WL_189 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=384800 $D=103
M1982 2922 WL_190 3304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=387710 $D=103
M1983 3306 WL_191 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=388200 $D=103
M1984 2922 WL_192 3308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=391110 $D=103
M1985 3310 WL_193 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=391600 $D=103
M1986 2922 WL_194 3312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=394510 $D=103
M1987 3314 WL_195 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=395000 $D=103
M1988 2922 WL_196 3316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=397910 $D=103
M1989 3318 WL_197 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=398400 $D=103
M1990 2922 WL_198 3320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=401310 $D=103
M1991 3322 WL_199 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=401800 $D=103
M1992 2922 WL_200 3324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=404710 $D=103
M1993 3326 WL_201 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=405200 $D=103
M1994 2922 WL_202 3328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=408110 $D=103
M1995 3330 WL_203 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=408600 $D=103
M1996 2922 WL_204 3332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=411510 $D=103
M1997 3334 WL_205 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=412000 $D=103
M1998 2922 WL_206 3336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=414910 $D=103
M1999 3338 WL_207 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=415400 $D=103
M2000 2922 WL_208 3340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=418310 $D=103
M2001 3342 WL_209 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=418800 $D=103
M2002 2922 WL_210 3344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=421710 $D=103
M2003 3346 WL_211 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=422200 $D=103
M2004 2922 WL_212 3348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=425110 $D=103
M2005 3350 WL_213 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=425600 $D=103
M2006 2922 WL_214 3352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=428510 $D=103
M2007 3354 WL_215 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=429000 $D=103
M2008 2922 WL_216 3356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=431910 $D=103
M2009 3358 WL_217 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=432400 $D=103
M2010 2922 WL_218 3360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=435310 $D=103
M2011 3362 WL_219 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=435800 $D=103
M2012 2922 WL_220 3364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=438710 $D=103
M2013 3366 WL_221 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=439200 $D=103
M2014 2922 WL_222 3368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=442110 $D=103
M2015 3370 WL_223 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=442600 $D=103
M2016 2922 WL_224 3372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=445510 $D=103
M2017 3374 WL_225 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=446000 $D=103
M2018 2922 WL_226 3376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=448910 $D=103
M2019 3378 WL_227 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=449400 $D=103
M2020 2922 WL_228 3380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=452310 $D=103
M2021 3382 WL_229 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=452800 $D=103
M2022 2922 WL_230 3384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=455710 $D=103
M2023 3386 WL_231 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=456200 $D=103
M2024 2922 WL_232 3388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=459110 $D=103
M2025 3390 WL_233 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=459600 $D=103
M2026 2922 WL_234 3392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=462510 $D=103
M2027 3394 WL_235 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=463000 $D=103
M2028 2922 WL_236 3396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=465910 $D=103
M2029 3398 WL_237 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=466400 $D=103
M2030 2922 WL_238 3400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=469310 $D=103
M2031 3402 WL_239 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=469800 $D=103
M2032 2922 WL_240 3404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=472710 $D=103
M2033 3406 WL_241 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=473200 $D=103
M2034 2922 WL_242 3408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=476110 $D=103
M2035 3410 WL_243 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=476600 $D=103
M2036 2922 WL_244 3412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=479510 $D=103
M2037 3414 WL_245 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=480000 $D=103
M2038 2922 WL_246 3416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=482910 $D=103
M2039 3418 WL_247 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=483400 $D=103
M2040 2922 WL_248 3420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=486310 $D=103
M2041 3422 WL_249 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=486800 $D=103
M2042 2922 WL_250 3424 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=489710 $D=103
M2043 3426 WL_251 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=490200 $D=103
M2044 2922 WL_252 3428 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=493110 $D=103
M2045 3430 WL_253 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=493600 $D=103
M2046 2922 WL_254 3432 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=496510 $D=103
M2047 3434 WL_255 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=497000 $D=103
M2048 2921 WL_0 2923 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=64710 $D=103
M2049 2925 WL_1 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=65200 $D=103
M2050 2921 WL_2 2927 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=68110 $D=103
M2051 2929 WL_3 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=68600 $D=103
M2052 2921 WL_4 2931 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=71510 $D=103
M2053 2933 WL_5 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=72000 $D=103
M2054 2921 WL_6 2935 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=74910 $D=103
M2055 2937 WL_7 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=75400 $D=103
M2056 2921 WL_8 2939 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=78310 $D=103
M2057 2941 WL_9 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=78800 $D=103
M2058 2921 WL_10 2943 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=81710 $D=103
M2059 2945 WL_11 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=82200 $D=103
M2060 2921 WL_12 2947 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=85110 $D=103
M2061 2949 WL_13 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=85600 $D=103
M2062 2921 WL_14 2951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=88510 $D=103
M2063 2953 WL_15 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=89000 $D=103
M2064 2921 WL_16 2955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=91910 $D=103
M2065 2957 WL_17 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=92400 $D=103
M2066 2921 WL_18 2959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=95310 $D=103
M2067 2961 WL_19 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=95800 $D=103
M2068 2921 WL_20 2963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=98710 $D=103
M2069 2965 WL_21 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=99200 $D=103
M2070 2921 WL_22 2967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=102110 $D=103
M2071 2969 WL_23 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=102600 $D=103
M2072 2921 WL_24 2971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=105510 $D=103
M2073 2973 WL_25 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=106000 $D=103
M2074 2921 WL_26 2975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=108910 $D=103
M2075 2977 WL_27 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=109400 $D=103
M2076 2921 WL_28 2979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=112310 $D=103
M2077 2981 WL_29 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=112800 $D=103
M2078 2921 WL_30 2983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=115710 $D=103
M2079 2985 WL_31 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=116200 $D=103
M2080 2921 WL_32 2987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=119110 $D=103
M2081 2989 WL_33 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=119600 $D=103
M2082 2921 WL_34 2991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=122510 $D=103
M2083 2993 WL_35 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=123000 $D=103
M2084 2921 WL_36 2995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=125910 $D=103
M2085 2997 WL_37 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=126400 $D=103
M2086 2921 WL_38 2999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=129310 $D=103
M2087 3001 WL_39 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=129800 $D=103
M2088 2921 WL_40 3003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=132710 $D=103
M2089 3005 WL_41 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=133200 $D=103
M2090 2921 WL_42 3007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=136110 $D=103
M2091 3009 WL_43 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=136600 $D=103
M2092 2921 WL_44 3011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=139510 $D=103
M2093 3013 WL_45 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=140000 $D=103
M2094 2921 WL_46 3015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=142910 $D=103
M2095 3017 WL_47 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=143400 $D=103
M2096 2921 WL_48 3019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=146310 $D=103
M2097 3021 WL_49 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=146800 $D=103
M2098 2921 WL_50 3023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=149710 $D=103
M2099 3025 WL_51 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=150200 $D=103
M2100 2921 WL_52 3027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=153110 $D=103
M2101 3029 WL_53 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=153600 $D=103
M2102 2921 WL_54 3031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=156510 $D=103
M2103 3033 WL_55 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=157000 $D=103
M2104 2921 WL_56 3035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=159910 $D=103
M2105 3037 WL_57 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=160400 $D=103
M2106 2921 WL_58 3039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=163310 $D=103
M2107 3041 WL_59 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=163800 $D=103
M2108 2921 WL_60 3043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=166710 $D=103
M2109 3045 WL_61 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=167200 $D=103
M2110 2921 WL_62 3047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=170110 $D=103
M2111 3049 WL_63 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=170600 $D=103
M2112 2921 WL_64 3051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=173510 $D=103
M2113 3053 WL_65 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=174000 $D=103
M2114 2921 WL_66 3055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=176910 $D=103
M2115 3057 WL_67 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=177400 $D=103
M2116 2921 WL_68 3059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=180310 $D=103
M2117 3061 WL_69 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=180800 $D=103
M2118 2921 WL_70 3063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=183710 $D=103
M2119 3065 WL_71 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=184200 $D=103
M2120 2921 WL_72 3067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=187110 $D=103
M2121 3069 WL_73 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=187600 $D=103
M2122 2921 WL_74 3071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=190510 $D=103
M2123 3073 WL_75 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=191000 $D=103
M2124 2921 WL_76 3075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=193910 $D=103
M2125 3077 WL_77 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=194400 $D=103
M2126 2921 WL_78 3079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=197310 $D=103
M2127 3081 WL_79 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=197800 $D=103
M2128 2921 WL_80 3083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=200710 $D=103
M2129 3085 WL_81 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=201200 $D=103
M2130 2921 WL_82 3087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=204110 $D=103
M2131 3089 WL_83 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=204600 $D=103
M2132 2921 WL_84 3091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=207510 $D=103
M2133 3093 WL_85 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=208000 $D=103
M2134 2921 WL_86 3095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=210910 $D=103
M2135 3097 WL_87 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=211400 $D=103
M2136 2921 WL_88 3099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=214310 $D=103
M2137 3101 WL_89 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=214800 $D=103
M2138 2921 WL_90 3103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=217710 $D=103
M2139 3105 WL_91 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=218200 $D=103
M2140 2921 WL_92 3107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=221110 $D=103
M2141 3109 WL_93 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=221600 $D=103
M2142 2921 WL_94 3111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=224510 $D=103
M2143 3113 WL_95 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=225000 $D=103
M2144 2921 WL_96 3115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=227910 $D=103
M2145 3117 WL_97 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=228400 $D=103
M2146 2921 WL_98 3119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=231310 $D=103
M2147 3121 WL_99 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=231800 $D=103
M2148 2921 WL_100 3123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=234710 $D=103
M2149 3125 WL_101 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=235200 $D=103
M2150 2921 WL_102 3127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=238110 $D=103
M2151 3129 WL_103 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=238600 $D=103
M2152 2921 WL_104 3131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=241510 $D=103
M2153 3133 WL_105 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=242000 $D=103
M2154 2921 WL_106 3135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=244910 $D=103
M2155 3137 WL_107 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=245400 $D=103
M2156 2921 WL_108 3139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=248310 $D=103
M2157 3141 WL_109 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=248800 $D=103
M2158 2921 WL_110 3143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=251710 $D=103
M2159 3145 WL_111 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=252200 $D=103
M2160 2921 WL_112 3147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=255110 $D=103
M2161 3149 WL_113 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=255600 $D=103
M2162 2921 WL_114 3151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=258510 $D=103
M2163 3153 WL_115 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=259000 $D=103
M2164 2921 WL_116 3155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=261910 $D=103
M2165 3157 WL_117 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=262400 $D=103
M2166 2921 WL_118 3159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=265310 $D=103
M2167 3161 WL_119 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=265800 $D=103
M2168 2921 WL_120 3163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=268710 $D=103
M2169 3165 WL_121 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=269200 $D=103
M2170 2921 WL_122 3167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=272110 $D=103
M2171 3169 WL_123 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=272600 $D=103
M2172 2921 WL_124 3171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=275510 $D=103
M2173 3173 WL_125 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=276000 $D=103
M2174 2921 WL_126 3175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=278910 $D=103
M2175 3177 WL_127 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=279400 $D=103
M2176 2921 WL_128 3179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=282310 $D=103
M2177 3181 WL_129 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=282800 $D=103
M2178 2921 WL_130 3183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=285710 $D=103
M2179 3185 WL_131 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=286200 $D=103
M2180 2921 WL_132 3187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=289110 $D=103
M2181 3189 WL_133 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=289600 $D=103
M2182 2921 WL_134 3191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=292510 $D=103
M2183 3193 WL_135 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=293000 $D=103
M2184 2921 WL_136 3195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=295910 $D=103
M2185 3197 WL_137 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=296400 $D=103
M2186 2921 WL_138 3199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=299310 $D=103
M2187 3201 WL_139 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=299800 $D=103
M2188 2921 WL_140 3203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=302710 $D=103
M2189 3205 WL_141 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=303200 $D=103
M2190 2921 WL_142 3207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=306110 $D=103
M2191 3209 WL_143 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=306600 $D=103
M2192 2921 WL_144 3211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=309510 $D=103
M2193 3213 WL_145 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=310000 $D=103
M2194 2921 WL_146 3215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=312910 $D=103
M2195 3217 WL_147 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=313400 $D=103
M2196 2921 WL_148 3219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=316310 $D=103
M2197 3221 WL_149 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=316800 $D=103
M2198 2921 WL_150 3223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=319710 $D=103
M2199 3225 WL_151 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=320200 $D=103
M2200 2921 WL_152 3227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=323110 $D=103
M2201 3229 WL_153 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=323600 $D=103
M2202 2921 WL_154 3231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=326510 $D=103
M2203 3233 WL_155 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=327000 $D=103
M2204 2921 WL_156 3235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=329910 $D=103
M2205 3237 WL_157 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=330400 $D=103
M2206 2921 WL_158 3239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=333310 $D=103
M2207 3241 WL_159 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=333800 $D=103
M2208 2921 WL_160 3243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=336710 $D=103
M2209 3245 WL_161 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=337200 $D=103
M2210 2921 WL_162 3247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=340110 $D=103
M2211 3249 WL_163 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=340600 $D=103
M2212 2921 WL_164 3251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=343510 $D=103
M2213 3253 WL_165 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=344000 $D=103
M2214 2921 WL_166 3255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=346910 $D=103
M2215 3257 WL_167 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=347400 $D=103
M2216 2921 WL_168 3259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=350310 $D=103
M2217 3261 WL_169 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=350800 $D=103
M2218 2921 WL_170 3263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=353710 $D=103
M2219 3265 WL_171 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=354200 $D=103
M2220 2921 WL_172 3267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=357110 $D=103
M2221 3269 WL_173 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=357600 $D=103
M2222 2921 WL_174 3271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=360510 $D=103
M2223 3273 WL_175 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=361000 $D=103
M2224 2921 WL_176 3275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=363910 $D=103
M2225 3277 WL_177 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=364400 $D=103
M2226 2921 WL_178 3279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=367310 $D=103
M2227 3281 WL_179 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=367800 $D=103
M2228 2921 WL_180 3283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=370710 $D=103
M2229 3285 WL_181 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=371200 $D=103
M2230 2921 WL_182 3287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=374110 $D=103
M2231 3289 WL_183 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=374600 $D=103
M2232 2921 WL_184 3291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=377510 $D=103
M2233 3293 WL_185 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=378000 $D=103
M2234 2921 WL_186 3295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=380910 $D=103
M2235 3297 WL_187 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=381400 $D=103
M2236 2921 WL_188 3299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=384310 $D=103
M2237 3301 WL_189 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=384800 $D=103
M2238 2921 WL_190 3303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=387710 $D=103
M2239 3305 WL_191 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=388200 $D=103
M2240 2921 WL_192 3307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=391110 $D=103
M2241 3309 WL_193 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=391600 $D=103
M2242 2921 WL_194 3311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=394510 $D=103
M2243 3313 WL_195 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=395000 $D=103
M2244 2921 WL_196 3315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=397910 $D=103
M2245 3317 WL_197 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=398400 $D=103
M2246 2921 WL_198 3319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=401310 $D=103
M2247 3321 WL_199 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=401800 $D=103
M2248 2921 WL_200 3323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=404710 $D=103
M2249 3325 WL_201 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=405200 $D=103
M2250 2921 WL_202 3327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=408110 $D=103
M2251 3329 WL_203 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=408600 $D=103
M2252 2921 WL_204 3331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=411510 $D=103
M2253 3333 WL_205 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=412000 $D=103
M2254 2921 WL_206 3335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=414910 $D=103
M2255 3337 WL_207 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=415400 $D=103
M2256 2921 WL_208 3339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=418310 $D=103
M2257 3341 WL_209 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=418800 $D=103
M2258 2921 WL_210 3343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=421710 $D=103
M2259 3345 WL_211 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=422200 $D=103
M2260 2921 WL_212 3347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=425110 $D=103
M2261 3349 WL_213 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=425600 $D=103
M2262 2921 WL_214 3351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=428510 $D=103
M2263 3353 WL_215 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=429000 $D=103
M2264 2921 WL_216 3355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=431910 $D=103
M2265 3357 WL_217 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=432400 $D=103
M2266 2921 WL_218 3359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=435310 $D=103
M2267 3361 WL_219 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=435800 $D=103
M2268 2921 WL_220 3363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=438710 $D=103
M2269 3365 WL_221 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=439200 $D=103
M2270 2921 WL_222 3367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=442110 $D=103
M2271 3369 WL_223 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=442600 $D=103
M2272 2921 WL_224 3371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=445510 $D=103
M2273 3373 WL_225 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=446000 $D=103
M2274 2921 WL_226 3375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=448910 $D=103
M2275 3377 WL_227 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=449400 $D=103
M2276 2921 WL_228 3379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=452310 $D=103
M2277 3381 WL_229 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=452800 $D=103
M2278 2921 WL_230 3383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=455710 $D=103
M2279 3385 WL_231 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=456200 $D=103
M2280 2921 WL_232 3387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=459110 $D=103
M2281 3389 WL_233 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=459600 $D=103
M2282 2921 WL_234 3391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=462510 $D=103
M2283 3393 WL_235 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=463000 $D=103
M2284 2921 WL_236 3395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=465910 $D=103
M2285 3397 WL_237 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=466400 $D=103
M2286 2921 WL_238 3399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=469310 $D=103
M2287 3401 WL_239 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=469800 $D=103
M2288 2921 WL_240 3403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=472710 $D=103
M2289 3405 WL_241 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=473200 $D=103
M2290 2921 WL_242 3407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=476110 $D=103
M2291 3409 WL_243 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=476600 $D=103
M2292 2921 WL_244 3411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=479510 $D=103
M2293 3413 WL_245 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=480000 $D=103
M2294 2921 WL_246 3415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=482910 $D=103
M2295 3417 WL_247 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=483400 $D=103
M2296 2921 WL_248 3419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=486310 $D=103
M2297 3421 WL_249 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=486800 $D=103
M2298 2921 WL_250 3423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=489710 $D=103
M2299 3425 WL_251 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=490200 $D=103
M2300 2921 WL_252 3427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=493110 $D=103
M2301 3429 WL_253 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=493600 $D=103
M2302 2921 WL_254 3431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=496510 $D=103
M2303 3433 WL_255 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=497000 $D=103
M2304 3435 WL_0 3438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=64710 $D=103
M2305 3440 WL_1 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=65200 $D=103
M2306 3435 WL_2 3442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=68110 $D=103
M2307 3444 WL_3 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=68600 $D=103
M2308 3435 WL_4 3446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=71510 $D=103
M2309 3448 WL_5 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=72000 $D=103
M2310 3435 WL_6 3450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=74910 $D=103
M2311 3452 WL_7 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=75400 $D=103
M2312 3435 WL_8 3454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=78310 $D=103
M2313 3456 WL_9 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=78800 $D=103
M2314 3435 WL_10 3458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=81710 $D=103
M2315 3460 WL_11 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=82200 $D=103
M2316 3435 WL_12 3462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=85110 $D=103
M2317 3464 WL_13 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=85600 $D=103
M2318 3435 WL_14 3466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=88510 $D=103
M2319 3468 WL_15 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=89000 $D=103
M2320 3435 WL_16 3470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=91910 $D=103
M2321 3472 WL_17 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=92400 $D=103
M2322 3435 WL_18 3474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=95310 $D=103
M2323 3476 WL_19 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=95800 $D=103
M2324 3435 WL_20 3478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=98710 $D=103
M2325 3480 WL_21 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=99200 $D=103
M2326 3435 WL_22 3482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=102110 $D=103
M2327 3484 WL_23 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=102600 $D=103
M2328 3435 WL_24 3486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=105510 $D=103
M2329 3488 WL_25 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=106000 $D=103
M2330 3435 WL_26 3490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=108910 $D=103
M2331 3492 WL_27 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=109400 $D=103
M2332 3435 WL_28 3494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=112310 $D=103
M2333 3496 WL_29 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=112800 $D=103
M2334 3435 WL_30 3498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=115710 $D=103
M2335 3500 WL_31 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=116200 $D=103
M2336 3435 WL_32 3502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=119110 $D=103
M2337 3504 WL_33 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=119600 $D=103
M2338 3435 WL_34 3506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=122510 $D=103
M2339 3508 WL_35 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=123000 $D=103
M2340 3435 WL_36 3510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=125910 $D=103
M2341 3512 WL_37 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=126400 $D=103
M2342 3435 WL_38 3514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=129310 $D=103
M2343 3516 WL_39 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=129800 $D=103
M2344 3435 WL_40 3518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=132710 $D=103
M2345 3520 WL_41 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=133200 $D=103
M2346 3435 WL_42 3522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=136110 $D=103
M2347 3524 WL_43 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=136600 $D=103
M2348 3435 WL_44 3526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=139510 $D=103
M2349 3528 WL_45 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=140000 $D=103
M2350 3435 WL_46 3530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=142910 $D=103
M2351 3532 WL_47 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=143400 $D=103
M2352 3435 WL_48 3534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=146310 $D=103
M2353 3536 WL_49 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=146800 $D=103
M2354 3435 WL_50 3538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=149710 $D=103
M2355 3540 WL_51 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=150200 $D=103
M2356 3435 WL_52 3542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=153110 $D=103
M2357 3544 WL_53 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=153600 $D=103
M2358 3435 WL_54 3546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=156510 $D=103
M2359 3548 WL_55 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=157000 $D=103
M2360 3435 WL_56 3550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=159910 $D=103
M2361 3552 WL_57 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=160400 $D=103
M2362 3435 WL_58 3554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=163310 $D=103
M2363 3556 WL_59 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=163800 $D=103
M2364 3435 WL_60 3558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=166710 $D=103
M2365 3560 WL_61 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=167200 $D=103
M2366 3435 WL_62 3562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=170110 $D=103
M2367 3564 WL_63 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=170600 $D=103
M2368 3435 WL_64 3566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=173510 $D=103
M2369 3568 WL_65 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=174000 $D=103
M2370 3435 WL_66 3570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=176910 $D=103
M2371 3572 WL_67 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=177400 $D=103
M2372 3435 WL_68 3574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=180310 $D=103
M2373 3576 WL_69 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=180800 $D=103
M2374 3435 WL_70 3578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=183710 $D=103
M2375 3580 WL_71 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=184200 $D=103
M2376 3435 WL_72 3582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=187110 $D=103
M2377 3584 WL_73 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=187600 $D=103
M2378 3435 WL_74 3586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=190510 $D=103
M2379 3588 WL_75 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=191000 $D=103
M2380 3435 WL_76 3590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=193910 $D=103
M2381 3592 WL_77 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=194400 $D=103
M2382 3435 WL_78 3594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=197310 $D=103
M2383 3596 WL_79 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=197800 $D=103
M2384 3435 WL_80 3598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=200710 $D=103
M2385 3600 WL_81 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=201200 $D=103
M2386 3435 WL_82 3602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=204110 $D=103
M2387 3604 WL_83 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=204600 $D=103
M2388 3435 WL_84 3606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=207510 $D=103
M2389 3608 WL_85 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=208000 $D=103
M2390 3435 WL_86 3610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=210910 $D=103
M2391 3612 WL_87 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=211400 $D=103
M2392 3435 WL_88 3614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=214310 $D=103
M2393 3616 WL_89 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=214800 $D=103
M2394 3435 WL_90 3618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=217710 $D=103
M2395 3620 WL_91 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=218200 $D=103
M2396 3435 WL_92 3622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=221110 $D=103
M2397 3624 WL_93 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=221600 $D=103
M2398 3435 WL_94 3626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=224510 $D=103
M2399 3628 WL_95 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=225000 $D=103
M2400 3435 WL_96 3630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=227910 $D=103
M2401 3632 WL_97 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=228400 $D=103
M2402 3435 WL_98 3634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=231310 $D=103
M2403 3636 WL_99 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=231800 $D=103
M2404 3435 WL_100 3638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=234710 $D=103
M2405 3640 WL_101 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=235200 $D=103
M2406 3435 WL_102 3642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=238110 $D=103
M2407 3644 WL_103 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=238600 $D=103
M2408 3435 WL_104 3646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=241510 $D=103
M2409 3648 WL_105 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=242000 $D=103
M2410 3435 WL_106 3650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=244910 $D=103
M2411 3652 WL_107 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=245400 $D=103
M2412 3435 WL_108 3654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=248310 $D=103
M2413 3656 WL_109 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=248800 $D=103
M2414 3435 WL_110 3658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=251710 $D=103
M2415 3660 WL_111 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=252200 $D=103
M2416 3435 WL_112 3662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=255110 $D=103
M2417 3664 WL_113 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=255600 $D=103
M2418 3435 WL_114 3666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=258510 $D=103
M2419 3668 WL_115 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=259000 $D=103
M2420 3435 WL_116 3670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=261910 $D=103
M2421 3672 WL_117 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=262400 $D=103
M2422 3435 WL_118 3674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=265310 $D=103
M2423 3676 WL_119 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=265800 $D=103
M2424 3435 WL_120 3678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=268710 $D=103
M2425 3680 WL_121 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=269200 $D=103
M2426 3435 WL_122 3682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=272110 $D=103
M2427 3684 WL_123 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=272600 $D=103
M2428 3435 WL_124 3686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=275510 $D=103
M2429 3688 WL_125 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=276000 $D=103
M2430 3435 WL_126 3690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=278910 $D=103
M2431 3692 WL_127 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=279400 $D=103
M2432 3435 WL_128 3694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=282310 $D=103
M2433 3696 WL_129 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=282800 $D=103
M2434 3435 WL_130 3698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=285710 $D=103
M2435 3700 WL_131 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=286200 $D=103
M2436 3435 WL_132 3702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=289110 $D=103
M2437 3704 WL_133 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=289600 $D=103
M2438 3435 WL_134 3706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=292510 $D=103
M2439 3708 WL_135 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=293000 $D=103
M2440 3435 WL_136 3710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=295910 $D=103
M2441 3712 WL_137 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=296400 $D=103
M2442 3435 WL_138 3714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=299310 $D=103
M2443 3716 WL_139 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=299800 $D=103
M2444 3435 WL_140 3718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=302710 $D=103
M2445 3720 WL_141 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=303200 $D=103
M2446 3435 WL_142 3722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=306110 $D=103
M2447 3724 WL_143 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=306600 $D=103
M2448 3435 WL_144 3726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=309510 $D=103
M2449 3728 WL_145 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=310000 $D=103
M2450 3435 WL_146 3730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=312910 $D=103
M2451 3732 WL_147 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=313400 $D=103
M2452 3435 WL_148 3734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=316310 $D=103
M2453 3736 WL_149 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=316800 $D=103
M2454 3435 WL_150 3738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=319710 $D=103
M2455 3740 WL_151 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=320200 $D=103
M2456 3435 WL_152 3742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=323110 $D=103
M2457 3744 WL_153 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=323600 $D=103
M2458 3435 WL_154 3746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=326510 $D=103
M2459 3748 WL_155 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=327000 $D=103
M2460 3435 WL_156 3750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=329910 $D=103
M2461 3752 WL_157 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=330400 $D=103
M2462 3435 WL_158 3754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=333310 $D=103
M2463 3756 WL_159 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=333800 $D=103
M2464 3435 WL_160 3758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=336710 $D=103
M2465 3760 WL_161 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=337200 $D=103
M2466 3435 WL_162 3762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=340110 $D=103
M2467 3764 WL_163 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=340600 $D=103
M2468 3435 WL_164 3766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=343510 $D=103
M2469 3768 WL_165 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=344000 $D=103
M2470 3435 WL_166 3770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=346910 $D=103
M2471 3772 WL_167 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=347400 $D=103
M2472 3435 WL_168 3774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=350310 $D=103
M2473 3776 WL_169 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=350800 $D=103
M2474 3435 WL_170 3778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=353710 $D=103
M2475 3780 WL_171 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=354200 $D=103
M2476 3435 WL_172 3782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=357110 $D=103
M2477 3784 WL_173 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=357600 $D=103
M2478 3435 WL_174 3786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=360510 $D=103
M2479 3788 WL_175 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=361000 $D=103
M2480 3435 WL_176 3790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=363910 $D=103
M2481 3792 WL_177 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=364400 $D=103
M2482 3435 WL_178 3794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=367310 $D=103
M2483 3796 WL_179 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=367800 $D=103
M2484 3435 WL_180 3798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=370710 $D=103
M2485 3800 WL_181 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=371200 $D=103
M2486 3435 WL_182 3802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=374110 $D=103
M2487 3804 WL_183 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=374600 $D=103
M2488 3435 WL_184 3806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=377510 $D=103
M2489 3808 WL_185 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=378000 $D=103
M2490 3435 WL_186 3810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=380910 $D=103
M2491 3812 WL_187 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=381400 $D=103
M2492 3435 WL_188 3814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=384310 $D=103
M2493 3816 WL_189 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=384800 $D=103
M2494 3435 WL_190 3818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=387710 $D=103
M2495 3820 WL_191 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=388200 $D=103
M2496 3435 WL_192 3822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=391110 $D=103
M2497 3824 WL_193 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=391600 $D=103
M2498 3435 WL_194 3826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=394510 $D=103
M2499 3828 WL_195 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=395000 $D=103
M2500 3435 WL_196 3830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=397910 $D=103
M2501 3832 WL_197 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=398400 $D=103
M2502 3435 WL_198 3834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=401310 $D=103
M2503 3836 WL_199 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=401800 $D=103
M2504 3435 WL_200 3838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=404710 $D=103
M2505 3840 WL_201 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=405200 $D=103
M2506 3435 WL_202 3842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=408110 $D=103
M2507 3844 WL_203 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=408600 $D=103
M2508 3435 WL_204 3846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=411510 $D=103
M2509 3848 WL_205 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=412000 $D=103
M2510 3435 WL_206 3850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=414910 $D=103
M2511 3852 WL_207 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=415400 $D=103
M2512 3435 WL_208 3854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=418310 $D=103
M2513 3856 WL_209 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=418800 $D=103
M2514 3435 WL_210 3858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=421710 $D=103
M2515 3860 WL_211 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=422200 $D=103
M2516 3435 WL_212 3862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=425110 $D=103
M2517 3864 WL_213 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=425600 $D=103
M2518 3435 WL_214 3866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=428510 $D=103
M2519 3868 WL_215 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=429000 $D=103
M2520 3435 WL_216 3870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=431910 $D=103
M2521 3872 WL_217 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=432400 $D=103
M2522 3435 WL_218 3874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=435310 $D=103
M2523 3876 WL_219 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=435800 $D=103
M2524 3435 WL_220 3878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=438710 $D=103
M2525 3880 WL_221 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=439200 $D=103
M2526 3435 WL_222 3882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=442110 $D=103
M2527 3884 WL_223 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=442600 $D=103
M2528 3435 WL_224 3886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=445510 $D=103
M2529 3888 WL_225 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=446000 $D=103
M2530 3435 WL_226 3890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=448910 $D=103
M2531 3892 WL_227 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=449400 $D=103
M2532 3435 WL_228 3894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=452310 $D=103
M2533 3896 WL_229 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=452800 $D=103
M2534 3435 WL_230 3898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=455710 $D=103
M2535 3900 WL_231 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=456200 $D=103
M2536 3435 WL_232 3902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=459110 $D=103
M2537 3904 WL_233 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=459600 $D=103
M2538 3435 WL_234 3906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=462510 $D=103
M2539 3908 WL_235 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=463000 $D=103
M2540 3435 WL_236 3910 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=465910 $D=103
M2541 3912 WL_237 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=466400 $D=103
M2542 3435 WL_238 3914 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=469310 $D=103
M2543 3916 WL_239 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=469800 $D=103
M2544 3435 WL_240 3918 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=472710 $D=103
M2545 3920 WL_241 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=473200 $D=103
M2546 3435 WL_242 3922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=476110 $D=103
M2547 3924 WL_243 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=476600 $D=103
M2548 3435 WL_244 3926 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=479510 $D=103
M2549 3928 WL_245 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=480000 $D=103
M2550 3435 WL_246 3930 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=482910 $D=103
M2551 3932 WL_247 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=483400 $D=103
M2552 3435 WL_248 3934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=486310 $D=103
M2553 3936 WL_249 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=486800 $D=103
M2554 3435 WL_250 3938 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=489710 $D=103
M2555 3940 WL_251 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=490200 $D=103
M2556 3435 WL_252 3942 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=493110 $D=103
M2557 3944 WL_253 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=493600 $D=103
M2558 3435 WL_254 3946 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=496510 $D=103
M2559 3948 WL_255 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=497000 $D=103
M2560 3436 WL_0 3437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=64710 $D=103
M2561 3439 WL_1 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=65200 $D=103
M2562 3436 WL_2 3441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=68110 $D=103
M2563 3443 WL_3 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=68600 $D=103
M2564 3436 WL_4 3445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=71510 $D=103
M2565 3447 WL_5 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=72000 $D=103
M2566 3436 WL_6 3449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=74910 $D=103
M2567 3451 WL_7 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=75400 $D=103
M2568 3436 WL_8 3453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=78310 $D=103
M2569 3455 WL_9 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=78800 $D=103
M2570 3436 WL_10 3457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=81710 $D=103
M2571 3459 WL_11 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=82200 $D=103
M2572 3436 WL_12 3461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=85110 $D=103
M2573 3463 WL_13 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=85600 $D=103
M2574 3436 WL_14 3465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=88510 $D=103
M2575 3467 WL_15 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=89000 $D=103
M2576 3436 WL_16 3469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=91910 $D=103
M2577 3471 WL_17 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=92400 $D=103
M2578 3436 WL_18 3473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=95310 $D=103
M2579 3475 WL_19 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=95800 $D=103
M2580 3436 WL_20 3477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=98710 $D=103
M2581 3479 WL_21 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=99200 $D=103
M2582 3436 WL_22 3481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=102110 $D=103
M2583 3483 WL_23 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=102600 $D=103
M2584 3436 WL_24 3485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=105510 $D=103
M2585 3487 WL_25 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=106000 $D=103
M2586 3436 WL_26 3489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=108910 $D=103
M2587 3491 WL_27 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=109400 $D=103
M2588 3436 WL_28 3493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=112310 $D=103
M2589 3495 WL_29 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=112800 $D=103
M2590 3436 WL_30 3497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=115710 $D=103
M2591 3499 WL_31 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=116200 $D=103
M2592 3436 WL_32 3501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=119110 $D=103
M2593 3503 WL_33 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=119600 $D=103
M2594 3436 WL_34 3505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=122510 $D=103
M2595 3507 WL_35 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=123000 $D=103
M2596 3436 WL_36 3509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=125910 $D=103
M2597 3511 WL_37 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=126400 $D=103
M2598 3436 WL_38 3513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=129310 $D=103
M2599 3515 WL_39 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=129800 $D=103
M2600 3436 WL_40 3517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=132710 $D=103
M2601 3519 WL_41 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=133200 $D=103
M2602 3436 WL_42 3521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=136110 $D=103
M2603 3523 WL_43 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=136600 $D=103
M2604 3436 WL_44 3525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=139510 $D=103
M2605 3527 WL_45 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=140000 $D=103
M2606 3436 WL_46 3529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=142910 $D=103
M2607 3531 WL_47 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=143400 $D=103
M2608 3436 WL_48 3533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=146310 $D=103
M2609 3535 WL_49 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=146800 $D=103
M2610 3436 WL_50 3537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=149710 $D=103
M2611 3539 WL_51 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=150200 $D=103
M2612 3436 WL_52 3541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=153110 $D=103
M2613 3543 WL_53 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=153600 $D=103
M2614 3436 WL_54 3545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=156510 $D=103
M2615 3547 WL_55 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=157000 $D=103
M2616 3436 WL_56 3549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=159910 $D=103
M2617 3551 WL_57 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=160400 $D=103
M2618 3436 WL_58 3553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=163310 $D=103
M2619 3555 WL_59 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=163800 $D=103
M2620 3436 WL_60 3557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=166710 $D=103
M2621 3559 WL_61 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=167200 $D=103
M2622 3436 WL_62 3561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=170110 $D=103
M2623 3563 WL_63 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=170600 $D=103
M2624 3436 WL_64 3565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=173510 $D=103
M2625 3567 WL_65 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=174000 $D=103
M2626 3436 WL_66 3569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=176910 $D=103
M2627 3571 WL_67 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=177400 $D=103
M2628 3436 WL_68 3573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=180310 $D=103
M2629 3575 WL_69 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=180800 $D=103
M2630 3436 WL_70 3577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=183710 $D=103
M2631 3579 WL_71 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=184200 $D=103
M2632 3436 WL_72 3581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=187110 $D=103
M2633 3583 WL_73 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=187600 $D=103
M2634 3436 WL_74 3585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=190510 $D=103
M2635 3587 WL_75 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=191000 $D=103
M2636 3436 WL_76 3589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=193910 $D=103
M2637 3591 WL_77 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=194400 $D=103
M2638 3436 WL_78 3593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=197310 $D=103
M2639 3595 WL_79 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=197800 $D=103
M2640 3436 WL_80 3597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=200710 $D=103
M2641 3599 WL_81 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=201200 $D=103
M2642 3436 WL_82 3601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=204110 $D=103
M2643 3603 WL_83 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=204600 $D=103
M2644 3436 WL_84 3605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=207510 $D=103
M2645 3607 WL_85 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=208000 $D=103
M2646 3436 WL_86 3609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=210910 $D=103
M2647 3611 WL_87 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=211400 $D=103
M2648 3436 WL_88 3613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=214310 $D=103
M2649 3615 WL_89 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=214800 $D=103
M2650 3436 WL_90 3617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=217710 $D=103
M2651 3619 WL_91 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=218200 $D=103
M2652 3436 WL_92 3621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=221110 $D=103
M2653 3623 WL_93 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=221600 $D=103
M2654 3436 WL_94 3625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=224510 $D=103
M2655 3627 WL_95 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=225000 $D=103
M2656 3436 WL_96 3629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=227910 $D=103
M2657 3631 WL_97 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=228400 $D=103
M2658 3436 WL_98 3633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=231310 $D=103
M2659 3635 WL_99 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=231800 $D=103
M2660 3436 WL_100 3637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=234710 $D=103
M2661 3639 WL_101 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=235200 $D=103
M2662 3436 WL_102 3641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=238110 $D=103
M2663 3643 WL_103 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=238600 $D=103
M2664 3436 WL_104 3645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=241510 $D=103
M2665 3647 WL_105 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=242000 $D=103
M2666 3436 WL_106 3649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=244910 $D=103
M2667 3651 WL_107 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=245400 $D=103
M2668 3436 WL_108 3653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=248310 $D=103
M2669 3655 WL_109 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=248800 $D=103
M2670 3436 WL_110 3657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=251710 $D=103
M2671 3659 WL_111 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=252200 $D=103
M2672 3436 WL_112 3661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=255110 $D=103
M2673 3663 WL_113 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=255600 $D=103
M2674 3436 WL_114 3665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=258510 $D=103
M2675 3667 WL_115 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=259000 $D=103
M2676 3436 WL_116 3669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=261910 $D=103
M2677 3671 WL_117 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=262400 $D=103
M2678 3436 WL_118 3673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=265310 $D=103
M2679 3675 WL_119 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=265800 $D=103
M2680 3436 WL_120 3677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=268710 $D=103
M2681 3679 WL_121 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=269200 $D=103
M2682 3436 WL_122 3681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=272110 $D=103
M2683 3683 WL_123 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=272600 $D=103
M2684 3436 WL_124 3685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=275510 $D=103
M2685 3687 WL_125 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=276000 $D=103
M2686 3436 WL_126 3689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=278910 $D=103
M2687 3691 WL_127 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=279400 $D=103
M2688 3436 WL_128 3693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=282310 $D=103
M2689 3695 WL_129 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=282800 $D=103
M2690 3436 WL_130 3697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=285710 $D=103
M2691 3699 WL_131 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=286200 $D=103
M2692 3436 WL_132 3701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=289110 $D=103
M2693 3703 WL_133 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=289600 $D=103
M2694 3436 WL_134 3705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=292510 $D=103
M2695 3707 WL_135 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=293000 $D=103
M2696 3436 WL_136 3709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=295910 $D=103
M2697 3711 WL_137 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=296400 $D=103
M2698 3436 WL_138 3713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=299310 $D=103
M2699 3715 WL_139 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=299800 $D=103
M2700 3436 WL_140 3717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=302710 $D=103
M2701 3719 WL_141 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=303200 $D=103
M2702 3436 WL_142 3721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=306110 $D=103
M2703 3723 WL_143 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=306600 $D=103
M2704 3436 WL_144 3725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=309510 $D=103
M2705 3727 WL_145 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=310000 $D=103
M2706 3436 WL_146 3729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=312910 $D=103
M2707 3731 WL_147 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=313400 $D=103
M2708 3436 WL_148 3733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=316310 $D=103
M2709 3735 WL_149 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=316800 $D=103
M2710 3436 WL_150 3737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=319710 $D=103
M2711 3739 WL_151 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=320200 $D=103
M2712 3436 WL_152 3741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=323110 $D=103
M2713 3743 WL_153 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=323600 $D=103
M2714 3436 WL_154 3745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=326510 $D=103
M2715 3747 WL_155 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=327000 $D=103
M2716 3436 WL_156 3749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=329910 $D=103
M2717 3751 WL_157 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=330400 $D=103
M2718 3436 WL_158 3753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=333310 $D=103
M2719 3755 WL_159 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=333800 $D=103
M2720 3436 WL_160 3757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=336710 $D=103
M2721 3759 WL_161 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=337200 $D=103
M2722 3436 WL_162 3761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=340110 $D=103
M2723 3763 WL_163 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=340600 $D=103
M2724 3436 WL_164 3765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=343510 $D=103
M2725 3767 WL_165 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=344000 $D=103
M2726 3436 WL_166 3769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=346910 $D=103
M2727 3771 WL_167 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=347400 $D=103
M2728 3436 WL_168 3773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=350310 $D=103
M2729 3775 WL_169 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=350800 $D=103
M2730 3436 WL_170 3777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=353710 $D=103
M2731 3779 WL_171 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=354200 $D=103
M2732 3436 WL_172 3781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=357110 $D=103
M2733 3783 WL_173 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=357600 $D=103
M2734 3436 WL_174 3785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=360510 $D=103
M2735 3787 WL_175 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=361000 $D=103
M2736 3436 WL_176 3789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=363910 $D=103
M2737 3791 WL_177 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=364400 $D=103
M2738 3436 WL_178 3793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=367310 $D=103
M2739 3795 WL_179 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=367800 $D=103
M2740 3436 WL_180 3797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=370710 $D=103
M2741 3799 WL_181 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=371200 $D=103
M2742 3436 WL_182 3801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=374110 $D=103
M2743 3803 WL_183 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=374600 $D=103
M2744 3436 WL_184 3805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=377510 $D=103
M2745 3807 WL_185 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=378000 $D=103
M2746 3436 WL_186 3809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=380910 $D=103
M2747 3811 WL_187 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=381400 $D=103
M2748 3436 WL_188 3813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=384310 $D=103
M2749 3815 WL_189 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=384800 $D=103
M2750 3436 WL_190 3817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=387710 $D=103
M2751 3819 WL_191 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=388200 $D=103
M2752 3436 WL_192 3821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=391110 $D=103
M2753 3823 WL_193 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=391600 $D=103
M2754 3436 WL_194 3825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=394510 $D=103
M2755 3827 WL_195 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=395000 $D=103
M2756 3436 WL_196 3829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=397910 $D=103
M2757 3831 WL_197 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=398400 $D=103
M2758 3436 WL_198 3833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=401310 $D=103
M2759 3835 WL_199 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=401800 $D=103
M2760 3436 WL_200 3837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=404710 $D=103
M2761 3839 WL_201 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=405200 $D=103
M2762 3436 WL_202 3841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=408110 $D=103
M2763 3843 WL_203 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=408600 $D=103
M2764 3436 WL_204 3845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=411510 $D=103
M2765 3847 WL_205 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=412000 $D=103
M2766 3436 WL_206 3849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=414910 $D=103
M2767 3851 WL_207 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=415400 $D=103
M2768 3436 WL_208 3853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=418310 $D=103
M2769 3855 WL_209 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=418800 $D=103
M2770 3436 WL_210 3857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=421710 $D=103
M2771 3859 WL_211 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=422200 $D=103
M2772 3436 WL_212 3861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=425110 $D=103
M2773 3863 WL_213 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=425600 $D=103
M2774 3436 WL_214 3865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=428510 $D=103
M2775 3867 WL_215 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=429000 $D=103
M2776 3436 WL_216 3869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=431910 $D=103
M2777 3871 WL_217 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=432400 $D=103
M2778 3436 WL_218 3873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=435310 $D=103
M2779 3875 WL_219 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=435800 $D=103
M2780 3436 WL_220 3877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=438710 $D=103
M2781 3879 WL_221 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=439200 $D=103
M2782 3436 WL_222 3881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=442110 $D=103
M2783 3883 WL_223 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=442600 $D=103
M2784 3436 WL_224 3885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=445510 $D=103
M2785 3887 WL_225 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=446000 $D=103
M2786 3436 WL_226 3889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=448910 $D=103
M2787 3891 WL_227 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=449400 $D=103
M2788 3436 WL_228 3893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=452310 $D=103
M2789 3895 WL_229 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=452800 $D=103
M2790 3436 WL_230 3897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=455710 $D=103
M2791 3899 WL_231 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=456200 $D=103
M2792 3436 WL_232 3901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=459110 $D=103
M2793 3903 WL_233 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=459600 $D=103
M2794 3436 WL_234 3905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=462510 $D=103
M2795 3907 WL_235 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=463000 $D=103
M2796 3436 WL_236 3909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=465910 $D=103
M2797 3911 WL_237 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=466400 $D=103
M2798 3436 WL_238 3913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=469310 $D=103
M2799 3915 WL_239 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=469800 $D=103
M2800 3436 WL_240 3917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=472710 $D=103
M2801 3919 WL_241 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=473200 $D=103
M2802 3436 WL_242 3921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=476110 $D=103
M2803 3923 WL_243 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=476600 $D=103
M2804 3436 WL_244 3925 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=479510 $D=103
M2805 3927 WL_245 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=480000 $D=103
M2806 3436 WL_246 3929 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=482910 $D=103
M2807 3931 WL_247 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=483400 $D=103
M2808 3436 WL_248 3933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=486310 $D=103
M2809 3935 WL_249 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=486800 $D=103
M2810 3436 WL_250 3937 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=489710 $D=103
M2811 3939 WL_251 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=490200 $D=103
M2812 3436 WL_252 3941 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=493110 $D=103
M2813 3943 WL_253 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=493600 $D=103
M2814 3436 WL_254 3945 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=496510 $D=103
M2815 3947 WL_255 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=497000 $D=103
M2816 3950 WL_0 3952 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=64710 $D=103
M2817 3954 WL_1 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=65200 $D=103
M2818 3950 WL_2 3956 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=68110 $D=103
M2819 3958 WL_3 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=68600 $D=103
M2820 3950 WL_4 3960 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=71510 $D=103
M2821 3962 WL_5 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=72000 $D=103
M2822 3950 WL_6 3964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=74910 $D=103
M2823 3966 WL_7 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=75400 $D=103
M2824 3950 WL_8 3968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=78310 $D=103
M2825 3970 WL_9 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=78800 $D=103
M2826 3950 WL_10 3972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=81710 $D=103
M2827 3974 WL_11 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=82200 $D=103
M2828 3950 WL_12 3976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=85110 $D=103
M2829 3978 WL_13 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=85600 $D=103
M2830 3950 WL_14 3980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=88510 $D=103
M2831 3982 WL_15 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=89000 $D=103
M2832 3950 WL_16 3984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=91910 $D=103
M2833 3986 WL_17 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=92400 $D=103
M2834 3950 WL_18 3988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=95310 $D=103
M2835 3990 WL_19 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=95800 $D=103
M2836 3950 WL_20 3992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=98710 $D=103
M2837 3994 WL_21 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=99200 $D=103
M2838 3950 WL_22 3996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=102110 $D=103
M2839 3998 WL_23 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=102600 $D=103
M2840 3950 WL_24 4000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=105510 $D=103
M2841 4002 WL_25 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=106000 $D=103
M2842 3950 WL_26 4004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=108910 $D=103
M2843 4006 WL_27 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=109400 $D=103
M2844 3950 WL_28 4008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=112310 $D=103
M2845 4010 WL_29 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=112800 $D=103
M2846 3950 WL_30 4012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=115710 $D=103
M2847 4014 WL_31 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=116200 $D=103
M2848 3950 WL_32 4016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=119110 $D=103
M2849 4018 WL_33 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=119600 $D=103
M2850 3950 WL_34 4020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=122510 $D=103
M2851 4022 WL_35 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=123000 $D=103
M2852 3950 WL_36 4024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=125910 $D=103
M2853 4026 WL_37 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=126400 $D=103
M2854 3950 WL_38 4028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=129310 $D=103
M2855 4030 WL_39 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=129800 $D=103
M2856 3950 WL_40 4032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=132710 $D=103
M2857 4034 WL_41 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=133200 $D=103
M2858 3950 WL_42 4036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=136110 $D=103
M2859 4038 WL_43 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=136600 $D=103
M2860 3950 WL_44 4040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=139510 $D=103
M2861 4042 WL_45 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=140000 $D=103
M2862 3950 WL_46 4044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=142910 $D=103
M2863 4046 WL_47 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=143400 $D=103
M2864 3950 WL_48 4048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=146310 $D=103
M2865 4050 WL_49 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=146800 $D=103
M2866 3950 WL_50 4052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=149710 $D=103
M2867 4054 WL_51 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=150200 $D=103
M2868 3950 WL_52 4056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=153110 $D=103
M2869 4058 WL_53 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=153600 $D=103
M2870 3950 WL_54 4060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=156510 $D=103
M2871 4062 WL_55 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=157000 $D=103
M2872 3950 WL_56 4064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=159910 $D=103
M2873 4066 WL_57 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=160400 $D=103
M2874 3950 WL_58 4068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=163310 $D=103
M2875 4070 WL_59 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=163800 $D=103
M2876 3950 WL_60 4072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=166710 $D=103
M2877 4074 WL_61 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=167200 $D=103
M2878 3950 WL_62 4076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=170110 $D=103
M2879 4078 WL_63 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=170600 $D=103
M2880 3950 WL_64 4080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=173510 $D=103
M2881 4082 WL_65 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=174000 $D=103
M2882 3950 WL_66 4084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=176910 $D=103
M2883 4086 WL_67 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=177400 $D=103
M2884 3950 WL_68 4088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=180310 $D=103
M2885 4090 WL_69 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=180800 $D=103
M2886 3950 WL_70 4092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=183710 $D=103
M2887 4094 WL_71 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=184200 $D=103
M2888 3950 WL_72 4096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=187110 $D=103
M2889 4098 WL_73 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=187600 $D=103
M2890 3950 WL_74 4100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=190510 $D=103
M2891 4102 WL_75 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=191000 $D=103
M2892 3950 WL_76 4104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=193910 $D=103
M2893 4106 WL_77 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=194400 $D=103
M2894 3950 WL_78 4108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=197310 $D=103
M2895 4110 WL_79 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=197800 $D=103
M2896 3950 WL_80 4112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=200710 $D=103
M2897 4114 WL_81 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=201200 $D=103
M2898 3950 WL_82 4116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=204110 $D=103
M2899 4118 WL_83 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=204600 $D=103
M2900 3950 WL_84 4120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=207510 $D=103
M2901 4122 WL_85 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=208000 $D=103
M2902 3950 WL_86 4124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=210910 $D=103
M2903 4126 WL_87 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=211400 $D=103
M2904 3950 WL_88 4128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=214310 $D=103
M2905 4130 WL_89 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=214800 $D=103
M2906 3950 WL_90 4132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=217710 $D=103
M2907 4134 WL_91 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=218200 $D=103
M2908 3950 WL_92 4136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=221110 $D=103
M2909 4138 WL_93 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=221600 $D=103
M2910 3950 WL_94 4140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=224510 $D=103
M2911 4142 WL_95 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=225000 $D=103
M2912 3950 WL_96 4144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=227910 $D=103
M2913 4146 WL_97 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=228400 $D=103
M2914 3950 WL_98 4148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=231310 $D=103
M2915 4150 WL_99 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=231800 $D=103
M2916 3950 WL_100 4152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=234710 $D=103
M2917 4154 WL_101 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=235200 $D=103
M2918 3950 WL_102 4156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=238110 $D=103
M2919 4158 WL_103 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=238600 $D=103
M2920 3950 WL_104 4160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=241510 $D=103
M2921 4162 WL_105 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=242000 $D=103
M2922 3950 WL_106 4164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=244910 $D=103
M2923 4166 WL_107 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=245400 $D=103
M2924 3950 WL_108 4168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=248310 $D=103
M2925 4170 WL_109 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=248800 $D=103
M2926 3950 WL_110 4172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=251710 $D=103
M2927 4174 WL_111 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=252200 $D=103
M2928 3950 WL_112 4176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=255110 $D=103
M2929 4178 WL_113 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=255600 $D=103
M2930 3950 WL_114 4180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=258510 $D=103
M2931 4182 WL_115 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=259000 $D=103
M2932 3950 WL_116 4184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=261910 $D=103
M2933 4186 WL_117 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=262400 $D=103
M2934 3950 WL_118 4188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=265310 $D=103
M2935 4190 WL_119 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=265800 $D=103
M2936 3950 WL_120 4192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=268710 $D=103
M2937 4194 WL_121 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=269200 $D=103
M2938 3950 WL_122 4196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=272110 $D=103
M2939 4198 WL_123 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=272600 $D=103
M2940 3950 WL_124 4200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=275510 $D=103
M2941 4202 WL_125 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=276000 $D=103
M2942 3950 WL_126 4204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=278910 $D=103
M2943 4206 WL_127 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=279400 $D=103
M2944 3950 WL_128 4208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=282310 $D=103
M2945 4210 WL_129 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=282800 $D=103
M2946 3950 WL_130 4212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=285710 $D=103
M2947 4214 WL_131 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=286200 $D=103
M2948 3950 WL_132 4216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=289110 $D=103
M2949 4218 WL_133 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=289600 $D=103
M2950 3950 WL_134 4220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=292510 $D=103
M2951 4222 WL_135 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=293000 $D=103
M2952 3950 WL_136 4224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=295910 $D=103
M2953 4226 WL_137 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=296400 $D=103
M2954 3950 WL_138 4228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=299310 $D=103
M2955 4230 WL_139 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=299800 $D=103
M2956 3950 WL_140 4232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=302710 $D=103
M2957 4234 WL_141 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=303200 $D=103
M2958 3950 WL_142 4236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=306110 $D=103
M2959 4238 WL_143 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=306600 $D=103
M2960 3950 WL_144 4240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=309510 $D=103
M2961 4242 WL_145 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=310000 $D=103
M2962 3950 WL_146 4244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=312910 $D=103
M2963 4246 WL_147 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=313400 $D=103
M2964 3950 WL_148 4248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=316310 $D=103
M2965 4250 WL_149 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=316800 $D=103
M2966 3950 WL_150 4252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=319710 $D=103
M2967 4254 WL_151 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=320200 $D=103
M2968 3950 WL_152 4256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=323110 $D=103
M2969 4258 WL_153 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=323600 $D=103
M2970 3950 WL_154 4260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=326510 $D=103
M2971 4262 WL_155 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=327000 $D=103
M2972 3950 WL_156 4264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=329910 $D=103
M2973 4266 WL_157 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=330400 $D=103
M2974 3950 WL_158 4268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=333310 $D=103
M2975 4270 WL_159 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=333800 $D=103
M2976 3950 WL_160 4272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=336710 $D=103
M2977 4274 WL_161 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=337200 $D=103
M2978 3950 WL_162 4276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=340110 $D=103
M2979 4278 WL_163 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=340600 $D=103
M2980 3950 WL_164 4280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=343510 $D=103
M2981 4282 WL_165 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=344000 $D=103
M2982 3950 WL_166 4284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=346910 $D=103
M2983 4286 WL_167 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=347400 $D=103
M2984 3950 WL_168 4288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=350310 $D=103
M2985 4290 WL_169 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=350800 $D=103
M2986 3950 WL_170 4292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=353710 $D=103
M2987 4294 WL_171 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=354200 $D=103
M2988 3950 WL_172 4296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=357110 $D=103
M2989 4298 WL_173 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=357600 $D=103
M2990 3950 WL_174 4300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=360510 $D=103
M2991 4302 WL_175 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=361000 $D=103
M2992 3950 WL_176 4304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=363910 $D=103
M2993 4306 WL_177 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=364400 $D=103
M2994 3950 WL_178 4308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=367310 $D=103
M2995 4310 WL_179 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=367800 $D=103
M2996 3950 WL_180 4312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=370710 $D=103
M2997 4314 WL_181 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=371200 $D=103
M2998 3950 WL_182 4316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=374110 $D=103
M2999 4318 WL_183 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=374600 $D=103
M3000 3950 WL_184 4320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=377510 $D=103
M3001 4322 WL_185 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=378000 $D=103
M3002 3950 WL_186 4324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=380910 $D=103
M3003 4326 WL_187 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=381400 $D=103
M3004 3950 WL_188 4328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=384310 $D=103
M3005 4330 WL_189 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=384800 $D=103
M3006 3950 WL_190 4332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=387710 $D=103
M3007 4334 WL_191 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=388200 $D=103
M3008 3950 WL_192 4336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=391110 $D=103
M3009 4338 WL_193 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=391600 $D=103
M3010 3950 WL_194 4340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=394510 $D=103
M3011 4342 WL_195 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=395000 $D=103
M3012 3950 WL_196 4344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=397910 $D=103
M3013 4346 WL_197 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=398400 $D=103
M3014 3950 WL_198 4348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=401310 $D=103
M3015 4350 WL_199 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=401800 $D=103
M3016 3950 WL_200 4352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=404710 $D=103
M3017 4354 WL_201 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=405200 $D=103
M3018 3950 WL_202 4356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=408110 $D=103
M3019 4358 WL_203 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=408600 $D=103
M3020 3950 WL_204 4360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=411510 $D=103
M3021 4362 WL_205 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=412000 $D=103
M3022 3950 WL_206 4364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=414910 $D=103
M3023 4366 WL_207 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=415400 $D=103
M3024 3950 WL_208 4368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=418310 $D=103
M3025 4370 WL_209 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=418800 $D=103
M3026 3950 WL_210 4372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=421710 $D=103
M3027 4374 WL_211 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=422200 $D=103
M3028 3950 WL_212 4376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=425110 $D=103
M3029 4378 WL_213 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=425600 $D=103
M3030 3950 WL_214 4380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=428510 $D=103
M3031 4382 WL_215 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=429000 $D=103
M3032 3950 WL_216 4384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=431910 $D=103
M3033 4386 WL_217 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=432400 $D=103
M3034 3950 WL_218 4388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=435310 $D=103
M3035 4390 WL_219 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=435800 $D=103
M3036 3950 WL_220 4392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=438710 $D=103
M3037 4394 WL_221 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=439200 $D=103
M3038 3950 WL_222 4396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=442110 $D=103
M3039 4398 WL_223 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=442600 $D=103
M3040 3950 WL_224 4400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=445510 $D=103
M3041 4402 WL_225 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=446000 $D=103
M3042 3950 WL_226 4404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=448910 $D=103
M3043 4406 WL_227 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=449400 $D=103
M3044 3950 WL_228 4408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=452310 $D=103
M3045 4410 WL_229 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=452800 $D=103
M3046 3950 WL_230 4412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=455710 $D=103
M3047 4414 WL_231 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=456200 $D=103
M3048 3950 WL_232 4416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=459110 $D=103
M3049 4418 WL_233 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=459600 $D=103
M3050 3950 WL_234 4420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=462510 $D=103
M3051 4422 WL_235 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=463000 $D=103
M3052 3950 WL_236 4424 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=465910 $D=103
M3053 4426 WL_237 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=466400 $D=103
M3054 3950 WL_238 4428 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=469310 $D=103
M3055 4430 WL_239 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=469800 $D=103
M3056 3950 WL_240 4432 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=472710 $D=103
M3057 4434 WL_241 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=473200 $D=103
M3058 3950 WL_242 4436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=476110 $D=103
M3059 4438 WL_243 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=476600 $D=103
M3060 3950 WL_244 4440 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=479510 $D=103
M3061 4442 WL_245 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=480000 $D=103
M3062 3950 WL_246 4444 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=482910 $D=103
M3063 4446 WL_247 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=483400 $D=103
M3064 3950 WL_248 4448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=486310 $D=103
M3065 4450 WL_249 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=486800 $D=103
M3066 3950 WL_250 4452 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=489710 $D=103
M3067 4454 WL_251 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=490200 $D=103
M3068 3950 WL_252 4456 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=493110 $D=103
M3069 4458 WL_253 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=493600 $D=103
M3070 3950 WL_254 4460 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=496510 $D=103
M3071 4462 WL_255 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=497000 $D=103
M3072 3949 WL_0 3951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=64710 $D=103
M3073 3953 WL_1 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=65200 $D=103
M3074 3949 WL_2 3955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=68110 $D=103
M3075 3957 WL_3 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=68600 $D=103
M3076 3949 WL_4 3959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=71510 $D=103
M3077 3961 WL_5 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=72000 $D=103
M3078 3949 WL_6 3963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=74910 $D=103
M3079 3965 WL_7 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=75400 $D=103
M3080 3949 WL_8 3967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=78310 $D=103
M3081 3969 WL_9 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=78800 $D=103
M3082 3949 WL_10 3971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=81710 $D=103
M3083 3973 WL_11 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=82200 $D=103
M3084 3949 WL_12 3975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=85110 $D=103
M3085 3977 WL_13 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=85600 $D=103
M3086 3949 WL_14 3979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=88510 $D=103
M3087 3981 WL_15 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=89000 $D=103
M3088 3949 WL_16 3983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=91910 $D=103
M3089 3985 WL_17 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=92400 $D=103
M3090 3949 WL_18 3987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=95310 $D=103
M3091 3989 WL_19 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=95800 $D=103
M3092 3949 WL_20 3991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=98710 $D=103
M3093 3993 WL_21 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=99200 $D=103
M3094 3949 WL_22 3995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=102110 $D=103
M3095 3997 WL_23 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=102600 $D=103
M3096 3949 WL_24 3999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=105510 $D=103
M3097 4001 WL_25 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=106000 $D=103
M3098 3949 WL_26 4003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=108910 $D=103
M3099 4005 WL_27 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=109400 $D=103
M3100 3949 WL_28 4007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=112310 $D=103
M3101 4009 WL_29 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=112800 $D=103
M3102 3949 WL_30 4011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=115710 $D=103
M3103 4013 WL_31 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=116200 $D=103
M3104 3949 WL_32 4015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=119110 $D=103
M3105 4017 WL_33 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=119600 $D=103
M3106 3949 WL_34 4019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=122510 $D=103
M3107 4021 WL_35 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=123000 $D=103
M3108 3949 WL_36 4023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=125910 $D=103
M3109 4025 WL_37 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=126400 $D=103
M3110 3949 WL_38 4027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=129310 $D=103
M3111 4029 WL_39 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=129800 $D=103
M3112 3949 WL_40 4031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=132710 $D=103
M3113 4033 WL_41 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=133200 $D=103
M3114 3949 WL_42 4035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=136110 $D=103
M3115 4037 WL_43 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=136600 $D=103
M3116 3949 WL_44 4039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=139510 $D=103
M3117 4041 WL_45 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=140000 $D=103
M3118 3949 WL_46 4043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=142910 $D=103
M3119 4045 WL_47 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=143400 $D=103
M3120 3949 WL_48 4047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=146310 $D=103
M3121 4049 WL_49 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=146800 $D=103
M3122 3949 WL_50 4051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=149710 $D=103
M3123 4053 WL_51 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=150200 $D=103
M3124 3949 WL_52 4055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=153110 $D=103
M3125 4057 WL_53 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=153600 $D=103
M3126 3949 WL_54 4059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=156510 $D=103
M3127 4061 WL_55 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=157000 $D=103
M3128 3949 WL_56 4063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=159910 $D=103
M3129 4065 WL_57 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=160400 $D=103
M3130 3949 WL_58 4067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=163310 $D=103
M3131 4069 WL_59 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=163800 $D=103
M3132 3949 WL_60 4071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=166710 $D=103
M3133 4073 WL_61 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=167200 $D=103
M3134 3949 WL_62 4075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=170110 $D=103
M3135 4077 WL_63 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=170600 $D=103
M3136 3949 WL_64 4079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=173510 $D=103
M3137 4081 WL_65 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=174000 $D=103
M3138 3949 WL_66 4083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=176910 $D=103
M3139 4085 WL_67 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=177400 $D=103
M3140 3949 WL_68 4087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=180310 $D=103
M3141 4089 WL_69 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=180800 $D=103
M3142 3949 WL_70 4091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=183710 $D=103
M3143 4093 WL_71 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=184200 $D=103
M3144 3949 WL_72 4095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=187110 $D=103
M3145 4097 WL_73 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=187600 $D=103
M3146 3949 WL_74 4099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=190510 $D=103
M3147 4101 WL_75 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=191000 $D=103
M3148 3949 WL_76 4103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=193910 $D=103
M3149 4105 WL_77 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=194400 $D=103
M3150 3949 WL_78 4107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=197310 $D=103
M3151 4109 WL_79 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=197800 $D=103
M3152 3949 WL_80 4111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=200710 $D=103
M3153 4113 WL_81 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=201200 $D=103
M3154 3949 WL_82 4115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=204110 $D=103
M3155 4117 WL_83 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=204600 $D=103
M3156 3949 WL_84 4119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=207510 $D=103
M3157 4121 WL_85 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=208000 $D=103
M3158 3949 WL_86 4123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=210910 $D=103
M3159 4125 WL_87 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=211400 $D=103
M3160 3949 WL_88 4127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=214310 $D=103
M3161 4129 WL_89 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=214800 $D=103
M3162 3949 WL_90 4131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=217710 $D=103
M3163 4133 WL_91 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=218200 $D=103
M3164 3949 WL_92 4135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=221110 $D=103
M3165 4137 WL_93 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=221600 $D=103
M3166 3949 WL_94 4139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=224510 $D=103
M3167 4141 WL_95 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=225000 $D=103
M3168 3949 WL_96 4143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=227910 $D=103
M3169 4145 WL_97 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=228400 $D=103
M3170 3949 WL_98 4147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=231310 $D=103
M3171 4149 WL_99 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=231800 $D=103
M3172 3949 WL_100 4151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=234710 $D=103
M3173 4153 WL_101 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=235200 $D=103
M3174 3949 WL_102 4155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=238110 $D=103
M3175 4157 WL_103 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=238600 $D=103
M3176 3949 WL_104 4159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=241510 $D=103
M3177 4161 WL_105 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=242000 $D=103
M3178 3949 WL_106 4163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=244910 $D=103
M3179 4165 WL_107 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=245400 $D=103
M3180 3949 WL_108 4167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=248310 $D=103
M3181 4169 WL_109 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=248800 $D=103
M3182 3949 WL_110 4171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=251710 $D=103
M3183 4173 WL_111 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=252200 $D=103
M3184 3949 WL_112 4175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=255110 $D=103
M3185 4177 WL_113 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=255600 $D=103
M3186 3949 WL_114 4179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=258510 $D=103
M3187 4181 WL_115 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=259000 $D=103
M3188 3949 WL_116 4183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=261910 $D=103
M3189 4185 WL_117 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=262400 $D=103
M3190 3949 WL_118 4187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=265310 $D=103
M3191 4189 WL_119 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=265800 $D=103
M3192 3949 WL_120 4191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=268710 $D=103
M3193 4193 WL_121 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=269200 $D=103
M3194 3949 WL_122 4195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=272110 $D=103
M3195 4197 WL_123 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=272600 $D=103
M3196 3949 WL_124 4199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=275510 $D=103
M3197 4201 WL_125 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=276000 $D=103
M3198 3949 WL_126 4203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=278910 $D=103
M3199 4205 WL_127 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=279400 $D=103
M3200 3949 WL_128 4207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=282310 $D=103
M3201 4209 WL_129 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=282800 $D=103
M3202 3949 WL_130 4211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=285710 $D=103
M3203 4213 WL_131 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=286200 $D=103
M3204 3949 WL_132 4215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=289110 $D=103
M3205 4217 WL_133 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=289600 $D=103
M3206 3949 WL_134 4219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=292510 $D=103
M3207 4221 WL_135 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=293000 $D=103
M3208 3949 WL_136 4223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=295910 $D=103
M3209 4225 WL_137 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=296400 $D=103
M3210 3949 WL_138 4227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=299310 $D=103
M3211 4229 WL_139 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=299800 $D=103
M3212 3949 WL_140 4231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=302710 $D=103
M3213 4233 WL_141 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=303200 $D=103
M3214 3949 WL_142 4235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=306110 $D=103
M3215 4237 WL_143 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=306600 $D=103
M3216 3949 WL_144 4239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=309510 $D=103
M3217 4241 WL_145 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=310000 $D=103
M3218 3949 WL_146 4243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=312910 $D=103
M3219 4245 WL_147 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=313400 $D=103
M3220 3949 WL_148 4247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=316310 $D=103
M3221 4249 WL_149 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=316800 $D=103
M3222 3949 WL_150 4251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=319710 $D=103
M3223 4253 WL_151 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=320200 $D=103
M3224 3949 WL_152 4255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=323110 $D=103
M3225 4257 WL_153 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=323600 $D=103
M3226 3949 WL_154 4259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=326510 $D=103
M3227 4261 WL_155 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=327000 $D=103
M3228 3949 WL_156 4263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=329910 $D=103
M3229 4265 WL_157 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=330400 $D=103
M3230 3949 WL_158 4267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=333310 $D=103
M3231 4269 WL_159 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=333800 $D=103
M3232 3949 WL_160 4271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=336710 $D=103
M3233 4273 WL_161 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=337200 $D=103
M3234 3949 WL_162 4275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=340110 $D=103
M3235 4277 WL_163 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=340600 $D=103
M3236 3949 WL_164 4279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=343510 $D=103
M3237 4281 WL_165 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=344000 $D=103
M3238 3949 WL_166 4283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=346910 $D=103
M3239 4285 WL_167 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=347400 $D=103
M3240 3949 WL_168 4287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=350310 $D=103
M3241 4289 WL_169 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=350800 $D=103
M3242 3949 WL_170 4291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=353710 $D=103
M3243 4293 WL_171 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=354200 $D=103
M3244 3949 WL_172 4295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=357110 $D=103
M3245 4297 WL_173 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=357600 $D=103
M3246 3949 WL_174 4299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=360510 $D=103
M3247 4301 WL_175 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=361000 $D=103
M3248 3949 WL_176 4303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=363910 $D=103
M3249 4305 WL_177 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=364400 $D=103
M3250 3949 WL_178 4307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=367310 $D=103
M3251 4309 WL_179 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=367800 $D=103
M3252 3949 WL_180 4311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=370710 $D=103
M3253 4313 WL_181 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=371200 $D=103
M3254 3949 WL_182 4315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=374110 $D=103
M3255 4317 WL_183 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=374600 $D=103
M3256 3949 WL_184 4319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=377510 $D=103
M3257 4321 WL_185 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=378000 $D=103
M3258 3949 WL_186 4323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=380910 $D=103
M3259 4325 WL_187 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=381400 $D=103
M3260 3949 WL_188 4327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=384310 $D=103
M3261 4329 WL_189 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=384800 $D=103
M3262 3949 WL_190 4331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=387710 $D=103
M3263 4333 WL_191 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=388200 $D=103
M3264 3949 WL_192 4335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=391110 $D=103
M3265 4337 WL_193 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=391600 $D=103
M3266 3949 WL_194 4339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=394510 $D=103
M3267 4341 WL_195 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=395000 $D=103
M3268 3949 WL_196 4343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=397910 $D=103
M3269 4345 WL_197 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=398400 $D=103
M3270 3949 WL_198 4347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=401310 $D=103
M3271 4349 WL_199 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=401800 $D=103
M3272 3949 WL_200 4351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=404710 $D=103
M3273 4353 WL_201 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=405200 $D=103
M3274 3949 WL_202 4355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=408110 $D=103
M3275 4357 WL_203 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=408600 $D=103
M3276 3949 WL_204 4359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=411510 $D=103
M3277 4361 WL_205 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=412000 $D=103
M3278 3949 WL_206 4363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=414910 $D=103
M3279 4365 WL_207 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=415400 $D=103
M3280 3949 WL_208 4367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=418310 $D=103
M3281 4369 WL_209 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=418800 $D=103
M3282 3949 WL_210 4371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=421710 $D=103
M3283 4373 WL_211 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=422200 $D=103
M3284 3949 WL_212 4375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=425110 $D=103
M3285 4377 WL_213 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=425600 $D=103
M3286 3949 WL_214 4379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=428510 $D=103
M3287 4381 WL_215 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=429000 $D=103
M3288 3949 WL_216 4383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=431910 $D=103
M3289 4385 WL_217 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=432400 $D=103
M3290 3949 WL_218 4387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=435310 $D=103
M3291 4389 WL_219 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=435800 $D=103
M3292 3949 WL_220 4391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=438710 $D=103
M3293 4393 WL_221 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=439200 $D=103
M3294 3949 WL_222 4395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=442110 $D=103
M3295 4397 WL_223 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=442600 $D=103
M3296 3949 WL_224 4399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=445510 $D=103
M3297 4401 WL_225 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=446000 $D=103
M3298 3949 WL_226 4403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=448910 $D=103
M3299 4405 WL_227 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=449400 $D=103
M3300 3949 WL_228 4407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=452310 $D=103
M3301 4409 WL_229 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=452800 $D=103
M3302 3949 WL_230 4411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=455710 $D=103
M3303 4413 WL_231 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=456200 $D=103
M3304 3949 WL_232 4415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=459110 $D=103
M3305 4417 WL_233 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=459600 $D=103
M3306 3949 WL_234 4419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=462510 $D=103
M3307 4421 WL_235 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=463000 $D=103
M3308 3949 WL_236 4423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=465910 $D=103
M3309 4425 WL_237 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=466400 $D=103
M3310 3949 WL_238 4427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=469310 $D=103
M3311 4429 WL_239 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=469800 $D=103
M3312 3949 WL_240 4431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=472710 $D=103
M3313 4433 WL_241 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=473200 $D=103
M3314 3949 WL_242 4435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=476110 $D=103
M3315 4437 WL_243 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=476600 $D=103
M3316 3949 WL_244 4439 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=479510 $D=103
M3317 4441 WL_245 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=480000 $D=103
M3318 3949 WL_246 4443 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=482910 $D=103
M3319 4445 WL_247 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=483400 $D=103
M3320 3949 WL_248 4447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=486310 $D=103
M3321 4449 WL_249 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=486800 $D=103
M3322 3949 WL_250 4451 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=489710 $D=103
M3323 4453 WL_251 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=490200 $D=103
M3324 3949 WL_252 4455 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=493110 $D=103
M3325 4457 WL_253 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=493600 $D=103
M3326 3949 WL_254 4459 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=496510 $D=103
M3327 4461 WL_255 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=497000 $D=103
M3328 608 WL_0 4463 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=64710 $D=103
M3329 4464 WL_1 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=65200 $D=103
M3330 608 WL_2 4465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=68110 $D=103
M3331 4466 WL_3 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=68600 $D=103
M3332 608 WL_4 4467 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=71510 $D=103
M3333 4468 WL_5 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=72000 $D=103
M3334 608 WL_6 4469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=74910 $D=103
M3335 4470 WL_7 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=75400 $D=103
M3336 608 WL_8 4471 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=78310 $D=103
M3337 4472 WL_9 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=78800 $D=103
M3338 608 WL_10 4473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=81710 $D=103
M3339 4474 WL_11 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=82200 $D=103
M3340 608 WL_12 4475 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=85110 $D=103
M3341 4476 WL_13 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=85600 $D=103
M3342 608 WL_14 4477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=88510 $D=103
M3343 4478 WL_15 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=89000 $D=103
M3344 608 WL_16 4479 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=91910 $D=103
M3345 4480 WL_17 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=92400 $D=103
M3346 608 WL_18 4481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=95310 $D=103
M3347 4482 WL_19 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=95800 $D=103
M3348 608 WL_20 4483 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=98710 $D=103
M3349 4484 WL_21 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=99200 $D=103
M3350 608 WL_22 4485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=102110 $D=103
M3351 4486 WL_23 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=102600 $D=103
M3352 608 WL_24 4487 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=105510 $D=103
M3353 4488 WL_25 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=106000 $D=103
M3354 608 WL_26 4489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=108910 $D=103
M3355 4490 WL_27 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=109400 $D=103
M3356 608 WL_28 4491 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=112310 $D=103
M3357 4492 WL_29 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=112800 $D=103
M3358 608 WL_30 4493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=115710 $D=103
M3359 4494 WL_31 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=116200 $D=103
M3360 608 WL_32 4495 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=119110 $D=103
M3361 4496 WL_33 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=119600 $D=103
M3362 608 WL_34 4497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=122510 $D=103
M3363 4498 WL_35 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=123000 $D=103
M3364 608 WL_36 4499 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=125910 $D=103
M3365 4500 WL_37 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=126400 $D=103
M3366 608 WL_38 4501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=129310 $D=103
M3367 4502 WL_39 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=129800 $D=103
M3368 608 WL_40 4503 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=132710 $D=103
M3369 4504 WL_41 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=133200 $D=103
M3370 608 WL_42 4505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=136110 $D=103
M3371 4506 WL_43 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=136600 $D=103
M3372 608 WL_44 4507 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=139510 $D=103
M3373 4508 WL_45 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=140000 $D=103
M3374 608 WL_46 4509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=142910 $D=103
M3375 4510 WL_47 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=143400 $D=103
M3376 608 WL_48 4511 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=146310 $D=103
M3377 4512 WL_49 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=146800 $D=103
M3378 608 WL_50 4513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=149710 $D=103
M3379 4514 WL_51 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=150200 $D=103
M3380 608 WL_52 4515 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=153110 $D=103
M3381 4516 WL_53 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=153600 $D=103
M3382 608 WL_54 4517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=156510 $D=103
M3383 4518 WL_55 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=157000 $D=103
M3384 608 WL_56 4519 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=159910 $D=103
M3385 4520 WL_57 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=160400 $D=103
M3386 608 WL_58 4521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=163310 $D=103
M3387 4522 WL_59 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=163800 $D=103
M3388 608 WL_60 4523 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=166710 $D=103
M3389 4524 WL_61 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=167200 $D=103
M3390 608 WL_62 4525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=170110 $D=103
M3391 4526 WL_63 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=170600 $D=103
M3392 608 WL_64 4527 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=173510 $D=103
M3393 4528 WL_65 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=174000 $D=103
M3394 608 WL_66 4529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=176910 $D=103
M3395 4530 WL_67 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=177400 $D=103
M3396 608 WL_68 4531 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=180310 $D=103
M3397 4532 WL_69 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=180800 $D=103
M3398 608 WL_70 4533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=183710 $D=103
M3399 4534 WL_71 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=184200 $D=103
M3400 608 WL_72 4535 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=187110 $D=103
M3401 4536 WL_73 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=187600 $D=103
M3402 608 WL_74 4537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=190510 $D=103
M3403 4538 WL_75 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=191000 $D=103
M3404 608 WL_76 4539 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=193910 $D=103
M3405 4540 WL_77 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=194400 $D=103
M3406 608 WL_78 4541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=197310 $D=103
M3407 4542 WL_79 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=197800 $D=103
M3408 608 WL_80 4543 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=200710 $D=103
M3409 4544 WL_81 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=201200 $D=103
M3410 608 WL_82 4545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=204110 $D=103
M3411 4546 WL_83 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=204600 $D=103
M3412 608 WL_84 4547 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=207510 $D=103
M3413 4548 WL_85 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=208000 $D=103
M3414 608 WL_86 4549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=210910 $D=103
M3415 4550 WL_87 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=211400 $D=103
M3416 608 WL_88 4551 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=214310 $D=103
M3417 4552 WL_89 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=214800 $D=103
M3418 608 WL_90 4553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=217710 $D=103
M3419 4554 WL_91 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=218200 $D=103
M3420 608 WL_92 4555 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=221110 $D=103
M3421 4556 WL_93 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=221600 $D=103
M3422 608 WL_94 4557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=224510 $D=103
M3423 4558 WL_95 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=225000 $D=103
M3424 608 WL_96 4559 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=227910 $D=103
M3425 4560 WL_97 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=228400 $D=103
M3426 608 WL_98 4561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=231310 $D=103
M3427 4562 WL_99 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=231800 $D=103
M3428 608 WL_100 4563 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=234710 $D=103
M3429 4564 WL_101 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=235200 $D=103
M3430 608 WL_102 4565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=238110 $D=103
M3431 4566 WL_103 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=238600 $D=103
M3432 608 WL_104 4567 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=241510 $D=103
M3433 4568 WL_105 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=242000 $D=103
M3434 608 WL_106 4569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=244910 $D=103
M3435 4570 WL_107 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=245400 $D=103
M3436 608 WL_108 4571 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=248310 $D=103
M3437 4572 WL_109 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=248800 $D=103
M3438 608 WL_110 4573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=251710 $D=103
M3439 4574 WL_111 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=252200 $D=103
M3440 608 WL_112 4575 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=255110 $D=103
M3441 4576 WL_113 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=255600 $D=103
M3442 608 WL_114 4577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=258510 $D=103
M3443 4578 WL_115 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=259000 $D=103
M3444 608 WL_116 4579 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=261910 $D=103
M3445 4580 WL_117 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=262400 $D=103
M3446 608 WL_118 4581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=265310 $D=103
M3447 4582 WL_119 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=265800 $D=103
M3448 608 WL_120 4583 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=268710 $D=103
M3449 4584 WL_121 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=269200 $D=103
M3450 608 WL_122 4585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=272110 $D=103
M3451 4586 WL_123 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=272600 $D=103
M3452 608 WL_124 4587 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=275510 $D=103
M3453 4588 WL_125 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=276000 $D=103
M3454 608 WL_126 4589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=278910 $D=103
M3455 4590 WL_127 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=279400 $D=103
M3456 608 WL_128 4591 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=282310 $D=103
M3457 4592 WL_129 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=282800 $D=103
M3458 608 WL_130 4593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=285710 $D=103
M3459 4594 WL_131 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=286200 $D=103
M3460 608 WL_132 4595 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=289110 $D=103
M3461 4596 WL_133 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=289600 $D=103
M3462 608 WL_134 4597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=292510 $D=103
M3463 4598 WL_135 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=293000 $D=103
M3464 608 WL_136 4599 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=295910 $D=103
M3465 4600 WL_137 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=296400 $D=103
M3466 608 WL_138 4601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=299310 $D=103
M3467 4602 WL_139 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=299800 $D=103
M3468 608 WL_140 4603 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=302710 $D=103
M3469 4604 WL_141 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=303200 $D=103
M3470 608 WL_142 4605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=306110 $D=103
M3471 4606 WL_143 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=306600 $D=103
M3472 608 WL_144 4607 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=309510 $D=103
M3473 4608 WL_145 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=310000 $D=103
M3474 608 WL_146 4609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=312910 $D=103
M3475 4610 WL_147 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=313400 $D=103
M3476 608 WL_148 4611 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=316310 $D=103
M3477 4612 WL_149 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=316800 $D=103
M3478 608 WL_150 4613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=319710 $D=103
M3479 4614 WL_151 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=320200 $D=103
M3480 608 WL_152 4615 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=323110 $D=103
M3481 4616 WL_153 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=323600 $D=103
M3482 608 WL_154 4617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=326510 $D=103
M3483 4618 WL_155 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=327000 $D=103
M3484 608 WL_156 4619 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=329910 $D=103
M3485 4620 WL_157 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=330400 $D=103
M3486 608 WL_158 4621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=333310 $D=103
M3487 4622 WL_159 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=333800 $D=103
M3488 608 WL_160 4623 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=336710 $D=103
M3489 4624 WL_161 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=337200 $D=103
M3490 608 WL_162 4625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=340110 $D=103
M3491 4626 WL_163 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=340600 $D=103
M3492 608 WL_164 4627 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=343510 $D=103
M3493 4628 WL_165 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=344000 $D=103
M3494 608 WL_166 4629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=346910 $D=103
M3495 4630 WL_167 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=347400 $D=103
M3496 608 WL_168 4631 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=350310 $D=103
M3497 4632 WL_169 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=350800 $D=103
M3498 608 WL_170 4633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=353710 $D=103
M3499 4634 WL_171 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=354200 $D=103
M3500 608 WL_172 4635 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=357110 $D=103
M3501 4636 WL_173 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=357600 $D=103
M3502 608 WL_174 4637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=360510 $D=103
M3503 4638 WL_175 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=361000 $D=103
M3504 608 WL_176 4639 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=363910 $D=103
M3505 4640 WL_177 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=364400 $D=103
M3506 608 WL_178 4641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=367310 $D=103
M3507 4642 WL_179 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=367800 $D=103
M3508 608 WL_180 4643 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=370710 $D=103
M3509 4644 WL_181 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=371200 $D=103
M3510 608 WL_182 4645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=374110 $D=103
M3511 4646 WL_183 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=374600 $D=103
M3512 608 WL_184 4647 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=377510 $D=103
M3513 4648 WL_185 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=378000 $D=103
M3514 608 WL_186 4649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=380910 $D=103
M3515 4650 WL_187 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=381400 $D=103
M3516 608 WL_188 4651 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=384310 $D=103
M3517 4652 WL_189 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=384800 $D=103
M3518 608 WL_190 4653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=387710 $D=103
M3519 4654 WL_191 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=388200 $D=103
M3520 608 WL_192 4655 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=391110 $D=103
M3521 4656 WL_193 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=391600 $D=103
M3522 608 WL_194 4657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=394510 $D=103
M3523 4658 WL_195 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=395000 $D=103
M3524 608 WL_196 4659 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=397910 $D=103
M3525 4660 WL_197 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=398400 $D=103
M3526 608 WL_198 4661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=401310 $D=103
M3527 4662 WL_199 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=401800 $D=103
M3528 608 WL_200 4663 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=404710 $D=103
M3529 4664 WL_201 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=405200 $D=103
M3530 608 WL_202 4665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=408110 $D=103
M3531 4666 WL_203 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=408600 $D=103
M3532 608 WL_204 4667 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=411510 $D=103
M3533 4668 WL_205 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=412000 $D=103
M3534 608 WL_206 4669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=414910 $D=103
M3535 4670 WL_207 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=415400 $D=103
M3536 608 WL_208 4671 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=418310 $D=103
M3537 4672 WL_209 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=418800 $D=103
M3538 608 WL_210 4673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=421710 $D=103
M3539 4674 WL_211 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=422200 $D=103
M3540 608 WL_212 4675 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=425110 $D=103
M3541 4676 WL_213 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=425600 $D=103
M3542 608 WL_214 4677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=428510 $D=103
M3543 4678 WL_215 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=429000 $D=103
M3544 608 WL_216 4679 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=431910 $D=103
M3545 4680 WL_217 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=432400 $D=103
M3546 608 WL_218 4681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=435310 $D=103
M3547 4682 WL_219 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=435800 $D=103
M3548 608 WL_220 4683 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=438710 $D=103
M3549 4684 WL_221 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=439200 $D=103
M3550 608 WL_222 4685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=442110 $D=103
M3551 4686 WL_223 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=442600 $D=103
M3552 608 WL_224 4687 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=445510 $D=103
M3553 4688 WL_225 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=446000 $D=103
M3554 608 WL_226 4689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=448910 $D=103
M3555 4690 WL_227 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=449400 $D=103
M3556 608 WL_228 4691 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=452310 $D=103
M3557 4692 WL_229 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=452800 $D=103
M3558 608 WL_230 4693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=455710 $D=103
M3559 4694 WL_231 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=456200 $D=103
M3560 608 WL_232 4695 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=459110 $D=103
M3561 4696 WL_233 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=459600 $D=103
M3562 608 WL_234 4697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=462510 $D=103
M3563 4698 WL_235 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=463000 $D=103
M3564 608 WL_236 4699 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=465910 $D=103
M3565 4700 WL_237 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=466400 $D=103
M3566 608 WL_238 4701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=469310 $D=103
M3567 4702 WL_239 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=469800 $D=103
M3568 608 WL_240 4703 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=472710 $D=103
M3569 4704 WL_241 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=473200 $D=103
M3570 608 WL_242 4705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=476110 $D=103
M3571 4706 WL_243 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=476600 $D=103
M3572 608 WL_244 4707 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=479510 $D=103
M3573 4708 WL_245 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=480000 $D=103
M3574 608 WL_246 4709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=482910 $D=103
M3575 4710 WL_247 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=483400 $D=103
M3576 608 WL_248 4711 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=486310 $D=103
M3577 4712 WL_249 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=486800 $D=103
M3578 608 WL_250 4713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=489710 $D=103
M3579 4714 WL_251 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=490200 $D=103
M3580 608 WL_252 4715 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=493110 $D=103
M3581 4716 WL_253 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=493600 $D=103
M3582 608 WL_254 4717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=496510 $D=103
M3583 4718 WL_255 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=497000 $D=103
X3584 Q_0 VDD D_0 VSS GTP_0 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14
+ WL_15 WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34
+ WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54
+ WL_55 WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74
+ WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94
+ WL_95 WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114
+ WL_115 WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134
+ WL_135 WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154
+ WL_155 WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174
+ WL_175 WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194
+ WL_195 WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214
+ WL_215 WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234
+ WL_235 WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254
+ WL_255 WE OE_ 545 546 547 548 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 1122 609 1123
+ 610 1124 611 1125 612 1126 613 1127 614 1128 615 1129 616 1130 617 1131 618 1132 619 1133
+ 620 1134 621 1135 622 1136 623 1137 624 1138 625 1139 626 1140 627 1141 628 1142 629 1143
+ 630 1144 631 1145 632 1146 633 1147 634 1148 635 1149 636 1150 637 1151 638 1152 639 1153
+ 640 1154 641 1155 642 1156 643 1157 644 1158 645 1159 646 1160 647 1161 648 1162 649 1163
+ 650 1164 651 1165 652 1166 653 1167 654 1168 655 1169 656 1170 657 1171 658 1172 659 1173
+ 660 1174 661 1175 662 1176 663 1177 664 1178 665 1179 666 1180 667 1181 668 1182 669 1183
+ 670 1184 671 1185 672 1186 673 1187 674 1188 675 1189 676 1190 677 1191 678 1192 679 1193
+ 680 1194 681 1195 682 1196 683 1197 684 1198 685 1199 686 1200 687 1201 688 1202 689 1203
+ 690 1204 691 1205 692 1206 693 1207 694 1208 695 1209 696 1210 697 1211 698 1212 699 1213
+ 700 1214 701 1215 702 1216 703 1217 704 1218 705 1219 706 1220 707 1221 708 1222 709 1223
+ 710 1224 711 1225 712 1226 713 1227 714 1228 715 1229 716 1230 717 1231 718 1232 719 1233
+ 720 1234 721 1235 722 1236 723 1237 724 1238 725 1239 726 1240 727 1241 728 1242 729 1243
+ 730 1244 731 1245 732 1246 733 1247 734 1248 735 1249 736 1250 737 1251 738 1252 739 1253
+ 740 1254 741 1255 742 1256 743 1257 744 1258 745 1259 746 1260 747 1261 748 1262 749 1263
+ 750 1264 751 1265 752 1266 753 1267 754 1268 755 1269 756 1270 757 1271 758 1272 759 1273
+ 760 1274 761 1275 762 1276 763 1277 764 1278 765 1279 766 1280 767 1281 768 1282 769 1283
+ 770 1284 771 1285 772 1286 773 1287 774 1288 775 1289 776 1290 777 1291 778 1292 779 1293
+ 780 1294 781 1295 782 1296 783 1297 784 1298 785 1299 786 1300 787 1301 788 1302 789 1303
+ 790 1304 791 1305 792 1306 793 1307 794 1308 795 1309 796 1310 797 1311 798 1312 799 1313
+ 800 1314 801 1315 802 1316 803 1317 804 1318 805 1319 806 1320 807 1321 808 1322 809 1323
+ 810 1324 811 1325 812 1326 813 1327 814 1328 815 1329 816 1330 817 1331 818 1332 819 1333
+ 820 1334 821 1335 822 1336 823 1337 824 1338 825 1339 826 1340 827 1341 828 1342 829 1343
+ 830 1344 831 1345 832 1346 833 1347 834 1348 835 1349 836 1350 837 1351 838 1352 839 1353
+ 840 1354 841 1355 842 1356 843 1357 844 1358 845 1359 846 1360 847 1361 848 1362 849 1363
+ 850 1364 851 1365 852 1366 853 1367 854 1368 855 1369 856 1370 857 1371 858 1372 859 1373
+ 860 1374 861 1375 862 1376 863 1377 864 1378 865
+ ICV_137 $T=0 0 0 0 $X=-1000 $Y=-1000
X3585 Q_1 VDD D_1 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 549 550 551 552 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 1379 1380 1381
+ 1382 1383 1384 1385 1386 1387 1388 1389 1390 1391 1392 1393 1394 1395 1396 1397 1398 1399 1400 1401
+ 1402 1403 1404 1405 1406 1407 1408 1409 1410 1411 1412 1413 1414 1415 1416 1417 1418 1419 1420 1421
+ 1422 1423 1424 1425 1426 1427 1428 1429 1430 1431 1432 1433 1434 1435 1436 1437 1438 1439 1440 1441
+ 1442 1443 1444 1445 1446 1447 1448 1449 1450 1451 1452 1453 1454 1455 1456 1457 1458 1459 1460 1461
+ 1462 1463 1464 1465 1466 1467 1468 1469 1470 1471 1472 1473 1474 1475 1476 1477 1478 1479 1480 1481
+ 1482 1483 1484 1485 1486 1487 1488 1489 1490 1491 1492 1493 1494 1495 1496 1497 1498 1499 1500 1501
+ 1502 1503 1504 1505 1506 1507 1508 1509 1510 1511 1512 1513 1514 1515 1516 1517 1518 1519 1520 1521
+ 1522 1523 1524 1525 1526 1527 1528 1529 1530 1531 1532 1533 1534 1535 1536 1537 1538 1539 1540 1541
+ 1542 1543 1544 1545 1546 1547 1548 1549 1550 1551 1552 1553 1554 1555 1556 1557 1558 1559 1560 1561
+ 1562 1563 1564 1565 1566 1567 1568 1569 1570 1571 1572 1573 1574 1575 1576 1577 1578 1579 1580 1581
+ 1582 1583 1584 1585 1586 1587 1588 1589 1590 1591 1592 1593 1594 1595 1596 1597 1598 1599 1600 1601
+ 1602 1603 1604 1605 1606 1607 1608 1609 1610 1611 1612 1613 1614 1615 1616 1617 1618 1619 1620 1621
+ 1622 1623 1624 1625 1626 1627 1628 1629 1630 1631 1632 1633 1634 1635 1636 1637 1638 1639 1640 1641
+ 1642 1643 1644 1645 1646 1647 1648 1649 1650 1651 1652 1653 1654 1655 1656 1657 1658 1659 1660 1661
+ 1662 1663 1664 1665 1666 1667 1668 1669 1670 1671 1672 1673 1674 1675 1676 1677 1678 1679 1680 1681
+ 1682 1683 1684 1685 1686 1687 1688 1689 1690 1691 1692 1693 1694 1695 1696 1697 1698 1699 1700 1701
+ 1702 1703 1704 1705 1706 1707 1708 1709 1710 1711 1712 1713 1714 1715 1716 1717 1718 1719 1720 1721
+ 1722 1723 1724 1725 1726 1727 1728 1729 1730 1731 1732 1733 1734 1735 1736 1737 1738 1739 1740 1741
+ 1742 1743 1744 1745 1746 1747 1748 1749 1750 1751 1752 1753 1754 1755 1756 1757 1758 1759 1760 1761
+ 1762 1763 1764 1765 1766 1767 1768 1769 1770 1771 1772 1773 1774 1775 1776 1777 1778 1779 1780 1781
+ 1782 1783 1784 1785 1786 1787 1788 1789 1790 1791 1792 1793 1794 1795 1796 1797 1798 1799 1800 1801
+ 1802 1803 1804 1805 1806 1807 1808 1809 1810 1811 1812 1813 1814 1815 1816 1817 1818 1819 1820 1821
+ 1822 1823 1824 1825 1826 1827 1828 1829 1830 1831 1832 1833 1834 1835 1836 1837 1838 1839 1840 1841
+ 1842 1843 1844 1845 1846 1847 1848 1849 1850 1851 1852 1853 1854 1855 1856 1857 1858 1859 1860 1861
+ 1862 1863 1864 1865 1866 1867 1868 1869 1870 1871 1872 1873 1874 1875 1876 1877 1878 1879 1880 1881
+ 1882 1883 1884 1885 1886 1887 1888 1889 1890 1891 1892
+ ICV_132 $T=38400 0 1 180 $X=18200 $Y=-1000
X3586 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_142 $T=0 0 0 90 $X=37400 $Y=62320
X3587 Q_2 VDD D_2 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 553 554 555 556 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 1893 1894 1895
+ 1896 1897 1898 1899 1900 1901 1902 1903 1904 1905 1906 1907 1908 1909 1910 1911 1912 1913 1914 1915
+ 1916 1917 1918 1919 1920 1921 1922 1923 1924 1925 1926 1927 1928 1929 1930 1931 1932 1933 1934 1935
+ 1936 1937 1938 1939 1940 1941 1942 1943 1944 1945 1946 1947 1948 1949 1950 1951 1952 1953 1954 1955
+ 1956 1957 1958 1959 1960 1961 1962 1963 1964 1965 1966 1967 1968 1969 1970 1971 1972 1973 1974 1975
+ 1976 1977 1978 1979 1980 1981 1982 1983 1984 1985 1986 1987 1988 1989 1990 1991 1992 1993 1994 1995
+ 1996 1997 1998 1999 2000 2001 2002 2003 2004 2005 2006 2007 2008 2009 2010 2011 2012 2013 2014 2015
+ 2016 2017 2018 2019 2020 2021 2022 2023 2024 2025 2026 2027 2028 2029 2030 2031 2032 2033 2034 2035
+ 2036 2037 2038 2039 2040 2041 2042 2043 2044 2045 2046 2047 2048 2049 2050 2051 2052 2053 2054 2055
+ 2056 2057 2058 2059 2060 2061 2062 2063 2064 2065 2066 2067 2068 2069 2070 2071 2072 2073 2074 2075
+ 2076 2077 2078 2079 2080 2081 2082 2083 2084 2085 2086 2087 2088 2089 2090 2091 2092 2093 2094 2095
+ 2096 2097 2098 2099 2100 2101 2102 2103 2104 2105 2106 2107 2108 2109 2110 2111 2112 2113 2114 2115
+ 2116 2117 2118 2119 2120 2121 2122 2123 2124 2125 2126 2127 2128 2129 2130 2131 2132 2133 2134 2135
+ 2136 2137 2138 2139 2140 2141 2142 2143 2144 2145 2146 2147 2148 2149 2150 2151 2152 2153 2154 2155
+ 2156 2157 2158 2159 2160 2161 2162 2163 2164 2165 2166 2167 2168 2169 2170 2171 2172 2173 2174 2175
+ 2176 2177 2178 2179 2180 2181 2182 2183 2184 2185 2186 2187 2188 2189 2190 2191 2192 2193 2194 2195
+ 2196 2197 2198 2199 2200 2201 2202 2203 2204 2205 2206 2207 2208 2209 2210 2211 2212 2213 2214 2215
+ 2216 2217 2218 2219 2220 2221 2222 2223 2224 2225 2226 2227 2228 2229 2230 2231 2232 2233 2234 2235
+ 2236 2237 2238 2239 2240 2241 2242 2243 2244 2245 2246 2247 2248 2249 2250 2251 2252 2253 2254 2255
+ 2256 2257 2258 2259 2260 2261 2262 2263 2264 2265 2266 2267 2268 2269 2270 2271 2272 2273 2274 2275
+ 2276 2277 2278 2279 2280 2281 2282 2283 2284 2285 2286 2287 2288 2289 2290 2291 2292 2293 2294 2295
+ 2296 2297 2298 2299 2300 2301 2302 2303 2304 2305 2306 2307 2308 2309 2310 2311 2312 2313 2314 2315
+ 2316 2317 2318 2319 2320 2321 2322 2323 2324 2325 2326 2327 2328 2329 2330 2331 2332 2333 2334 2335
+ 2336 2337 2338 2339 2340 2341 2342 2343 2344 2345 2346 2347 2348 2349 2350 2351 2352 2353 2354 2355
+ 2356 2357 2358 2359 2360 2361 2362 2363 2364 2365 2366 2367 2368 2369 2370 2371 2372 2373 2374 2375
+ 2376 2377 2378 2379 2380 2381 2382 2383 2384 2385 2386 2387 2388 2389 2390 2391 2392 2393 2394 2395
+ 2396 2397 2398 2399 2400 2401 2402 2403 2404 2405 2406
+ ICV_127 $T=39600 0 0 0 $X=38600 $Y=-1000
X3588 Q_3 VDD D_3 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 557 558 559 560 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 2407 2408 2409
+ 2410 2411 2412 2413 2414 2415 2416 2417 2418 2419 2420 2421 2422 2423 2424 2425 2426 2427 2428 2429
+ 2430 2431 2432 2433 2434 2435 2436 2437 2438 2439 2440 2441 2442 2443 2444 2445 2446 2447 2448 2449
+ 2450 2451 2452 2453 2454 2455 2456 2457 2458 2459 2460 2461 2462 2463 2464 2465 2466 2467 2468 2469
+ 2470 2471 2472 2473 2474 2475 2476 2477 2478 2479 2480 2481 2482 2483 2484 2485 2486 2487 2488 2489
+ 2490 2491 2492 2493 2494 2495 2496 2497 2498 2499 2500 2501 2502 2503 2504 2505 2506 2507 2508 2509
+ 2510 2511 2512 2513 2514 2515 2516 2517 2518 2519 2520 2521 2522 2523 2524 2525 2526 2527 2528 2529
+ 2530 2531 2532 2533 2534 2535 2536 2537 2538 2539 2540 2541 2542 2543 2544 2545 2546 2547 2548 2549
+ 2550 2551 2552 2553 2554 2555 2556 2557 2558 2559 2560 2561 2562 2563 2564 2565 2566 2567 2568 2569
+ 2570 2571 2572 2573 2574 2575 2576 2577 2578 2579 2580 2581 2582 2583 2584 2585 2586 2587 2588 2589
+ 2590 2591 2592 2593 2594 2595 2596 2597 2598 2599 2600 2601 2602 2603 2604 2605 2606 2607 2608 2609
+ 2610 2611 2612 2613 2614 2615 2616 2617 2618 2619 2620 2621 2622 2623 2624 2625 2626 2627 2628 2629
+ 2630 2631 2632 2633 2634 2635 2636 2637 2638 2639 2640 2641 2642 2643 2644 2645 2646 2647 2648 2649
+ 2650 2651 2652 2653 2654 2655 2656 2657 2658 2659 2660 2661 2662 2663 2664 2665 2666 2667 2668 2669
+ 2670 2671 2672 2673 2674 2675 2676 2677 2678 2679 2680 2681 2682 2683 2684 2685 2686 2687 2688 2689
+ 2690 2691 2692 2693 2694 2695 2696 2697 2698 2699 2700 2701 2702 2703 2704 2705 2706 2707 2708 2709
+ 2710 2711 2712 2713 2714 2715 2716 2717 2718 2719 2720 2721 2722 2723 2724 2725 2726 2727 2728 2729
+ 2730 2731 2732 2733 2734 2735 2736 2737 2738 2739 2740 2741 2742 2743 2744 2745 2746 2747 2748 2749
+ 2750 2751 2752 2753 2754 2755 2756 2757 2758 2759 2760 2761 2762 2763 2764 2765 2766 2767 2768 2769
+ 2770 2771 2772 2773 2774 2775 2776 2777 2778 2779 2780 2781 2782 2783 2784 2785 2786 2787 2788 2789
+ 2790 2791 2792 2793 2794 2795 2796 2797 2798 2799 2800 2801 2802 2803 2804 2805 2806 2807 2808 2809
+ 2810 2811 2812 2813 2814 2815 2816 2817 2818 2819 2820 2821 2822 2823 2824 2825 2826 2827 2828 2829
+ 2830 2831 2832 2833 2834 2835 2836 2837 2838 2839 2840 2841 2842 2843 2844 2845 2846 2847 2848 2849
+ 2850 2851 2852 2853 2854 2855 2856 2857 2858 2859 2860 2861 2862 2863 2864 2865 2866 2867 2868 2869
+ 2870 2871 2872 2873 2874 2875 2876 2877 2878 2879 2880 2881 2882 2883 2884 2885 2886 2887 2888 2889
+ 2890 2891 2892 2893 2894 2895 2896 2897 2898 2899 2900 2901 2902 2903 2904 2905 2906 2907 2908 2909
+ 2910 2911 2912 2913 2914 2915 2916 2917 2918 2919 2920
+ ICV_122 $T=78000 0 1 180 $X=57800 $Y=-1000
X3589 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_141 $T=0 0 0 90 $X=77000 $Y=62320
X3590 Q_4 VDD D_4 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 561 562 563 564 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 2921 2922 2923
+ 2924 2925 2926 2927 2928 2929 2930 2931 2932 2933 2934 2935 2936 2937 2938 2939 2940 2941 2942 2943
+ 2944 2945 2946 2947 2948 2949 2950 2951 2952 2953 2954 2955 2956 2957 2958 2959 2960 2961 2962 2963
+ 2964 2965 2966 2967 2968 2969 2970 2971 2972 2973 2974 2975 2976 2977 2978 2979 2980 2981 2982 2983
+ 2984 2985 2986 2987 2988 2989 2990 2991 2992 2993 2994 2995 2996 2997 2998 2999 3000 3001 3002 3003
+ 3004 3005 3006 3007 3008 3009 3010 3011 3012 3013 3014 3015 3016 3017 3018 3019 3020 3021 3022 3023
+ 3024 3025 3026 3027 3028 3029 3030 3031 3032 3033 3034 3035 3036 3037 3038 3039 3040 3041 3042 3043
+ 3044 3045 3046 3047 3048 3049 3050 3051 3052 3053 3054 3055 3056 3057 3058 3059 3060 3061 3062 3063
+ 3064 3065 3066 3067 3068 3069 3070 3071 3072 3073 3074 3075 3076 3077 3078 3079 3080 3081 3082 3083
+ 3084 3085 3086 3087 3088 3089 3090 3091 3092 3093 3094 3095 3096 3097 3098 3099 3100 3101 3102 3103
+ 3104 3105 3106 3107 3108 3109 3110 3111 3112 3113 3114 3115 3116 3117 3118 3119 3120 3121 3122 3123
+ 3124 3125 3126 3127 3128 3129 3130 3131 3132 3133 3134 3135 3136 3137 3138 3139 3140 3141 3142 3143
+ 3144 3145 3146 3147 3148 3149 3150 3151 3152 3153 3154 3155 3156 3157 3158 3159 3160 3161 3162 3163
+ 3164 3165 3166 3167 3168 3169 3170 3171 3172 3173 3174 3175 3176 3177 3178 3179 3180 3181 3182 3183
+ 3184 3185 3186 3187 3188 3189 3190 3191 3192 3193 3194 3195 3196 3197 3198 3199 3200 3201 3202 3203
+ 3204 3205 3206 3207 3208 3209 3210 3211 3212 3213 3214 3215 3216 3217 3218 3219 3220 3221 3222 3223
+ 3224 3225 3226 3227 3228 3229 3230 3231 3232 3233 3234 3235 3236 3237 3238 3239 3240 3241 3242 3243
+ 3244 3245 3246 3247 3248 3249 3250 3251 3252 3253 3254 3255 3256 3257 3258 3259 3260 3261 3262 3263
+ 3264 3265 3266 3267 3268 3269 3270 3271 3272 3273 3274 3275 3276 3277 3278 3279 3280 3281 3282 3283
+ 3284 3285 3286 3287 3288 3289 3290 3291 3292 3293 3294 3295 3296 3297 3298 3299 3300 3301 3302 3303
+ 3304 3305 3306 3307 3308 3309 3310 3311 3312 3313 3314 3315 3316 3317 3318 3319 3320 3321 3322 3323
+ 3324 3325 3326 3327 3328 3329 3330 3331 3332 3333 3334 3335 3336 3337 3338 3339 3340 3341 3342 3343
+ 3344 3345 3346 3347 3348 3349 3350 3351 3352 3353 3354 3355 3356 3357 3358 3359 3360 3361 3362 3363
+ 3364 3365 3366 3367 3368 3369 3370 3371 3372 3373 3374 3375 3376 3377 3378 3379 3380 3381 3382 3383
+ 3384 3385 3386 3387 3388 3389 3390 3391 3392 3393 3394 3395 3396 3397 3398 3399 3400 3401 3402 3403
+ 3404 3405 3406 3407 3408 3409 3410 3411 3412 3413 3414 3415 3416 3417 3418 3419 3420 3421 3422 3423
+ 3424 3425 3426 3427 3428 3429 3430 3431 3432 3433 3434
+ ICV_117 $T=79200 0 0 0 $X=78200 $Y=-1000
X3591 Q_5 VDD D_5 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 565 566 567 568 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 3435 3436 3437
+ 3438 3439 3440 3441 3442 3443 3444 3445 3446 3447 3448 3449 3450 3451 3452 3453 3454 3455 3456 3457
+ 3458 3459 3460 3461 3462 3463 3464 3465 3466 3467 3468 3469 3470 3471 3472 3473 3474 3475 3476 3477
+ 3478 3479 3480 3481 3482 3483 3484 3485 3486 3487 3488 3489 3490 3491 3492 3493 3494 3495 3496 3497
+ 3498 3499 3500 3501 3502 3503 3504 3505 3506 3507 3508 3509 3510 3511 3512 3513 3514 3515 3516 3517
+ 3518 3519 3520 3521 3522 3523 3524 3525 3526 3527 3528 3529 3530 3531 3532 3533 3534 3535 3536 3537
+ 3538 3539 3540 3541 3542 3543 3544 3545 3546 3547 3548 3549 3550 3551 3552 3553 3554 3555 3556 3557
+ 3558 3559 3560 3561 3562 3563 3564 3565 3566 3567 3568 3569 3570 3571 3572 3573 3574 3575 3576 3577
+ 3578 3579 3580 3581 3582 3583 3584 3585 3586 3587 3588 3589 3590 3591 3592 3593 3594 3595 3596 3597
+ 3598 3599 3600 3601 3602 3603 3604 3605 3606 3607 3608 3609 3610 3611 3612 3613 3614 3615 3616 3617
+ 3618 3619 3620 3621 3622 3623 3624 3625 3626 3627 3628 3629 3630 3631 3632 3633 3634 3635 3636 3637
+ 3638 3639 3640 3641 3642 3643 3644 3645 3646 3647 3648 3649 3650 3651 3652 3653 3654 3655 3656 3657
+ 3658 3659 3660 3661 3662 3663 3664 3665 3666 3667 3668 3669 3670 3671 3672 3673 3674 3675 3676 3677
+ 3678 3679 3680 3681 3682 3683 3684 3685 3686 3687 3688 3689 3690 3691 3692 3693 3694 3695 3696 3697
+ 3698 3699 3700 3701 3702 3703 3704 3705 3706 3707 3708 3709 3710 3711 3712 3713 3714 3715 3716 3717
+ 3718 3719 3720 3721 3722 3723 3724 3725 3726 3727 3728 3729 3730 3731 3732 3733 3734 3735 3736 3737
+ 3738 3739 3740 3741 3742 3743 3744 3745 3746 3747 3748 3749 3750 3751 3752 3753 3754 3755 3756 3757
+ 3758 3759 3760 3761 3762 3763 3764 3765 3766 3767 3768 3769 3770 3771 3772 3773 3774 3775 3776 3777
+ 3778 3779 3780 3781 3782 3783 3784 3785 3786 3787 3788 3789 3790 3791 3792 3793 3794 3795 3796 3797
+ 3798 3799 3800 3801 3802 3803 3804 3805 3806 3807 3808 3809 3810 3811 3812 3813 3814 3815 3816 3817
+ 3818 3819 3820 3821 3822 3823 3824 3825 3826 3827 3828 3829 3830 3831 3832 3833 3834 3835 3836 3837
+ 3838 3839 3840 3841 3842 3843 3844 3845 3846 3847 3848 3849 3850 3851 3852 3853 3854 3855 3856 3857
+ 3858 3859 3860 3861 3862 3863 3864 3865 3866 3867 3868 3869 3870 3871 3872 3873 3874 3875 3876 3877
+ 3878 3879 3880 3881 3882 3883 3884 3885 3886 3887 3888 3889 3890 3891 3892 3893 3894 3895 3896 3897
+ 3898 3899 3900 3901 3902 3903 3904 3905 3906 3907 3908 3909 3910 3911 3912 3913 3914 3915 3916 3917
+ 3918 3919 3920 3921 3922 3923 3924 3925 3926 3927 3928 3929 3930 3931 3932 3933 3934 3935 3936 3937
+ 3938 3939 3940 3941 3942 3943 3944 3945 3946 3947 3948
+ ICV_112 $T=117600 0 1 180 $X=97400 $Y=-1000
X3592 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_140 $T=0 0 0 90 $X=116600 $Y=62320
X3593 Q_6 VDD D_6 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ 569 570 571 572 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 3949 3950 3951
+ 3952 3953 3954 3955 3956 3957 3958 3959 3960 3961 3962 3963 3964 3965 3966 3967 3968 3969 3970 3971
+ 3972 3973 3974 3975 3976 3977 3978 3979 3980 3981 3982 3983 3984 3985 3986 3987 3988 3989 3990 3991
+ 3992 3993 3994 3995 3996 3997 3998 3999 4000 4001 4002 4003 4004 4005 4006 4007 4008 4009 4010 4011
+ 4012 4013 4014 4015 4016 4017 4018 4019 4020 4021 4022 4023 4024 4025 4026 4027 4028 4029 4030 4031
+ 4032 4033 4034 4035 4036 4037 4038 4039 4040 4041 4042 4043 4044 4045 4046 4047 4048 4049 4050 4051
+ 4052 4053 4054 4055 4056 4057 4058 4059 4060 4061 4062 4063 4064 4065 4066 4067 4068 4069 4070 4071
+ 4072 4073 4074 4075 4076 4077 4078 4079 4080 4081 4082 4083 4084 4085 4086 4087 4088 4089 4090 4091
+ 4092 4093 4094 4095 4096 4097 4098 4099 4100 4101 4102 4103 4104 4105 4106 4107 4108 4109 4110 4111
+ 4112 4113 4114 4115 4116 4117 4118 4119 4120 4121 4122 4123 4124 4125 4126 4127 4128 4129 4130 4131
+ 4132 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149 4150 4151
+ 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4165 4166 4167 4168 4169 4170 4171
+ 4172 4173 4174 4175 4176 4177 4178 4179 4180 4181 4182 4183 4184 4185 4186 4187 4188 4189 4190 4191
+ 4192 4193 4194 4195 4196 4197 4198 4199 4200 4201 4202 4203 4204 4205 4206 4207 4208 4209 4210 4211
+ 4212 4213 4214 4215 4216 4217 4218 4219 4220 4221 4222 4223 4224 4225 4226 4227 4228 4229 4230 4231
+ 4232 4233 4234 4235 4236 4237 4238 4239 4240 4241 4242 4243 4244 4245 4246 4247 4248 4249 4250 4251
+ 4252 4253 4254 4255 4256 4257 4258 4259 4260 4261 4262 4263 4264 4265 4266 4267 4268 4269 4270 4271
+ 4272 4273 4274 4275 4276 4277 4278 4279 4280 4281 4282 4283 4284 4285 4286 4287 4288 4289 4290 4291
+ 4292 4293 4294 4295 4296 4297 4298 4299 4300 4301 4302 4303 4304 4305 4306 4307 4308 4309 4310 4311
+ 4312 4313 4314 4315 4316 4317 4318 4319 4320 4321 4322 4323 4324 4325 4326 4327 4328 4329 4330 4331
+ 4332 4333 4334 4335 4336 4337 4338 4339 4340 4341 4342 4343 4344 4345 4346 4347 4348 4349 4350 4351
+ 4352 4353 4354 4355 4356 4357 4358 4359 4360 4361 4362 4363 4364 4365 4366 4367 4368 4369 4370 4371
+ 4372 4373 4374 4375 4376 4377 4378 4379 4380 4381 4382 4383 4384 4385 4386 4387 4388 4389 4390 4391
+ 4392 4393 4394 4395 4396 4397 4398 4399 4400 4401 4402 4403 4404 4405 4406 4407 4408 4409 4410 4411
+ 4412 4413 4414 4415 4416 4417 4418 4419 4420 4421 4422 4423 4424 4425 4426 4427 4428 4429 4430 4431
+ 4432 4433 4434 4435 4436 4437 4438 4439 4440 4441 4442 4443 4444 4445 4446 4447 4448 4449 4450 4451
+ 4452 4453 4454 4455 4456 4457 4458 4459 4460 4461 4462
+ ICV_107 $T=118800 0 0 0 $X=117800 $Y=-1000
X3594 VSS VDD D_7 Q_7 STUBDW_0 STUBDW__0 STUBDR_0 STUBDR__0 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_0 WE
+ OE_ 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595
+ 596 597 598 599 600 601 602 603 604 605 606 607 608
+ ICV_139 $T=0 0 0 90 $X=137000 $Y=-1000
X3595 VSS VDD WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17
+ WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37
+ WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57
+ WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77
+ WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97
+ WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117
+ WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137
+ WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157
+ WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177
+ WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197
+ WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217
+ WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237
+ WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255 578 579
+ 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599
+ 600 601 602 603 604 605 606 607 866 4463 867 4464 868 4465 869 4466 870 4467 871 4468
+ 872 4469 873 4470 874 4471 875 4472 876 4473 877 4474 878 4475 879 4476 880 4477 881 4478
+ 882 4479 883 4480 884 4481 885 4482 886 4483 887 4484 888 4485 889 4486 890 4487 891 4488
+ 892 4489 893 4490 894 4491 895 4492 896 4493 897 4494 898 4495 899 4496 900 4497 901 4498
+ 902 4499 903 4500 904 4501 905 4502 906 4503 907 4504 908 4505 909 4506 910 4507 911 4508
+ 912 4509 913 4510 914 4511 915 4512 916 4513 917 4514 918 4515 919 4516 920 4517 921 4518
+ 922 4519 923 4520 924 4521 925 4522 926 4523 927 4524 928 4525 929 4526 930 4527 931 4528
+ 932 4529 933 4530 934 4531 935 4532 936 4533 937 4534 938 4535 939 4536 940 4537 941 4538
+ 942 4539 943 4540 944 4541 945 4542 946 4543 947 4544 948 4545 949 4546 950 4547 951 4548
+ 952 4549 953 4550 954 4551 955 4552 956 4553 957 4554 958 4555 959 4556 960 4557 961 4558
+ 962 4559 963 4560 964 4561 965 4562 966 4563 967 4564 968 4565 969 4566 970 4567 971 4568
+ 972 4569 973 4570 974 4571 975 4572 976 4573 977 4574 978 4575 979 4576 980 4577 981 4578
+ 982 4579 983 4580 984 4581 985 4582 986 4583 987 4584 988 4585 989 4586 990 4587 991 4588
+ 992 4589 993 4590 994 4591 995 4592 996 4593 997 4594 998 4595 999 4596 1000 4597 1001 4598
+ 1002 4599 1003 4600 1004 4601 1005 4602 1006 4603 1007 4604 1008 4605 1009 4606 1010 4607 1011 4608
+ 1012 4609 1013 4610 1014 4611 1015 4612 1016 4613 1017 4614 1018 4615 1019 4616 1020 4617 1021 4618
+ 1022 4619 1023 4620 1024 4621 1025 4622 1026 4623 1027 4624 1028 4625 1029 4626 1030 4627 1031 4628
+ 1032 4629 1033 4630 1034 4631 1035 4632 1036 4633 1037 4634 1038 4635 1039 4636 1040 4637 1041 4638
+ 1042 4639 1043 4640 1044 4641 1045 4642 1046 4643 1047 4644 1048 4645 1049 4646 1050 4647 1051 4648
+ 1052 4649 1053 4650 1054 4651 1055 4652 1056 4653 1057 4654 1058 4655 1059 4656 1060 4657 1061 4658
+ 1062 4659 1063 4660 1064 4661 1065 4662 1066 4663 1067 4664 1068 4665 1069 4666 1070 4667 1071 4668
+ 1072 4669 1073 4670 1074 4671 1075 4672 1076 4673 1077 4674 1078 4675 1079 4676 1080 4677 1081 4678
+ 1082 4679 1083 4680 1084 4681 1085 4682 1086 4683 1087 4684 1088 4685 1089 4686 1090 4687 1091 4688
+ 1092 4689 1093 4690 1094 4691 1095 4692 1096 4693 1097 4694 1098 4695 1099 4696 1100 4697 1101 4698
+ 1102 4699 1103 4700 1104 4701 1105 4702 1106 4703 1107 4704 1108 4705 1109 4706 1110 4707 1111 4708
+ 1112 4709 1113 4710 1114 4711 1115 4712 1116 4713 1117 4714 1118 4715 1119 4716 1120 4717 1121 4718
+ ICV_138 $T=0 0 0 90 $X=137000 $Y=61500
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT SIGN_MEMFC4T
** N=22 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD BL0 BL0_ BL1 BL1_ BL2 BL2_ BL3 BL3_
.ENDS
***************************************
.SUBCKT base_flmo_nvpv 2 4 7 8
** N=18 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 2 8 7 2 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=380 $Y=850 $D=103
M1 8 7 2 2 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=850 $D=103
M2 4 8 7 4 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=370 $Y=260 $D=192
M3 8 7 4 4 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=260 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMFC1TL
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS
.ENDS
***************************************
.SUBCKT ntapCont_0_16_0_16_8_1_0_4_0_4_center_center
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCWD
** N=4 EP=0 IP=2 FDC=0
*.CALIBRE ISOLATED NETS: VDD WL0 VSS WL1
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT ai 1 2 3 4 5 6
** N=89 EP=6 IP=0 FDC=14
M0 4 9 1 1 lpnfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=6980 $D=103
M1 1 9 4 1 lpnfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=6980 $D=103
M2 9 2 1 1 lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=6980 $D=103
M3 1 2 9 1 lpnfet w=9.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=6980 $D=103
M4 5 2 1 1 lpnfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2620 $Y=6980 $D=103
M5 1 2 5 1 lpnfet w=1.22e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=6980 $D=103
M6 4 9 3 3 lppfet w=2.42e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=3370 $D=192
M7 3 9 4 3 lppfet w=2.42e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=3370 $D=192
M8 9 2 3 3 lppfet w=1.94e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=3850 $D=192
M9 3 2 9 3 lppfet w=1.94e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=3850 $D=192
M10 5 2 3 3 lppfet w=2.42e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2620 $Y=3370 $D=192
M11 3 2 5 3 lppfet w=2.42e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=3370 $D=192
D12 1 2 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1540 $Y=140 $D=558
D13 1 6 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1550 $Y=800 $D=558
.ENDS
***************************************
.SUBCKT ap 1 2 3 4 5 16 17 18 19 20
** N=613 EP=10 IP=0 FDC=76
M0 3 24 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=0 $D=103
M1 4 25 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=49910 $D=103
M2 1 17 21 1 lpnfet w=1.76e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=520 $Y=23290 $D=103
M3 31 21 1 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=760 $Y=12370 $D=103
M4 32 21 1 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=760 $Y=35540 $D=103
M5 1 24 3 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=0 $D=103
M6 1 25 4 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=49910 $D=103
M7 22 18 1 1 lpnfet w=1.76e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1000 $Y=23290 $D=103
M8 24 29 27 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1020 $Y=9720 $D=103
M9 25 30 28 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1020 $Y=40530 $D=103
M10 33 26 31 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1080 $Y=12370 $D=103
M11 34 26 32 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1080 $Y=35540 $D=103
M12 3 24 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=0 $D=103
M13 27 23 33 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=12370 $D=103
M14 28 22 34 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=35540 $D=103
M15 4 25 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=49910 $D=103
M16 27 29 24 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1500 $Y=9720 $D=103
M17 28 30 25 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1500 $Y=40530 $D=103
M18 1 24 3 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=0 $D=103
M19 35 23 27 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=12370 $D=103
M20 36 22 28 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=35540 $D=103
M21 1 25 4 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=49910 $D=103
M22 24 29 27 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1980 $Y=9720 $D=103
M23 25 30 28 1 lpnfet w=1.28e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1980 $Y=40530 $D=103
M24 37 26 35 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2200 $Y=12370 $D=103
M25 38 26 36 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2200 $Y=35540 $D=103
M26 1 19 23 1 lpnfet w=1.76e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2280 $Y=23290 $D=103
M27 3 24 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=0 $D=103
M28 4 25 1 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=49910 $D=103
M29 1 3 24 1 lpnfet w=1.6e-07 l=3.6e-07 m=1 par=1 nf=1 ngcon=1 $X=2500 $Y=10840 $D=103
M30 1 4 25 1 lpnfet w=1.6e-07 l=3.6e-07 m=1 par=1 nf=1 ngcon=1 $X=2500 $Y=40530 $D=103
M31 1 21 37 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=12370 $D=103
M32 1 21 38 1 lpnfet w=3.82e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=35540 $D=103
M33 26 20 1 1 lpnfet w=1.76e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2760 $Y=23290 $D=103
M34 1 24 3 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=0 $D=103
M35 1 25 4 1 lpnfet w=1.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=49910 $D=103
M36 1 5 29 1 lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=9950 $D=103
M37 1 16 30 1 lpnfet w=5.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=41000 $D=103
M38 3 24 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=2770 $D=192
M39 27 21 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=17570 $D=192
M40 28 21 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=30960 $D=192
M41 4 25 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=440 $Y=45840 $D=192
M42 2 17 21 2 lppfet w=3.56e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=520 $Y=26330 $D=192
M43 2 24 3 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=2770 $D=192
M44 2 21 27 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=17570 $D=192
M45 2 21 28 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=30960 $D=192
M46 2 25 4 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=920 $Y=45840 $D=192
M47 22 18 2 2 lppfet w=3.56e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1000 $Y=26330 $D=192
M48 24 5 27 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1020 $Y=6390 $D=192
M49 25 16 28 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1020 $Y=42960 $D=192
M50 3 24 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=2770 $D=192
M51 27 23 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=17570 $D=192
M52 28 22 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=30960 $D=192
M53 4 25 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1400 $Y=45840 $D=192
M54 27 5 24 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1500 $Y=6390 $D=192
M55 28 16 25 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1500 $Y=42960 $D=192
M56 2 24 3 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=2770 $D=192
M57 2 23 27 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=17570 $D=192
M58 2 22 28 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=30960 $D=192
M59 2 25 4 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1880 $Y=45840 $D=192
M60 24 5 27 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1980 $Y=6390 $D=192
M61 25 16 28 2 lppfet w=2.14e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1980 $Y=42960 $D=192
M62 2 19 23 2 lppfet w=3.56e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2280 $Y=26330 $D=192
M63 3 24 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=2770 $D=192
M64 27 26 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=17570 $D=192
M65 28 26 2 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=30960 $D=192
M66 4 25 2 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2360 $Y=45840 $D=192
M67 2 3 24 2 lppfet w=1.6e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=7040 $D=192
M68 2 4 25 2 lppfet w=1.6e-07 l=1.8e-07 m=1 par=1 nf=1 ngcon=1 $X=2520 $Y=44290 $D=192
M69 26 20 2 2 lppfet w=3.56e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2760 $Y=26330 $D=192
M70 2 24 3 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=2770 $D=192
M71 2 26 27 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=17570 $D=192
M72 2 26 28 2 lppfet w=3.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=30960 $D=192
M73 2 25 4 2 lppfet w=2.88e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2840 $Y=45840 $D=192
M74 2 5 29 2 lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=7630 $D=192
M75 2 16 30 2 lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=42960 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDG0T
** N=43 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WL0 WL1 G0 XP1F XP0F
.ENDS
***************************************
.SUBCKT ptapCont_0_16_0_16_6_2_0_4_0_4_center_center
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDGF VSS
** N=18 EP=1 IP=1 FDC=1
*.CALIBRE ISOLATED NETS: VDD WL0 WL1 XP1 XP0
M0 VSS VSS VSS VSS nfet L=9.2e-07 W=2.36e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=300 $Y=1880 $D=97
.ENDS
***************************************
.SUBCKT ndiffCont_0_16_0_16_5_1_0_4_0_4_center_center
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ptapCont_0_16_0_16_5_2_0_4_0_4_center_center
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDG1M
** N=9 EP=0 IP=1 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WL0 WL1 XP1F XP0F G1
.ENDS
***************************************
.SUBCKT ptapCont_0_16_0_16_14_2_0_4_0_4_center_center
** N=29 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SIGN_MEMWD VSS VDD G0 WL0 WL1 GTP G1 G2_W0 G2_W1
** N=488 EP=9 IP=3 FDC=47
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0
M0 26 G2_W0 22 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=810 $D=103
M1 27 G1 26 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=1130 $D=103
M2 VSS G0 27 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=1450 $D=103
M3 28 G0 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=1930 $D=103
M4 29 G1 28 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=2250 $D=103
M5 23 G2_W1 29 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=2570 $D=103
M6 18 22 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=880 $D=103
M7 GTP 25 18 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=1400 $D=103
M8 19 24 GTP VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=1880 $D=103
M9 VSS 23 19 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=2400 $D=103
M10 VSS 23 24 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14790 $Y=2950 $D=103
M11 25 22 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14810 $Y=360 $D=103
M12 20 18 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=180 $D=103
M13 VSS 18 20 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=660 $D=103
M14 20 18 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=1140 $D=103
M15 VSS 19 21 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=2140 $D=103
M16 21 19 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=2620 $D=103
M17 VSS 19 21 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=3100 $D=103
M18 WL0 20 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=180 $D=103
M19 VSS 20 WL0 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=660 $D=103
M20 WL0 20 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=1140 $D=103
M21 VSS 21 WL1 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=2140 $D=103
M22 WL1 21 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=2620 $D=103
M23 VSS 21 WL1 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=3100 $D=103
M24 VSS VSS VSS VSS nfet L=9.2e-07 W=5.44e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=1880 $D=97
M25 22 G2_W0 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=180 $D=192
M26 VDD G1 22 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=660 $D=192
M27 22 G0 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=1140 $D=192
M28 VDD G0 23 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=2140 $D=192
M29 23 G1 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=2620 $D=192
M30 VDD G2_W1 23 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=3100 $D=192
M31 GTP 22 18 VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11960 $Y=1400 $D=192
M32 19 23 GTP VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11960 $Y=1880 $D=192
M33 VDD 23 24 VDD lppfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=12320 $Y=3100 $D=192
M34 25 22 VDD VDD lppfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=12400 $Y=180 $D=192
M35 20 18 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=180 $D=192
M36 VDD 18 20 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=660 $D=192
M37 20 18 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=1140 $D=192
M38 VDD 19 21 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=2140 $D=192
M39 21 19 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=2620 $D=192
M40 VDD 19 21 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=3100 $D=192
M41 WL0 20 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=180 $D=192
M42 VDD 20 WL0 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=660 $D=192
M43 WL0 20 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=1140 $D=192
M44 VDD 21 WL1 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=2140 $D=192
M45 WL1 21 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=2620 $D=192
M46 VDD 21 WL1 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=3100 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMWD0 VSS VDD XP2_1 XP2_0 G0 WL0 WL1 GTP G1
** N=15 EP=9 IP=17 FDC=47
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2
X0 VSS VDD G0 WL0 WL1 GTP G1 XP2_0 XP2_1 SIGN_MEMWD $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMROW_8 VSS VDD WL0 WL1 G0 XP2_1 XP2_0 GTP G1
** N=32 EP=9 IP=44 FDC=50
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP1F_0 XP0F_0 XP1F_3 XP0F_3 G1B XP1_0 XP0_0 XP1_1 XP0_1 XP1F_1 XP0F_1 XP1F_2 XP0F_2
M0 VSS VSS VSS VSS nfet L=9.2e-07 W=2.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=7660 $Y=620 $D=97
X1 VSS SIGN_MEMFLWDGF $T=0 0 0 0 $X=-1000 $Y=-1000
X2 VSS SIGN_MEMFLWDGF $T=3400 0 0 0 $X=2400 $Y=-1000
X8 VSS VDD XP2_1 XP2_0 G0 WL0 WL1 GTP G1 SIGN_MEMWD0 $T=20400 0 0 0 $X=19400 $Y=-1000
.ENDS
***************************************
.SUBCKT VPC_M1_CDNS_6479038850981
** N=25 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDMMM
** N=8 EP=0 IP=2 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WL0 WL1 G0 XP1F XP0F G1
.ENDS
***************************************
.SUBCKT SIGN_MEMROW_FILLER3 VSS VDD XP2_7 XP2_6 WL0 WL1 G0 GTP G1
** N=27 EP=9 IP=55 FDC=52
*.CALIBRE ISOLATED NETS: XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 XP1_0 XP0_0 XP1_1 XP0_1 XP1_2 XP0_2 XP1_3 XP0_3 XP1_4 XP0_4 XP1F XP0F
X0 VSS SIGN_MEMFLWDGF $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS SIGN_MEMFLWDGF $T=3400 0 0 0 $X=2400 $Y=-1000
X2 VSS SIGN_MEMFLWDGF $T=6800 0 0 0 $X=5800 $Y=-1000
X3 VSS SIGN_MEMFLWDGF $T=10200 0 0 0 $X=9200 $Y=-1000
X4 VSS SIGN_MEMFLWDGF $T=13600 0 0 0 $X=12600 $Y=-1000
X5 VSS VDD G0 WL0 WL1 GTP G1 XP2_7 XP2_6 SIGN_MEMWD $T=20400 0 0 0 $X=19400 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMROW_FILLER2 VSS VDD XP2_5 XP2_4 WL0 WL1 G0 GTP G1
** N=27 EP=9 IP=55 FDC=52
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_3 XP2_2 XP2_1 XP2_0 XP1_0 XP0_0 XP1_1 XP0_1 XP1_2 XP0_2 XP1_3 XP0_3 XP1_4 XP0_4 XP1F XP0F
X0 VSS SIGN_MEMFLWDGF $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS SIGN_MEMFLWDGF $T=3400 0 0 0 $X=2400 $Y=-1000
X2 VSS SIGN_MEMFLWDGF $T=6800 0 0 0 $X=5800 $Y=-1000
X3 VSS SIGN_MEMFLWDGF $T=10200 0 0 0 $X=9200 $Y=-1000
X4 VSS SIGN_MEMFLWDGF $T=13600 0 0 0 $X=12600 $Y=-1000
X5 VSS VDD G0 WL0 WL1 GTP G1 XP2_4 XP2_5 SIGN_MEMWD $T=20400 0 0 0 $X=19400 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMROW_FILLER1 VSS VDD XP2_3 XP2_2 WL0 WL1 G0 GTP G1
** N=27 EP=9 IP=55 FDC=52
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_1 XP2_0 XP1_0 XP0_0 XP1_1 XP0_1 XP1_2 XP0_2 XP1_3 XP0_3 XP1_4 XP0_4 XP1F XP0F
X0 VSS SIGN_MEMFLWDGF $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS SIGN_MEMFLWDGF $T=3400 0 0 0 $X=2400 $Y=-1000
X2 VSS SIGN_MEMFLWDGF $T=6800 0 0 0 $X=5800 $Y=-1000
X3 VSS SIGN_MEMFLWDGF $T=10200 0 0 0 $X=9200 $Y=-1000
X4 VSS SIGN_MEMFLWDGF $T=13600 0 0 0 $X=12600 $Y=-1000
X5 VSS VDD G0 WL0 WL1 GTP G1 XP2_3 XP2_2 SIGN_MEMWD $T=20400 0 0 0 $X=19400 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_99 1 2 3 4 7 8 9 10 13 14 15 26 29
** N=29 EP=13 IP=54 FDC=104
X0 1 2 7 8 3 4 26 13 29 SIGN_MEMROW_FILLER2 $T=0 0 1 0 $X=-1000 $Y=-4400
X1 1 2 9 10 14 15 26 13 29 SIGN_MEMROW_FILLER1 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_100 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 30
+ 33 34
** N=34 EP=22 IP=84 FDC=206
X0 1 2 3 4 30 11 12 13 34 SIGN_MEMROW_8 $T=0 -6800 1 0 $X=-1000 $Y=-11200
X1 1 2 5 6 14 15 30 13 33 SIGN_MEMROW_FILLER3 $T=0 -6800 0 0 $X=-1000 $Y=-7800
X2 1 2 17 16 7 8 9 10 13 18 19 30 33 ICV_99 $T=0 0 0 0 $X=-1000 $Y=-4400
.ENDS
***************************************
.SUBCKT ICV_101 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 38 41 42 43
** N=43 EP=31 IP=68 FDC=412
X0 1 2 4 3 11 12 13 14 15 16 17 18 19 5 6 7 8 9 10 38
+ 42 41
+ ICV_100 $T=0 -13600 0 0 $X=-1000 $Y=-24800
X1 1 2 21 20 11 12 13 14 15 16 17 18 19 22 23 24 25 26 27 38
+ 43 42
+ ICV_100 $T=0 0 0 0 $X=-1000 $Y=-11200
.ENDS
***************************************
.SUBCKT ICV_102 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 51 52 53 54 55 56
** N=56 EP=49 IP=86 FDC=824
X0 1 2 3 4 5 6 7 8 9 10 19 20 21 22 23 24 25 26 27 11
+ 12 13 14 15 16 17 18 54 51 52 53
+ ICV_101 $T=0 -27200 0 0 $X=-1000 $Y=-52000
X1 1 2 28 29 30 31 32 33 34 35 19 20 21 22 23 24 25 26 27 36
+ 37 38 39 40 41 42 43 54 53 55 56
+ ICV_101 $T=0 0 0 0 $X=-1000 $Y=-24800
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDG0B
** N=43 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WL0 G0 WL1 XP1F XP0F
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDG1T VSS
** N=12 EP=1 IP=2 FDC=1
*.CALIBRE ISOLATED NETS: VDD WL0 G0 WL1 XP1F XP0F G1
M0 VSS VSS VSS VSS nfet L=9.2e-07 W=2.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=860 $Y=620 $D=97
.ENDS
***************************************
.SUBCKT SIGN_MEMFLWDG1B
** N=10 EP=0 IP=1 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD WL0 G0 WL1 XP1F XP0F G1
.ENDS
***************************************
.SUBCKT SIGN_MEMROW_64 VSS VDD WL0 G0 WL1 XP2_1 XP2_0 GTP G1
** N=29 EP=9 IP=54 FDC=48
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 G0B XP1F_5 XP0F_5 G1B XP1F_0 XP0F_0 XP1F_1 XP0F_1 XP1F_2 XP0F_2 XP1F_3 XP0F_3 XP1F_4 XP0F_4
X2 VSS VDD XP2_1 XP2_0 G0 WL0 WL1 GTP G1 SIGN_MEMWD0 $T=20400 0 0 0 $X=19400 $Y=-1000
X4 VSS SIGN_MEMFLWDG1T $T=6800 0 0 0 $X=5800 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMFCMWDX VSS XP1 XP0
** N=14 EP=3 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: VDD MWL
D0 VSS XP1 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1110 $Y=520 $D=558
D1 VSS XP0 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=1890 $Y=520 $D=558
.ENDS
***************************************
.SUBCKT SIGN_MEMHWDB0 VSS VDD G0 WL0 WL1 XP2_1 XP2_0 GTP G1
** N=488 EP=9 IP=3 FDC=47
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2
M0 24 XP2_0 20 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=3740 $D=103
M1 25 G1 24 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=4060 $D=103
M2 VSS G0 25 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=4380 $D=103
M3 26 G0 VSS VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=4860 $D=103
M4 27 G1 26 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=5180 $D=103
M5 21 XP2_1 27 VSS lpnfet w=8.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7570 $Y=5500 $D=103
M6 16 20 VSS VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=3810 $D=103
M7 GTP 23 16 VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=4330 $D=103
M8 17 22 GTP VSS lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=4810 $D=103
M9 VSS 21 17 VSS lpnfet w=2.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14110 $Y=5330 $D=103
M10 VSS 21 22 VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14790 $Y=5880 $D=103
M11 23 20 VSS VSS lpnfet w=2.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=14810 $Y=3290 $D=103
M12 18 16 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=3110 $D=103
M13 VSS 16 18 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=3590 $D=103
M14 18 16 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=4070 $D=103
M15 VSS 17 19 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=5070 $D=103
M16 19 17 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=5550 $D=103
M17 VSS 17 19 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=6030 $D=103
M18 WL0 18 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=3110 $D=103
M19 VSS 18 WL0 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=3590 $D=103
M20 WL0 18 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=4070 $D=103
M21 VSS 19 WL1 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=5070 $D=103
M22 WL1 19 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=5550 $D=103
M23 VSS 19 WL1 VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=6030 $D=103
M24 VSS VSS VSS VSS nfet L=9.2e-07 W=5.44e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=420 $Y=4810 $D=97
M25 20 XP2_0 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=3110 $D=192
M26 VDD G1 20 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=3590 $D=192
M27 20 G0 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=4070 $D=192
M28 VDD G0 21 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=5070 $D=192
M29 21 G1 VDD VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=5550 $D=192
M30 VDD XP2_1 21 VDD lppfet w=6.8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10510 $Y=6030 $D=192
M31 GTP 20 16 VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11960 $Y=4330 $D=192
M32 17 21 GTP VDD lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11960 $Y=4810 $D=192
M33 VDD 21 22 VDD lppfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=12320 $Y=6030 $D=192
M34 23 20 VDD VDD lppfet w=4.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=12400 $Y=3110 $D=192
M35 18 16 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=3110 $D=192
M36 VDD 16 18 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=3590 $D=192
M37 18 16 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=4070 $D=192
M38 VDD 17 19 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=5070 $D=192
M39 19 17 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=5550 $D=192
M40 VDD 17 19 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=6030 $D=192
M41 WL0 18 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=3110 $D=192
M42 VDD 18 WL0 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=3590 $D=192
M43 WL0 18 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=4070 $D=192
M44 VDD 19 WL1 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=5070 $D=192
M45 WL1 19 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=5550 $D=192
M46 VDD 19 WL1 VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=6030 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMMWDX VSS VDD MWL GTP MBL MWLD MBL_
** N=461 EP=7 IP=0 FDC=49
*.CALIBRE ISOLATED NETS: XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0
M0 GTP VDD 17 VSS lpnfet w=7e-07 l=2.4e-07 m=1 par=1 nf=1 ngcon=1 $X=14670 $Y=980 $D=103
M1 VSS 17 18 VSS lpnfet w=2.8e-07 l=1.6e-07 m=1 par=1 nf=1 ngcon=1 $X=17390 $Y=1180 $D=103
M2 19 18 VSS VSS lpnfet w=2.8e-07 l=1.6e-07 m=1 par=1 nf=1 ngcon=1 $X=17390 $Y=1860 $D=103
M3 16 19 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=180 $D=103
M4 VSS 19 16 VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=660 $D=103
M5 16 19 VSS VSS lpnfet w=1.68e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=18470 $Y=1140 $D=103
M6 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=28300 $Y=2860 $D=103
M7 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=28300 $Y=3860 $D=103
M8 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=29060 $Y=2860 $D=103
M9 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=29060 $Y=3860 $D=103
M10 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=30040 $Y=2860 $D=103
M11 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=30040 $Y=3860 $D=103
M12 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=30800 $Y=2860 $D=103
M13 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=30800 $Y=3860 $D=103
M14 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=31780 $Y=2860 $D=103
M15 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=31780 $Y=3860 $D=103
M16 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=32540 $Y=2860 $D=103
M17 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=32540 $Y=3860 $D=103
M18 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=33520 $Y=2860 $D=103
M19 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=33520 $Y=3860 $D=103
M20 MBL VSS VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=34280 $Y=2860 $D=103
M21 VSS VSS MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=34280 $Y=3860 $D=103
M22 MBL MWLD VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=35260 $Y=2860 $D=103
M23 VSS MWLD MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=35260 $Y=3860 $D=103
M24 MWL 16 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=180 $D=103
M25 VSS 16 MWL VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=660 $D=103
M26 MWL 16 VSS VSS lpnfet w=4.18e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=36010 $Y=1140 $D=103
M27 MBL MWLD VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=36020 $Y=2860 $D=103
M28 VSS MWLD MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=36020 $Y=3860 $D=103
M29 MBL MWLD VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=37000 $Y=2860 $D=103
M30 VSS MWLD MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=37000 $Y=3860 $D=103
M31 MBL MWLD VSS VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=37760 $Y=2860 $D=103
M32 VSS MWLD MBL VSS lpnfet w=2.1e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=37760 $Y=3860 $D=103
M33 MBL MWLD VSS VSS lpnfet w=1.6e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=38760 $Y=2860 $D=103
M34 VSS MWLD MBL VSS lpnfet w=1.6e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=38760 $Y=3860 $D=103
M35 MBL MWLD VSS VSS lpnfet w=1.6e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=39520 $Y=2860 $D=103
M36 VSS MWLD MBL VSS lpnfet w=1.6e-07 l=5.6e-07 m=1 par=1 nf=1 ngcon=1 $X=39520 $Y=3860 $D=103
M37 MBL_ GTP VDD VDD lppfet w=6.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5730 $Y=1780 $D=192
M38 MBL GTP MBL_ VDD lppfet w=6.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5730 $Y=2260 $D=192
M39 VDD GTP MBL VDD lppfet w=6.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5730 $Y=2740 $D=192
M40 GTP VSS 17 VDD lppfet w=7e-07 l=2.4e-07 m=1 par=1 nf=1 ngcon=1 $X=12670 $Y=980 $D=192
M41 VDD 17 18 VDD lppfet w=4.6e-07 l=1.6e-07 m=1 par=1 nf=1 ngcon=1 $X=16330 $Y=1180 $D=192
M42 19 18 VDD VDD lppfet w=4.6e-07 l=1.6e-07 m=1 par=1 nf=1 ngcon=1 $X=16330 $Y=1860 $D=192
M43 16 19 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=180 $D=192
M44 VDD 19 16 VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=660 $D=192
M45 16 19 VDD VDD lppfet w=3.52e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=22060 $Y=1140 $D=192
M46 MWL 16 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=180 $D=192
M47 VDD 16 MWL VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=660 $D=192
M48 MWL 16 VDD VDD lppfet w=7.58e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=26590 $Y=1180 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMWORD_ROWS VSS VDD XP1_0 XP0_0 XP1_1 XP0_1 WL0_0 WL1_0 MWL WL0_31 WL1_31 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP
+ WL0_63 WL1_63 WL0_95 WL1_95 WL0_127 WL1_127 WL1_30 WL0_30 WL0_29 WL1_29 WL1_62 WL0_62 WL0_61 WL1_61 WL1_94 WL0_94 WL0_93 WL1_93 WL1_126 WL0_126
+ WL0_125 WL1_125 WL1_28 WL0_28 WL0_27 WL1_27 WL1_26 WL0_26 WL0_25 WL1_25 WL1_60 WL0_60 WL0_59 WL1_59 WL1_58 WL0_58 WL0_57 WL1_57 WL1_92 WL0_92
+ WL0_91 WL1_91 WL1_90 WL0_90 WL0_89 WL1_89 WL1_124 WL0_124 WL0_123 WL1_123 WL1_122 WL0_122 WL0_121 WL1_121 WL1_24 WL0_24 WL0_23 WL1_23 WL1_22 WL0_22
+ WL0_21 WL1_21 WL1_20 WL0_20 WL0_19 WL1_19 WL1_18 WL0_18 WL0_17 WL1_17 WL1_56 WL0_56 WL0_55 WL1_55 WL1_54 WL0_54 WL0_53 WL1_53 WL1_52 WL0_52
+ WL0_51 WL1_51 WL1_50 WL0_50 WL0_49 WL1_49 WL1_88 WL0_88 WL0_87 WL1_87 WL1_86 WL0_86 WL0_85 WL1_85 WL1_84 WL0_84 WL0_83 WL1_83 WL1_82 WL0_82
+ WL0_81 WL1_81 WL1_120 WL0_120 WL0_119 WL1_119 WL1_118 WL0_118 WL0_117 WL1_117 WL1_116 WL0_116 WL0_115 WL1_115 WL1_114 WL0_114 WL0_113 WL1_113 WL1_16 WL0_16
+ WL0_15 WL1_15 WL1_14 WL0_14 WL0_13 WL1_13 WL1_12 WL0_12 WL0_11 WL1_11 WL1_10 WL0_10 WL0_9 WL1_9 WL1_8 WL0_8 WL0_7 WL1_7 WL1_6 WL0_6
+ WL0_5 WL1_5 WL1_4 WL0_4 WL0_3 WL1_3 WL1_2 WL0_2 WL0_1 WL1_1 WL1_48 WL0_48 WL0_47 WL1_47 WL1_46 WL0_46 WL0_45 WL1_45 WL1_44 WL0_44
+ WL0_43 WL1_43 WL1_42 WL0_42 WL0_41 WL1_41 WL1_40 WL0_40 WL0_39 WL1_39 WL1_38 WL0_38 WL0_37 WL1_37 WL1_36 WL0_36 WL0_35 WL1_35 WL1_34 WL0_34
+ WL0_33 WL1_33 WL1_80 WL0_80 WL0_79 WL1_79 WL1_78 WL0_78 WL0_77 WL1_77 WL1_76 WL0_76 WL0_75 WL1_75 WL1_74 WL0_74 WL0_73 WL1_73 WL1_72 WL0_72
+ WL0_71 WL1_71 WL1_70 WL0_70 WL0_69 WL1_69 WL1_68 WL0_68 WL0_67 WL1_67 WL1_66 WL0_66 WL0_65 WL1_65 WL1_112 WL0_112 WL0_111 WL1_111 WL1_110 WL0_110
+ WL0_109 WL1_109 WL1_108 WL0_108 WL0_107 WL1_107 WL1_106 WL0_106 WL0_105 WL1_105 WL1_104 WL0_104 WL0_103 WL1_103 WL1_102 WL0_102 WL0_101 WL1_101 WL1_100 WL0_100
+ WL0_99 WL1_99 WL1_98 WL0_98 WL0_97 WL1_97 WL0_32 WL1_32 WL0_64 WL1_64 WL0_96 WL1_96 MBL MWLD MBL_ XP1_2 XP0_2 XP1_3 XP0_3 XP1_4
+ XP0_4 XP1_5 XP0_5
** N=292 EP=283 IP=936 FDC=6645
D0 VSS XP1_5 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=18110 $Y=438650 $D=558
D1 VSS XP0_5 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=18890 $Y=438650 $D=558
X3 VSS VDD XP2_7 XP2_6 WL0_31 WL1_31 XP0_1 GTP XP1_2 SIGN_MEMROW_FILLER3 $T=0 111730 1 0 $X=-1000 $Y=107330
X4 VSS VDD XP2_7 XP2_6 WL0_63 WL1_63 XP1_1 GTP XP1_2 SIGN_MEMROW_FILLER3 $T=0 220530 1 0 $X=-1000 $Y=216130
X5 VSS VDD XP2_7 XP2_6 WL0_95 WL1_95 XP0_0 GTP XP1_2 SIGN_MEMROW_FILLER3 $T=0 329330 1 0 $X=-1000 $Y=324930
X6 VSS VDD XP2_7 XP2_6 WL0_127 WL1_127 XP1_0 GTP XP1_2 SIGN_MEMROW_FILLER3 $T=0 438130 1 0 $X=-1000 $Y=433730
X7 VSS VDD WL0_30 WL1_30 XP2_5 XP2_4 XP2_3 XP2_2 GTP WL0_29 WL1_29 XP0_1 XP1_2 ICV_99 $T=0 104930 1 0 $X=-1000 $Y=100530
X8 VSS VDD WL0_62 WL1_62 XP2_5 XP2_4 XP2_3 XP2_2 GTP WL0_61 WL1_61 XP1_1 XP1_2 ICV_99 $T=0 213730 1 0 $X=-1000 $Y=209330
X9 VSS VDD WL0_94 WL1_94 XP2_5 XP2_4 XP2_3 XP2_2 GTP WL0_93 WL1_93 XP0_0 XP1_2 ICV_99 $T=0 322530 1 0 $X=-1000 $Y=318130
X10 VSS VDD WL0_126 WL1_126 XP2_5 XP2_4 XP2_3 XP2_2 GTP WL0_125 WL1_125 XP1_0 XP1_2 ICV_99 $T=0 431330 1 0 $X=-1000 $Y=426930
X11 VSS VDD WL0_28 WL1_28 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL0_27 WL1_27 WL1_26 WL0_26 WL0_25 WL1_25 XP0_1
+ XP0_2 XP1_2
+ ICV_100 $T=0 91330 1 0 $X=-1000 $Y=86930
X12 VSS VDD WL0_60 WL1_60 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL0_59 WL1_59 WL1_58 WL0_58 WL0_57 WL1_57 XP1_1
+ XP0_2 XP1_2
+ ICV_100 $T=0 200130 1 0 $X=-1000 $Y=195730
X13 VSS VDD WL0_92 WL1_92 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL0_91 WL1_91 WL1_90 WL0_90 WL0_89 WL1_89 XP0_0
+ XP0_2 XP1_2
+ ICV_100 $T=0 308930 1 0 $X=-1000 $Y=304530
X14 VSS VDD WL0_124 WL1_124 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL0_123 WL1_123 WL1_122 WL0_122 WL0_121 WL1_121 XP1_0
+ XP0_2 XP1_2
+ ICV_100 $T=0 417730 1 0 $X=-1000 $Y=413330
X15 VSS VDD WL1_24 WL0_24 WL0_23 WL1_23 WL1_22 WL0_22 WL0_21 WL1_21 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_20
+ WL0_20 WL0_19 WL1_19 WL1_18 WL0_18 WL0_17 WL1_17 XP0_1 XP0_2 XP1_3 XP0_3
+ ICV_101 $T=0 64130 1 0 $X=-1000 $Y=59730
X16 VSS VDD WL1_56 WL0_56 WL0_55 WL1_55 WL1_54 WL0_54 WL0_53 WL1_53 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_52
+ WL0_52 WL0_51 WL1_51 WL1_50 WL0_50 WL0_49 WL1_49 XP1_1 XP0_2 XP1_3 XP0_3
+ ICV_101 $T=0 172930 1 0 $X=-1000 $Y=168530
X17 VSS VDD WL1_88 WL0_88 WL0_87 WL1_87 WL1_86 WL0_86 WL0_85 WL1_85 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_84
+ WL0_84 WL0_83 WL1_83 WL1_82 WL0_82 WL0_81 WL1_81 XP0_0 XP0_2 XP1_3 XP0_3
+ ICV_101 $T=0 281730 1 0 $X=-1000 $Y=277330
X18 VSS VDD WL1_120 WL0_120 WL0_119 WL1_119 WL1_118 WL0_118 WL0_117 WL1_117 XP2_7 XP2_6 XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_116
+ WL0_116 WL0_115 WL1_115 WL1_114 WL0_114 WL0_113 WL1_113 XP1_0 XP0_2 XP1_3 XP0_3
+ ICV_101 $T=0 390530 1 0 $X=-1000 $Y=386130
X19 VSS VDD WL1_16 WL0_16 WL0_15 WL1_15 WL1_14 WL0_14 WL0_13 WL1_13 WL1_12 WL0_12 WL0_11 WL1_11 WL1_10 WL0_10 WL0_9 WL1_9 XP2_7 XP2_6
+ XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_8 WL0_8 WL0_7 WL1_7 WL1_6 WL0_6 WL0_5 WL1_5 WL1_4 WL0_4 WL0_3 WL1_3 WL1_2
+ WL0_2 WL0_1 WL1_1 XP0_3 XP1_4 XP0_4 XP0_1 XP1_5 XP0_5
+ ICV_102 $T=0 9730 1 0 $X=-1000 $Y=5330
X20 VSS VDD WL1_48 WL0_48 WL0_47 WL1_47 WL1_46 WL0_46 WL0_45 WL1_45 WL1_44 WL0_44 WL0_43 WL1_43 WL1_42 WL0_42 WL0_41 WL1_41 XP2_7 XP2_6
+ XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_40 WL0_40 WL0_39 WL1_39 WL1_38 WL0_38 WL0_37 WL1_37 WL1_36 WL0_36 WL0_35 WL1_35 WL1_34
+ WL0_34 WL0_33 WL1_33 XP0_3 XP1_4 XP0_4 XP1_1 XP1_5 XP0_5
+ ICV_102 $T=0 118530 1 0 $X=-1000 $Y=114130
X21 VSS VDD WL1_80 WL0_80 WL0_79 WL1_79 WL1_78 WL0_78 WL0_77 WL1_77 WL1_76 WL0_76 WL0_75 WL1_75 WL1_74 WL0_74 WL0_73 WL1_73 XP2_7 XP2_6
+ XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_72 WL0_72 WL0_71 WL1_71 WL1_70 WL0_70 WL0_69 WL1_69 WL1_68 WL0_68 WL0_67 WL1_67 WL1_66
+ WL0_66 WL0_65 WL1_65 XP0_3 XP1_4 XP0_4 XP0_0 XP1_5 XP0_5
+ ICV_102 $T=0 227330 1 0 $X=-1000 $Y=222930
X22 VSS VDD WL1_112 WL0_112 WL0_111 WL1_111 WL1_110 WL0_110 WL0_109 WL1_109 WL1_108 WL0_108 WL0_107 WL1_107 WL1_106 WL0_106 WL0_105 WL1_105 XP2_7 XP2_6
+ XP2_5 XP2_4 XP2_3 XP2_2 XP2_1 XP2_0 GTP WL1_104 WL0_104 WL0_103 WL1_103 WL1_102 WL0_102 WL0_101 WL1_101 WL1_100 WL0_100 WL0_99 WL1_99 WL1_98
+ WL0_98 WL0_97 WL1_97 XP0_3 XP1_4 XP0_4 XP1_0 XP1_5 XP0_5
+ ICV_102 $T=0 336130 1 0 $X=-1000 $Y=331730
X24 VSS SIGN_MEMFLWDG1T $T=6800 2930 0 0 $X=5800 $Y=1930
X27 VSS VDD WL0_32 XP1_1 WL1_32 XP2_1 XP2_0 GTP XP0_5 SIGN_MEMROW_64 $T=0 111730 0 0 $X=-1000 $Y=110730
X28 VSS VDD WL0_64 XP0_0 WL1_64 XP2_1 XP2_0 GTP XP0_5 SIGN_MEMROW_64 $T=0 220530 0 0 $X=-1000 $Y=219530
X29 VSS VDD WL0_96 XP1_0 WL1_96 XP2_1 XP2_0 GTP XP0_5 SIGN_MEMROW_64 $T=0 329330 0 0 $X=-1000 $Y=328330
X30 VSS XP1_0 XP0_0 SIGN_MEMFCMWDX $T=0 438130 0 0 $X=-1000 $Y=437130
X31 VSS XP1_1 XP0_1 SIGN_MEMFCMWDX $T=3400 438130 0 0 $X=2400 $Y=437130
X32 VSS XP1_2 XP0_2 SIGN_MEMFCMWDX $T=6800 438130 0 0 $X=5800 $Y=437130
X33 VSS XP1_3 XP0_3 SIGN_MEMFCMWDX $T=10200 438130 0 0 $X=9200 $Y=437130
X34 VSS XP1_4 XP0_4 SIGN_MEMFCMWDX $T=13600 438130 0 0 $X=12600 $Y=437130
X35 VSS VDD XP0_1 WL0_0 WL1_0 XP2_1 XP2_0 GTP XP0_5 SIGN_MEMHWDB0 $T=20400 0 0 0 $X=19400 $Y=-1000
X36 VSS VDD MWL GTP MBL MWLD MBL_ SIGN_MEMMWDX $T=20400 438130 0 0 $X=19400 $Y=437130
.ENDS
***************************************
.SUBCKT SIGN_MEMHXP38X VSS VDD A2 A1 A0 XP_7 XP_6 XP_5 XP_4 XP_3 XP_2 XP_1 XP_0 BWEN AGTPB AGTPT
** N=41 EP=16 IP=109 FDC=348
*.CALIBRE ISOLATED NETS: WEI OEI_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 AY0 AY0_
M0 VSS VSS VSS VSS nfet L=9.2e-07 W=2.02e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1280 $Y=3380 $D=97
M1 VSS VSS VSS VSS nfet L=9.2e-07 W=2.03e-06 m=1 par=1 nf=1 ngcon=1 psp=0 $X=1280 $Y=6050 $D=97
X2 VSS A2 VDD 33 29 BWEN ai $T=6800 0 1 180 $X=2400 $Y=-1000
X3 VSS A1 VDD 32 31 BWEN ai $T=6800 0 0 0 $X=5800 $Y=-1000
X4 VSS A0 VDD 30 34 BWEN ai $T=13600 0 1 180 $X=9200 $Y=-1000
X5 VSS VDD XP_6 XP_7 AGTPB AGTPT 29 34 30 31 ap $T=0 9040 0 0 $X=-1000 $Y=8040
X6 VSS VDD XP_4 XP_5 AGTPB AGTPT 29 34 30 32 ap $T=6800 9040 1 180 $X=2400 $Y=8040
X7 VSS VDD XP_2 XP_3 AGTPB AGTPT 33 34 30 31 ap $T=6800 9040 0 0 $X=5800 $Y=8040
X8 VSS VDD XP_0 XP_1 AGTPB AGTPT 33 34 30 32 ap $T=13600 9040 1 180 $X=9200 $Y=8040
.ENDS
***************************************
.SUBCKT SIGN_MEMHYP38X VSS VDD A2 A1 A0 YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 BWEN AGTPB AGTPT
** N=27 EP=16 IP=104 FDC=346
*.CALIBRE ISOLATED NETS: WEI OEI_ AY0 AY0_
X0 VSS A2 VDD 25 21 BWEN ai $T=6800 0 1 180 $X=2400 $Y=-1000
X1 VSS A1 VDD 24 23 BWEN ai $T=6800 0 0 0 $X=5800 $Y=-1000
X2 VSS A0 VDD 22 26 BWEN ai $T=13600 0 1 180 $X=9200 $Y=-1000
X3 VSS VDD YP1_2 YP1_3 AGTPB AGTPT 21 26 22 23 ap $T=0 9040 0 0 $X=-1000 $Y=8040
X4 VSS VDD YP1_0 YP1_1 AGTPB AGTPT 21 26 22 24 ap $T=6800 9040 1 180 $X=2400 $Y=8040
X5 VSS VDD YP0_2 YP0_3 AGTPB AGTPT 25 26 22 23 ap $T=6800 9040 0 0 $X=5800 $Y=8040
X6 VSS VDD YP0_0 YP0_1 AGTPB AGTPT 25 26 22 24 ap $T=13600 9040 1 180 $X=9200 $Y=8040
.ENDS
***************************************
.SUBCKT SIGN_MEMHYP12RX VSS VDD A0 AY0 AY0_ AGTP BWEN
** N=24 EP=7 IP=28 FDC=90
*.CALIBRE ISOLATED NETS: WEI OEI_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GSRCN RST CLK GTPN
X0 VSS A0 VDD 22 23 BWEN ai $T=0 0 0 0 $X=-1000 $Y=-1000
X1 VSS VDD AY0 AY0_ AGTP AGTP VSS 22 23 VSS ap $T=0 9040 0 0 $X=-1000 $Y=8040
.ENDS
***************************************
.SUBCKT VPC_M1_CDNS_6479038850985
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT bf 1 2 3 4 5 6 7 8 9 10 11
** N=607 EP=11 IP=4 FDC=89
M0 19 2 20 2 lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1130 $Y=20160 $D=103
M1 18 13 2 2 lpnfet w=2.05e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1260 $Y=14610 $D=103
M2 20 12 19 2 lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1610 $Y=20160 $D=103
M3 2 13 18 2 lpnfet w=2.05e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1740 $Y=14610 $D=103
M4 2 17 19 2 lpnfet w=5.4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2120 $Y=19300 $D=103
M5 29 18 2 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2220 $Y=14460 $D=103
M6 27 8 20 2 lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2220 $Y=20540 $D=103
M7 2 16 27 2 lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2540 $Y=20540 $D=103
M8 5 24 29 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2620 $Y=14960 $D=103
M9 16 20 2 2 lpnfet w=8.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3060 $Y=19840 $D=103
M10 30 24 5 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3100 $Y=14960 $D=103
M11 2 3 12 2 lpnfet w=3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3440 $Y=6900 $D=103
M12 2 18 30 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3500 $Y=14540 $D=103
M13 31 18 2 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3980 $Y=14540 $D=103
M14 2 8 17 2 lpnfet w=9.2e-07 l=3.6e-07 m=1 par=1 nf=1 ngcon=1 $X=4040 $Y=19780 $D=103
M15 5 24 31 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4380 $Y=14960 $D=103
M16 32 17 2 2 lpnfet w=2.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4800 $Y=18600 $D=103
M17 33 24 5 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4860 $Y=14960 $D=103
M18 14 4 2 2 lpnfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4870 $Y=6070 $D=103
M19 10 16 32 2 lpnfet w=2.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5120 $Y=18600 $D=103
M20 2 18 33 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5260 $Y=14460 $D=103
M21 34 16 10 2 lpnfet w=2.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5600 $Y=18600 $D=103
M22 35 18 2 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5740 $Y=14460 $D=103
M23 2 17 34 2 lpnfet w=2.1e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5920 $Y=18600 $D=103
M24 5 24 35 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6140 $Y=14960 $D=103
M25 36 24 5 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6620 $Y=14960 $D=103
M26 37 8 22 2 lpnfet w=1.54e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6880 $Y=19070 $D=103
M27 2 18 36 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7020 $Y=14460 $D=103
M28 2 11 21 2 lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7070 $Y=7290 $D=103
M29 2 2 37 2 lpnfet w=1.54e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7200 $Y=19070 $D=103
M30 40 18 2 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7500 $Y=14460 $D=103
M31 38 23 2 2 lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7630 $Y=7170 $D=103
M32 39 6 2 2 lpnfet w=1.62e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7680 $Y=18990 $D=103
M33 5 24 40 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7900 $Y=14960 $D=103
M34 11 21 38 2 lpnfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7950 $Y=7170 $D=103
M35 13 22 39 2 lpnfet w=1.62e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8000 $Y=18990 $D=103
M36 41 24 5 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8380 $Y=14960 $D=103
M37 42 22 13 2 lpnfet w=1.62e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8480 $Y=18990 $D=103
M38 2 18 41 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8780 $Y=14460 $D=103
M39 2 6 42 2 lpnfet w=1.62e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8800 $Y=18990 $D=103
M40 43 18 2 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9260 $Y=14460 $D=103
M41 15 14 2 2 lpnfet w=2.02e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9320 $Y=18590 $D=103
M42 5 24 43 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9660 $Y=14960 $D=103
M43 44 24 5 2 lpnfet w=1.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10140 $Y=14960 $D=103
M44 2 18 44 2 lpnfet w=2.2e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10540 $Y=14460 $D=103
M45 7 15 2 2 lpnfet w=3.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10720 $Y=17720 $D=103
M46 24 9 2 2 lpnfet w=1.94e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11060 $Y=14720 $D=103
M47 2 15 7 2 lpnfet w=3.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=11200 $Y=17720 $D=103
M48 25 8 1 1 lppfet w=1.34e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1090 $Y=22030 $D=192
M49 26 2 25 1 lppfet w=1.34e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1410 $Y=22030 $D=192
M50 20 12 26 1 lppfet w=1.34e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1730 $Y=22030 $D=192
M51 18 13 1 1 lppfet w=2.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2000 $Y=10480 $D=192
M52 28 17 20 1 lppfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2330 $Y=22140 $D=192
M53 1 13 18 1 lppfet w=2.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2480 $Y=10480 $D=192
M54 1 16 28 1 lppfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2650 $Y=22140 $D=192
M55 18 13 1 1 lppfet w=2.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=2960 $Y=10480 $D=192
M56 16 20 1 1 lppfet w=1.62e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3170 $Y=21890 $D=192
M57 1 3 12 1 lppfet w=6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3440 $Y=7800 $D=192
M58 1 13 18 1 lppfet w=2.15e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=3440 $Y=10480 $D=192
M59 1 8 17 1 lppfet w=1.9e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4280 $Y=21890 $D=192
M60 5 18 1 1 lppfet w=3.44e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4380 $Y=9130 $D=192
M61 10 17 1 1 lppfet w=1.78e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4800 $Y=21890 $D=192
M62 1 18 5 1 lppfet w=3.44e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4860 $Y=9130 $D=192
M63 14 4 1 1 lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=4870 $Y=7570 $D=192
M64 1 17 10 1 lppfet w=1.78e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5280 $Y=21890 $D=192
M65 5 18 1 1 lppfet w=3.44e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5340 $Y=9130 $D=192
M66 1 4 14 1 lppfet w=9e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5350 $Y=7570 $D=192
M67 10 16 1 1 lppfet w=1.78e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5760 $Y=21890 $D=192
M68 1 18 5 1 lppfet w=3.44e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=5820 $Y=9130 $D=192
M69 1 16 10 1 lppfet w=1.78e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6240 $Y=21890 $D=192
M70 22 8 1 1 lppfet w=1.6e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6720 $Y=21890 $D=192
M71 5 24 1 1 lppfet w=2.4e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=6760 $Y=10230 $D=192
M72 1 11 21 1 lppfet w=3.2e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7070 $Y=8330 $D=192
M73 1 2 22 1 lppfet w=1.6e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7200 $Y=21890 $D=192
M74 11 21 1 1 lppfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7590 $Y=8330 $D=192
M75 13 6 1 1 lppfet w=1.72e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7700 $Y=21890 $D=192
M76 24 9 1 1 lppfet w=2.85e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=7920 $Y=9620 $D=192
M77 1 6 13 1 lppfet w=1.72e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8180 $Y=21890 $D=192
M78 1 9 24 1 lppfet w=2.85e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8400 $Y=9620 $D=192
M79 13 22 1 1 lppfet w=1.72e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8660 $Y=21890 $D=192
M80 7 15 1 1 lppfet w=3.01e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=8880 $Y=9620 $D=192
M81 1 22 13 1 lppfet w=1.72e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9140 $Y=21890 $D=192
M82 1 15 7 1 lppfet w=3.01e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9360 $Y=9620 $D=192
M83 15 14 1 1 lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9660 $Y=21890 $D=192
M84 23 23 1 1 lppfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9720 $Y=8670 $D=192
M85 7 15 1 1 lppfet w=3.01e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=9840 $Y=9620 $D=192
M86 1 14 15 1 lppfet w=2.12e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10140 $Y=21890 $D=192
M87 1 1 23 1 lppfet w=1.6e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10280 $Y=8550 $D=192
M88 1 15 7 1 lppfet w=3.01e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=10320 $Y=9620 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMHBFX VDD VSS CEN WEN CLK WEI RST GTP MBL GSRCN GTPN
** N=82 EP=11 IP=11 FDC=94
*.CALIBRE ISOLATED NETS: STUBWE
D0 VSS VSS tdndsx AREA=1.024e-13 perim=1.28e-06 $X=770 $Y=140 $D=558
D1 VSS CEN tdndsx AREA=1.024e-13 perim=1.28e-06 $X=3160 $Y=140 $D=558
D2 VSS WEN tdndsx AREA=1.024e-13 perim=1.28e-06 $X=8420 $Y=140 $D=558
D3 VSS VSS tdndsx AREA=1.024e-13 perim=1.28e-06 $X=10440 $Y=140 $D=558
D4 VSS CLK tdndsx AREA=1.024e-13 perim=1.28e-06 $X=12040 $Y=140 $D=558
X5 VDD VSS CEN WEN RST GTP WEI CLK MBL GSRCN GTPN bf $T=0 2500 0 0 $X=-1000 $Y=1500
.ENDS
***************************************
.SUBCKT SIGN_MEMCK VDD VSS GTPN GSRCN CLK RST GTP
** N=347 EP=7 IP=0 FDC=30
*.CALIBRE ISOLATED NETS: A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0
M0 84 GSRCN VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=3080 $D=103
M1 82 84 VSS VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=4410 $D=103
M2 83 CLK GTPN VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=9930 $D=103
M3 GTP GTPN VSS VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=30710 $D=103
M4 VSS GSRCN 84 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=3080 $D=103
M5 VSS 84 82 VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=4410 $D=103
M6 82 CLK 83 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=9930 $D=103
M7 VSS GTPN GTP VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=30710 $D=103
M8 84 GSRCN VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=3080 $D=103
M9 82 84 VSS VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=4410 $D=103
M10 83 CLK 82 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=9930 $D=103
M11 83 GTPN VDD VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=13880 $D=103
M12 GTP GTPN VSS VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=30710 $D=103
M13 VSS GSRCN 84 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=3080 $D=103
M14 VSS 84 82 VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=4410 $D=103
M15 GTPN CLK 83 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=9930 $D=103
M16 VDD GTPN 83 VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=13880 $D=103
M17 VSS GTPN GTP VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=30710 $D=103
M18 84 GSRCN VDD VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=1120 $D=192
M19 GTPN RST VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=15490 $D=192
M20 GTP GTPN VDD VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=19430 $D=192
M21 VDD GSRCN 84 VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=1120 $D=192
M22 VDD RST GTPN VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=15490 $D=192
M23 VDD GTPN GTP VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=19430 $D=192
M24 84 GSRCN VDD VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=1120 $D=192
M25 GTPN RST VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=15490 $D=192
M26 GTP GTPN VDD VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=19430 $D=192
M27 VDD GSRCN 84 VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=1120 $D=192
M28 VDD RST GTPN VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=15490 $D=192
M29 VDD GTPN GTP VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=19430 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEMCLK_DRVS VDD VSS GTPN GSRCN CLK RST AGTP GTP_0 GTP_1 GTP_2 GTP_3
** N=543 EP=11 IP=324 FDC=150
*.CALIBRE ISOLATED NETS: A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0
M0 24 GSRCN VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=3080 $D=103
M1 22 24 VSS VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=4410 $D=103
M2 23 CLK GTPN VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=9930 $D=103
M3 AGTP GTPN VSS VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=30710 $D=103
M4 VSS GSRCN 24 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=3080 $D=103
M5 VSS 24 22 VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=4410 $D=103
M6 22 CLK 23 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=9930 $D=103
M7 VSS GTPN AGTP VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=30710 $D=103
M8 24 GSRCN VSS VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=3080 $D=103
M9 22 24 VSS VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=4410 $D=103
M10 23 CLK 22 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=9930 $D=103
M11 23 GTPN VDD VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=13880 $D=103
M12 AGTP GTPN VSS VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=30710 $D=103
M13 VSS GSRCN 24 VSS lpnfet w=4e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=3080 $D=103
M14 VSS 24 22 VSS lpnfet w=4.7e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=4410 $D=103
M15 GTPN CLK 23 VSS lpnfet w=3.13e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=9930 $D=103
M16 VDD GTPN 23 VSS lpnfet w=8e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=13880 $D=103
M17 VSS GTPN AGTP VSS lpnfet w=2.8e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=30710 $D=103
M18 24 GSRCN VDD VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=1120 $D=192
M19 GTPN RST VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=15490 $D=192
M20 AGTP GTPN VDD VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=180 $Y=19430 $D=192
M21 VDD GSRCN 24 VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=1120 $D=192
M22 VDD RST GTPN VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=15490 $D=192
M23 VDD GTPN AGTP VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=660 $Y=19430 $D=192
M24 24 GSRCN VDD VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=1120 $D=192
M25 GTPN RST VDD VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=15490 $D=192
M26 AGTP GTPN VDD VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1140 $Y=19430 $D=192
M27 VDD GSRCN 24 VDD lppfet w=5.3e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=1120 $D=192
M28 VDD RST GTPN VDD lppfet w=3e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=15490 $D=192
M29 VDD GTPN AGTP VDD lppfet w=9.5e-06 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=1620 $Y=19430 $D=192
X30 VDD VSS GTPN GSRCN CLK RST GTP_0 SIGN_MEMCK $T=3840 0 1 180 $X=920 $Y=-1000
X31 VDD VSS GTPN GSRCN CLK RST GTP_1 SIGN_MEMCK $T=3840 0 0 0 $X=2840 $Y=-1000
X32 VDD VSS GTPN GSRCN CLK RST GTP_2 SIGN_MEMCK $T=7680 0 1 180 $X=4760 $Y=-1000
X33 VDD VSS GTPN GSRCN CLK RST GTP_3 SIGN_MEMCK $T=7680 0 0 0 $X=6680 $Y=-1000
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCCMBLST2 VSS 4
** N=7 EP=2 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD WL
M0 4 VSS VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1390 $D=103
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCCMBLST VSS WL NDL NDR WP
** N=9 EP=5 IP=0 FDC=2
*.CALIBRE ISOLATED NETS: VDD
M0 NDL WP VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=90 $Y=1390 $D=103
M1 NDR WL VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1390 $D=103
.ENDS
***************************************
.SUBCKT SIGN_MEMFLCCMBLSTU VSS WL 4
** N=7 EP=3 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD
M0 4 WL VSS VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=950 $Y=1390 $D=103
.ENDS
***************************************
.SUBCKT ICV_88 1 2 3 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 22
+ 24 26 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45
+ 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
** N=68 EP=55 IP=59 FDC=616
X0 1 3 4 2 22 28 26 24 17 18 19 20 7 6 8 9 10 11 12 13
+ 14 15 16 60 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44
+ 43 42 41 40 39 38 37 36 35 34 33 32 31 30 29
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_87
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_85 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_86
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_89 1 2 3 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 268 270 272 274 275 276 277 278 279 280 281 282 283 284 325
+ 356 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439
+ 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459
+ 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479
+ 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499
+ 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519
+ 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539
+ 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559
+ 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579
+ 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599
+ 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619
+ 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639
+ 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659
+ 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679
+ 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699
+ 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719
+ 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739
+ 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759
+ 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779
+ 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799
+ 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819
+ 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839
+ 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859
+ 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879
+ 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899
+ 900 901 902 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919
+ 920 921 922 923 924 925 926 927 928 929 930 931 932
** N=932 EP=793 IP=971 FDC=24680
*.SEEDPROM
X0 4 1 2 3 274 275 276 277 278 279 280 281 282 283 284 262 263 264 265 266
+ 268 270 272 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356
+ ICV_88 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 355 354
+ 353 352 351 350 349 348 347 346 345 344 343 342 341 340 339 338 337 336 335 334
+ 333 332 331 330 329 328 327 326 421 422 423 424 425 426 427 428 429 430 431 432
+ 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452
+ 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472
+ 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492
+ 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512
+ 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532
+ 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552
+ 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572
+ 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592
+ 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612
+ 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631 632
+ 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651 652
+ 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670 671 672
+ 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691 692
+ 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710 711 712
+ 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730 731 732
+ 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750 751 752
+ 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771 772
+ 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792
+ 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810 811 812
+ 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830 831 832
+ 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850 851 852
+ 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870 871 872
+ 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890 891 892
+ 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910 911 912
+ 913 914 915 916 917 918 919 920 921 922 923 924 925 926 927 928 929 930 931 932
+ ICV_85 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_83 1 2 3 4 5 6 7 8 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=59 EP=55 IP=59 FDC=616
X0 1 3 4 2 24 27 26 25 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_82
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_80 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_81
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_84 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 282 283 316
+ 347 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923
** N=923 EP=793 IP=961 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 273 274 275 276 277 278 279 280 281 282 283 266
+ 268 270 272 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ ICV_83 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 317 318
+ 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338
+ 339 340 341 342 343 344 345 346 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503
+ 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683
+ 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703
+ 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723
+ 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743
+ 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763
+ 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783
+ 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803
+ 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823
+ 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863
+ 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883
+ 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903
+ 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923
+ ICV_80 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_98 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -38400 0 270 $X=62320 $Y=-40600
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -38400 0 270 $X=89520 $Y=-40600
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -38400 0 270 $X=116720 $Y=-40600
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -38400 0 270 $X=143920 $Y=-40600
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -38400 0 270 $X=171120 $Y=-40600
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -38400 0 270 $X=198320 $Y=-40600
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -38400 0 270 $X=225520 $Y=-40600
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -38400 0 270 $X=252720 $Y=-40600
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -38400 0 270 $X=279920 $Y=-40600
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -38400 0 270 $X=307120 $Y=-40600
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -38400 0 270 $X=334320 $Y=-40600
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -38400 0 270 $X=361520 $Y=-40600
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -38400 0 270 $X=388720 $Y=-40600
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -38400 0 270 $X=415920 $Y=-40600
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -38400 0 270 $X=443120 $Y=-40600
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -38400 0 270 $X=470320 $Y=-40600
.ENDS
***************************************
.SUBCKT ICV_78 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=65 EP=55 IP=59 FDC=616
X0 1 3 4 2 9 12 11 10 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_77
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_75 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_76
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_79 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 267 269 271 273 274 275 276 277 278 279 280 281 282 283 316
+ 347 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923
** N=923 EP=793 IP=961 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 265 267 269 271 273 274 275 276 277 278 279 280
+ 281 282 283 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ ICV_78 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 346 345
+ 344 343 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326 325
+ 324 323 322 321 320 319 318 317 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503
+ 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683
+ 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703
+ 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723
+ 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743
+ 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763
+ 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783
+ 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803
+ 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823
+ 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863
+ 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883
+ 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903
+ 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923
+ ICV_75 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_73 1 2 3 4 5 6 7 8 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=59 EP=55 IP=59 FDC=616
X0 1 3 4 2 24 27 26 25 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_72
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_70 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_71
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_74 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 282 283 316
+ 347 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923
** N=923 EP=793 IP=961 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 273 274 275 276 277 278 279 280 281 282 283 266
+ 268 270 272 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ ICV_73 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 317 318
+ 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338
+ 339 340 341 342 343 344 345 346 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503
+ 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683
+ 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703
+ 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723
+ 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743
+ 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763
+ 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783
+ 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803
+ 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823
+ 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863
+ 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883
+ 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903
+ 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923
+ ICV_70 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_97 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -78000 0 270 $X=62320 $Y=-80200
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -78000 0 270 $X=89520 $Y=-80200
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -78000 0 270 $X=116720 $Y=-80200
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -78000 0 270 $X=143920 $Y=-80200
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -78000 0 270 $X=171120 $Y=-80200
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -78000 0 270 $X=198320 $Y=-80200
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -78000 0 270 $X=225520 $Y=-80200
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -78000 0 270 $X=252720 $Y=-80200
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -78000 0 270 $X=279920 $Y=-80200
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -78000 0 270 $X=307120 $Y=-80200
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -78000 0 270 $X=334320 $Y=-80200
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -78000 0 270 $X=361520 $Y=-80200
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -78000 0 270 $X=388720 $Y=-80200
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -78000 0 270 $X=415920 $Y=-80200
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -78000 0 270 $X=443120 $Y=-80200
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -78000 0 270 $X=470320 $Y=-80200
.ENDS
***************************************
.SUBCKT ICV_68 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=65 EP=55 IP=59 FDC=616
X0 1 3 4 2 9 12 11 10 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_67
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_65 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_66
** N=67 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 262 263 264 265 266 268 270 272 274 275 276 277 278 279 280 281 282 283 284 317
+ 348 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431
+ 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451
+ 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471
+ 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491
+ 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511
+ 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531
+ 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551
+ 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571
+ 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591
+ 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611
+ 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631
+ 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651
+ 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670 671
+ 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691
+ 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710 711
+ 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730 731
+ 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750 751
+ 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771
+ 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791
+ 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810 811
+ 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830 831
+ 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850 851
+ 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870 871
+ 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890 891
+ 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910 911
+ 912 913 914 915 916 917 918 919 920 921 922 923 924
** N=924 EP=793 IP=962 FDC=24680
*.SEEDPROM
X0 4 1 2 3 262 263 264 265 266 268 270 272 274 275 276 277 278 279 280 281
+ 282 283 284 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333
+ 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348
+ ICV_68 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 347 346
+ 345 344 343 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326
+ 325 324 323 322 321 320 319 318 413 414 415 416 417 418 419 420 421 422 423 424
+ 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444
+ 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464
+ 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484
+ 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504
+ 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524
+ 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544
+ 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564
+ 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584
+ 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604
+ 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624
+ 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644
+ 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664
+ 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683 684
+ 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703 704
+ 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724
+ 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743 744
+ 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763 764
+ 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783 784
+ 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803 804
+ 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823 824
+ 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843 844
+ 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863 864
+ 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883 884
+ 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903 904
+ 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923 924
+ ICV_65 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_63 1 2 3 4 5 6 7 8 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=59 EP=55 IP=59 FDC=616
X0 1 3 4 2 24 27 26 25 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_62 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_61
** N=35 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_56 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_59
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 266 268 270 272 273 274 275 276 277 278 279 280 281 282 283 316
+ 347 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923
** N=923 EP=793 IP=961 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 273 274 275 276 277 278 279 280 281 282 283 266
+ 268 270 272 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ ICV_63 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 317 318
+ 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338
+ 339 340 341 342 343 344 345 346 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503
+ 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683
+ 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703
+ 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723
+ 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743
+ 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763
+ 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783
+ 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803
+ 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823
+ 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863
+ 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883
+ 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903
+ 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923
+ ICV_57 $T=19200 63320 1 180 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_96 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
** N=258 EP=257 IP=288 FDC=512
X0 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_95 $T=63320 -117600 0 270 $X=62320 $Y=-119800
X1 1 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_95 $T=90520 -117600 0 270 $X=89520 $Y=-119800
X2 1 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 ICV_95 $T=117720 -117600 0 270 $X=116720 $Y=-119800
X3 1 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 ICV_95 $T=144920 -117600 0 270 $X=143920 $Y=-119800
X4 1 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 ICV_95 $T=172120 -117600 0 270 $X=171120 $Y=-119800
X5 1 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 ICV_95 $T=199320 -117600 0 270 $X=198320 $Y=-119800
X6 1 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 ICV_95 $T=226520 -117600 0 270 $X=225520 $Y=-119800
X7 1 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 ICV_95 $T=253720 -117600 0 270 $X=252720 $Y=-119800
X8 1 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 ICV_95 $T=280920 -117600 0 270 $X=279920 $Y=-119800
X9 1 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 ICV_95 $T=308120 -117600 0 270 $X=307120 $Y=-119800
X10 1 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 ICV_95 $T=335320 -117600 0 270 $X=334320 $Y=-119800
X11 1 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 ICV_95 $T=362520 -117600 0 270 $X=361520 $Y=-119800
X12 1 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 ICV_95 $T=389720 -117600 0 270 $X=388720 $Y=-119800
X13 1 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 ICV_95 $T=416920 -117600 0 270 $X=415920 $Y=-119800
X14 1 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 ICV_95 $T=444120 -117600 0 270 $X=443120 $Y=-119800
X15 1 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 ICV_95 $T=471320 -117600 0 270 $X=470320 $Y=-119800
.ENDS
***************************************
.SUBCKT ICV_54 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
** N=65 EP=55 IP=59 FDC=616
X0 1 3 4 2 9 12 11 10 5 6 7 8 14 13 15 16 17 18 19 20
+ 21 22 23 59 58 57 56 55 54 53 52 51 50 49 48 47 46 45 44 43
+ 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28
+ ICV_53 $T=0 0 0 0 $X=-1000 $Y=-20200
.ENDS
***************************************
.SUBCKT ICV_52
** N=36 EP=0 IP=34 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
** N=802 EP=800 IP=802 FDC=24064
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662
+ 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682
+ 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702
+ 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722
+ 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742
+ 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762
+ 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782
+ 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802
+ ICV_47 $T=0 0 0 0 $X=-1000 $Y=-1000
.ENDS
***************************************
.SUBCKT ICV_50
** N=66 EP=0 IP=66 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 267 269 271 273 274 275 276 277 278 279 280 281 282 283 316
+ 347 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530
+ 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550
+ 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570
+ 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590
+ 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923
** N=923 EP=793 IP=961 FDC=24680
*.SEEDPROM
X0 4 1 2 3 261 262 263 264 265 267 269 271 273 274 275 276 277 278 279 280
+ 281 282 283 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332
+ 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347
+ ICV_54 $T=0 0 0 90 $X=-1000 $Y=-1000
X2 4 2 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 346 345
+ 344 343 342 341 340 339 338 337 336 335 334 333 332 331 330 329 328 327 326 325
+ 324 323 322 321 320 319 318 317 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503
+ 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683
+ 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703
+ 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723
+ 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743
+ 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758 759 760 761 762 763
+ 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778 779 780 781 782 783
+ 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798 799 800 801 802 803
+ 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818 819 820 821 822 823
+ 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838 839 840 841 842 843
+ 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858 859 860 861 862 863
+ 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878 879 880 881 882 883
+ 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 903
+ 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 922 923
+ ICV_48 $T=0 63320 0 0 $X=-1000 $Y=62320
.ENDS
***************************************
.SUBCKT ICV_91 1 2 3 4 5 6 7 8 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56
** N=66 EP=55 IP=95 FDC=616
D0 1 3 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=140 $Y=-141760 $D=558
D1 1 4 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=140 $Y=-139360 $D=558
X2 1 2 57 5 6 58 4 59 21 22 23 3 SIGN_MEMIOX $T=1200 -147600 1 90 $X=200 $Y=-148600
X3 1 21 22 23 SIGN_MEMFLIO $T=1200 -157200 1 90 $X=200 $Y=-158200
X4 1 2 57 58 7 8 59 24 SIGN_MEMSA8 $T=12470 -147600 1 90 $X=11470 $Y=-148600
X5 1 24 SIGN_MEMFLSA $T=12470 -157200 1 90 $X=11470 $Y=-158200
X6 1 2 5 7 8 6 12 13 14 15 16 17 18 19 11 10 20 25 26 27
+ 28 33 34 35 36 41 42 43 44 49 50 51 52 32 31 30 29 40 39 38
+ 37 48 47 46 45 56 55 54 53
+ SIGN_MEMMUX_CD_ODD $T=22810 -157200 1 90 $X=21810 $Y=-158200
.ENDS
***************************************
.SUBCKT ICV_90 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 387 388 389 390 391 392 393 394 395 396 397 398
+ 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418
+ 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438
+ 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458
+ 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478
+ 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498
+ 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518
+ 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538
+ 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558
+ 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578
+ 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598
+ 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618
+ 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658
+ 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678
+ 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
+ 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718
+ 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738
+ 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758
+ 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778
+ 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798
+ 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878
+ 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898
** N=898 EP=800 IP=1158 FDC=24064
*.SEEDPROM
X1 1 2 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277
+ 278 279 280 281 282 283 284 285 286 287 288 289 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150
+ 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210
+ 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230
+ 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250
+ 251 252 253 254 255 256 257 258 387 388 389 390 391 392 393 394 395 396 397 398
+ 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418
+ 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438
+ 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458
+ 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478
+ 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498
+ 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518
+ 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538
+ 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558
+ 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578
+ 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598
+ 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618
+ 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658
+ 659 660 661 662 663 664 665 666 667 668 669 670 671 672 673 674 675 676 677 678
+ 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693 694 695 696 697 698
+ 699 700 701 702 703 704 705 706 707 708 709 710 711 712 713 714 715 716 717 718
+ 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734 735 736 737 738
+ 739 740 741 742 743 744 745 746 747 748 749 750 751 752 753 754 755 756 757 758
+ 759 760 761 762 763 764 765 766 767 768 769 770 771 772 773 774 775 776 777 778
+ 779 780 781 782 783 784 785 786 787 788 789 790 791 792 793 794 795 796 797 798
+ 799 800 801 802 803 804 805 806 807 808 809 810 811 812 813 814 815 816 817 818
+ 819 820 821 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837 838
+ 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 854 855 856 857 858
+ 859 860 861 862 863 864 865 866 867 868 869 870 871 872 873 874 875 876 877 878
+ 879 880 881 882 883 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898
+ SIGN_MEMBIT_COL $T=63320 -138000 0 270 $X=62320 $Y=-158200
.ENDS
***************************************
.SUBCKT SIGN_MEMWING_8_RIGHT VSS VDD D_0 Q_0 D_1 Q_1 D_2 Q_2 D_3 Q_3 D_4 Q_4 D_5 Q_5 D_6 Q_6 D_7 Q_7 WL_0 WL_1
+ WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 WL_20 WL_21
+ WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41
+ WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 WL_59 WL_60 WL_61
+ WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81
+ WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98 WL_99 WL_100 WL_101
+ WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 WL_119 WL_120 WL_121
+ WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138 WL_139 WL_140 WL_141
+ WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158 WL_159 WL_160 WL_161
+ WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178 WL_179 WL_180 WL_181
+ WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198 WL_199 WL_200 WL_201
+ WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218 WL_219 WL_220 WL_221
+ WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238 WL_239 WL_240 WL_241
+ WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0
+ YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 WE GTP_0 OE_ GTP_1 589 621 622 623 624 625 626 627 628 629 630
+ 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650
+ 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 666 667 668 669 670
+ 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690
+ 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705 706 707 708 709 710
+ 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725 726 727 728 729 730
+ 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745 746 747 748 749 750
+ 751 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770
+ 771 772 773 774 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790
+ 791 792 793 794 795 796 797 798 799 800 801 802 803 804 805 806 807 808 809 810
+ 811 812 813 814 815 816 817 818 819 820 821 822 823 824 825 826 827 828 829 830
+ 831 832 833 834 835 836 837 838 839 840 841 842 843 844 845 846 847 848 849 850
+ 851 852 853 854 855 856 857 858 859 860 861 862 863 864 865 866 867 868 869 870
+ 871 872 873 874 875 876 877 878 879 880 881 882 883 884 885 886 887 888 889 890
+ 891 892 893 894 895 896 897 898 899 900 901 902 903 904 905 906 907 908 909 910
+ 911 912 913 914 915 916 917 918 919 920 921 922 923 924 925 926 927 928 929 930
+ 931 932 933 934 935 936 937 938 939 940 941 942 943 944 945 946 947 948 949 950
+ 951 952 953 954 955 956 957 958 959 960 961 962 963 964 965 966 967 968 969 970
+ 971 972 973 974 975 976 977 978 979 980 981 982 983 984 985 986 987 988 989 990
+ 991 992 993 994 995 996 997 998 999 1000 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010
+ 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030
+ 1031 1032 1033 1034 1035 1036 1037 1038 1039 1040 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050
+ 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060 1061 1062 1063 1064 1065 1066 1067 1068 1069 1070
+ 1071 1072 1073 1074 1075 1076 1077 1078 1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089 1090
+ 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100 1101 1102 1103 1104 1105 1106 1107 1108 1109 1110
+ 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130
+ 1131 1132 1133
** N=4730 EP=803 IP=7477 FDC=202560
*.SEEDPROM
*.CALIBRE ISOLATED NETS: BLT_0 BLT__0 BLT_1 BLT__1 BLT_2 BLT__2 BLT_3 BLT__3 BLT_4 BLT__4 BLT_5 BLT__5 BLT_6 BLT__6 BLT_7 BLT__7 BLT_8 BLT__8 BLT_9 BLT__9
*+ BLT_10 BLT__10 BLT_11 BLT__11 BLT_12 BLT__12 BLT_13 BLT__13 BLT_14 BLT__14 BLT_15 BLT__15 BLT__31 BLT_31 BLT__30 BLT_30 BLT__29 BLT_29 BLT__28 BLT_28
*+ BLT__27 BLT_27 BLT__26 BLT_26 BLT__25 BLT_25 BLT__24 BLT_24 BLT__23 BLT_23 BLT__22 BLT_22 BLT__21 BLT_21 BLT__20 BLT_20 BLT__19 BLT_19 BLT__18 BLT_18
*+ BLT__17 BLT_17 BLT__16 BLT_16 BLT_32 BLT__32 BLT_33 BLT__33 BLT_34 BLT__34 BLT_35 BLT__35 BLT_36 BLT__36 BLT_37 BLT__37 BLT_38 BLT__38 BLT_39 BLT__39
*+ BLT_40 BLT__40 BLT_41 BLT__41 BLT_42 BLT__42 BLT_43 BLT__43 BLT_44 BLT__44 BLT_45 BLT__45 BLT_46 BLT__46 BLT_47 BLT__47 BLT__63 BLT_63 BLT__62 BLT_62
*+ BLT__61 BLT_61 BLT__60 BLT_60 BLT__59 BLT_59 BLT__58 BLT_58 BLT__57 BLT_57 BLT__56 BLT_56 BLT__55 BLT_55 BLT__54 BLT_54 BLT__53 BLT_53 BLT__52 BLT_52
*+ BLT__51 BLT_51 BLT__50 BLT_50 BLT__49 BLT_49 BLT__48 BLT_48 BLT_64 BLT__64 BLT_65 BLT__65 BLT_66 BLT__66 BLT_67 BLT__67 BLT_68 BLT__68 BLT_69 BLT__69
*+ BLT_70 BLT__70 BLT_71 BLT__71 BLT_72 BLT__72 BLT_73 BLT__73 BLT_74 BLT__74 BLT_75 BLT__75 BLT_76 BLT__76 BLT_77 BLT__77 BLT_78 BLT__78 BLT_79 BLT__79
*+ BLT__95 BLT_95 BLT__94 BLT_94 BLT__93 BLT_93 BLT__92 BLT_92 BLT__91 BLT_91 BLT__90 BLT_90 BLT__89 BLT_89 BLT__88 BLT_88 BLT__87 BLT_87 BLT__86 BLT_86
*+ BLT__85 BLT_85 BLT__84 BLT_84 BLT__83 BLT_83 BLT__82 BLT_82 BLT__81 BLT_81 BLT__80 BLT_80 BLT_96 BLT__96 BLT_97 BLT__97 BLT_98 BLT__98 BLT_99 BLT__99
*+ BLT_100 BLT__100 BLT_101 BLT__101 BLT_102 BLT__102 BLT_103 BLT__103 BLT_104 BLT__104 BLT_105 BLT__105 BLT_106 BLT__106 BLT_107 BLT__107 BLT_108 BLT__108 BLT_109 BLT__109
*+ BLT_110 BLT__110 BLT_111 BLT__111 STUBDR_0 BLT__127 BLT_127 BLT__126 BLT_126 BLT__125 BLT_125 BLT__124 BLT_124 BLT__123 BLT_123 BLT__122 BLT_122 BLT__121 BLT_121 BLT__120
*+ BLT_120 BLT__119 BLT_119 BLT__118 BLT_118 BLT__117 BLT_117 BLT__116 BLT_116 BLT__115 BLT_115 BLT__114 BLT_114 BLT__113 BLT_113 BLT__112 BLT_112
M0 1134 WL_0 1135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=64710 $D=103
M1 1136 WL_1 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=65200 $D=103
M2 1134 WL_2 1137 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=68110 $D=103
M3 1138 WL_3 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=68600 $D=103
M4 1134 WL_4 1139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=71510 $D=103
M5 1140 WL_5 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=72000 $D=103
M6 1134 WL_6 1141 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=74910 $D=103
M7 1142 WL_7 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=75400 $D=103
M8 1134 WL_8 1143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=78310 $D=103
M9 1144 WL_9 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=78800 $D=103
M10 1134 WL_10 1145 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=81710 $D=103
M11 1146 WL_11 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=82200 $D=103
M12 1134 WL_12 1147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=85110 $D=103
M13 1148 WL_13 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=85600 $D=103
M14 1134 WL_14 1149 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=88510 $D=103
M15 1150 WL_15 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=89000 $D=103
M16 1134 WL_16 1151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=91910 $D=103
M17 1152 WL_17 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=92400 $D=103
M18 1134 WL_18 1153 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=95310 $D=103
M19 1154 WL_19 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=95800 $D=103
M20 1134 WL_20 1155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=98710 $D=103
M21 1156 WL_21 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=99200 $D=103
M22 1134 WL_22 1157 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=102110 $D=103
M23 1158 WL_23 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=102600 $D=103
M24 1134 WL_24 1159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=105510 $D=103
M25 1160 WL_25 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=106000 $D=103
M26 1134 WL_26 1161 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=108910 $D=103
M27 1162 WL_27 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=109400 $D=103
M28 1134 WL_28 1163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=112310 $D=103
M29 1164 WL_29 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=112800 $D=103
M30 1134 WL_30 1165 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=115710 $D=103
M31 1166 WL_31 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=116200 $D=103
M32 1134 WL_32 1167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=119110 $D=103
M33 1168 WL_33 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=119600 $D=103
M34 1134 WL_34 1169 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=122510 $D=103
M35 1170 WL_35 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=123000 $D=103
M36 1134 WL_36 1171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=125910 $D=103
M37 1172 WL_37 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=126400 $D=103
M38 1134 WL_38 1173 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=129310 $D=103
M39 1174 WL_39 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=129800 $D=103
M40 1134 WL_40 1175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=132710 $D=103
M41 1176 WL_41 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=133200 $D=103
M42 1134 WL_42 1177 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=136110 $D=103
M43 1178 WL_43 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=136600 $D=103
M44 1134 WL_44 1179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=139510 $D=103
M45 1180 WL_45 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=140000 $D=103
M46 1134 WL_46 1181 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=142910 $D=103
M47 1182 WL_47 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=143400 $D=103
M48 1134 WL_48 1183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=146310 $D=103
M49 1184 WL_49 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=146800 $D=103
M50 1134 WL_50 1185 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=149710 $D=103
M51 1186 WL_51 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=150200 $D=103
M52 1134 WL_52 1187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=153110 $D=103
M53 1188 WL_53 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=153600 $D=103
M54 1134 WL_54 1189 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=156510 $D=103
M55 1190 WL_55 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=157000 $D=103
M56 1134 WL_56 1191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=159910 $D=103
M57 1192 WL_57 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=160400 $D=103
M58 1134 WL_58 1193 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=163310 $D=103
M59 1194 WL_59 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=163800 $D=103
M60 1134 WL_60 1195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=166710 $D=103
M61 1196 WL_61 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=167200 $D=103
M62 1134 WL_62 1197 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=170110 $D=103
M63 1198 WL_63 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=170600 $D=103
M64 1134 WL_64 1199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=173510 $D=103
M65 1200 WL_65 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=174000 $D=103
M66 1134 WL_66 1201 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=176910 $D=103
M67 1202 WL_67 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=177400 $D=103
M68 1134 WL_68 1203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=180310 $D=103
M69 1204 WL_69 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=180800 $D=103
M70 1134 WL_70 1205 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=183710 $D=103
M71 1206 WL_71 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=184200 $D=103
M72 1134 WL_72 1207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=187110 $D=103
M73 1208 WL_73 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=187600 $D=103
M74 1134 WL_74 1209 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=190510 $D=103
M75 1210 WL_75 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=191000 $D=103
M76 1134 WL_76 1211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=193910 $D=103
M77 1212 WL_77 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=194400 $D=103
M78 1134 WL_78 1213 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=197310 $D=103
M79 1214 WL_79 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=197800 $D=103
M80 1134 WL_80 1215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=200710 $D=103
M81 1216 WL_81 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=201200 $D=103
M82 1134 WL_82 1217 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=204110 $D=103
M83 1218 WL_83 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=204600 $D=103
M84 1134 WL_84 1219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=207510 $D=103
M85 1220 WL_85 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=208000 $D=103
M86 1134 WL_86 1221 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=210910 $D=103
M87 1222 WL_87 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=211400 $D=103
M88 1134 WL_88 1223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=214310 $D=103
M89 1224 WL_89 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=214800 $D=103
M90 1134 WL_90 1225 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=217710 $D=103
M91 1226 WL_91 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=218200 $D=103
M92 1134 WL_92 1227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=221110 $D=103
M93 1228 WL_93 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=221600 $D=103
M94 1134 WL_94 1229 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=224510 $D=103
M95 1230 WL_95 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=225000 $D=103
M96 1134 WL_96 1231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=227910 $D=103
M97 1232 WL_97 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=228400 $D=103
M98 1134 WL_98 1233 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=231310 $D=103
M99 1234 WL_99 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=231800 $D=103
M100 1134 WL_100 1235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=234710 $D=103
M101 1236 WL_101 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=235200 $D=103
M102 1134 WL_102 1237 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=238110 $D=103
M103 1238 WL_103 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=238600 $D=103
M104 1134 WL_104 1239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=241510 $D=103
M105 1240 WL_105 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=242000 $D=103
M106 1134 WL_106 1241 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=244910 $D=103
M107 1242 WL_107 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=245400 $D=103
M108 1134 WL_108 1243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=248310 $D=103
M109 1244 WL_109 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=248800 $D=103
M110 1134 WL_110 1245 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=251710 $D=103
M111 1246 WL_111 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=252200 $D=103
M112 1134 WL_112 1247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=255110 $D=103
M113 1248 WL_113 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=255600 $D=103
M114 1134 WL_114 1249 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=258510 $D=103
M115 1250 WL_115 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=259000 $D=103
M116 1134 WL_116 1251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=261910 $D=103
M117 1252 WL_117 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=262400 $D=103
M118 1134 WL_118 1253 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=265310 $D=103
M119 1254 WL_119 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=265800 $D=103
M120 1134 WL_120 1255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=268710 $D=103
M121 1256 WL_121 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=269200 $D=103
M122 1134 WL_122 1257 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=272110 $D=103
M123 1258 WL_123 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=272600 $D=103
M124 1134 WL_124 1259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=275510 $D=103
M125 1260 WL_125 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=276000 $D=103
M126 1134 WL_126 1261 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=278910 $D=103
M127 1262 WL_127 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=279400 $D=103
M128 1134 WL_128 1263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=282310 $D=103
M129 1264 WL_129 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=282800 $D=103
M130 1134 WL_130 1265 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=285710 $D=103
M131 1266 WL_131 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=286200 $D=103
M132 1134 WL_132 1267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=289110 $D=103
M133 1268 WL_133 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=289600 $D=103
M134 1134 WL_134 1269 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=292510 $D=103
M135 1270 WL_135 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=293000 $D=103
M136 1134 WL_136 1271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=295910 $D=103
M137 1272 WL_137 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=296400 $D=103
M138 1134 WL_138 1273 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=299310 $D=103
M139 1274 WL_139 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=299800 $D=103
M140 1134 WL_140 1275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=302710 $D=103
M141 1276 WL_141 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=303200 $D=103
M142 1134 WL_142 1277 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=306110 $D=103
M143 1278 WL_143 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=306600 $D=103
M144 1134 WL_144 1279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=309510 $D=103
M145 1280 WL_145 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=310000 $D=103
M146 1134 WL_146 1281 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=312910 $D=103
M147 1282 WL_147 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=313400 $D=103
M148 1134 WL_148 1283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=316310 $D=103
M149 1284 WL_149 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=316800 $D=103
M150 1134 WL_150 1285 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=319710 $D=103
M151 1286 WL_151 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=320200 $D=103
M152 1134 WL_152 1287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=323110 $D=103
M153 1288 WL_153 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=323600 $D=103
M154 1134 WL_154 1289 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=326510 $D=103
M155 1290 WL_155 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=327000 $D=103
M156 1134 WL_156 1291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=329910 $D=103
M157 1292 WL_157 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=330400 $D=103
M158 1134 WL_158 1293 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=333310 $D=103
M159 1294 WL_159 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=333800 $D=103
M160 1134 WL_160 1295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=336710 $D=103
M161 1296 WL_161 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=337200 $D=103
M162 1134 WL_162 1297 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=340110 $D=103
M163 1298 WL_163 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=340600 $D=103
M164 1134 WL_164 1299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=343510 $D=103
M165 1300 WL_165 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=344000 $D=103
M166 1134 WL_166 1301 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=346910 $D=103
M167 1302 WL_167 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=347400 $D=103
M168 1134 WL_168 1303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=350310 $D=103
M169 1304 WL_169 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=350800 $D=103
M170 1134 WL_170 1305 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=353710 $D=103
M171 1306 WL_171 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=354200 $D=103
M172 1134 WL_172 1307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=357110 $D=103
M173 1308 WL_173 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=357600 $D=103
M174 1134 WL_174 1309 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=360510 $D=103
M175 1310 WL_175 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=361000 $D=103
M176 1134 WL_176 1311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=363910 $D=103
M177 1312 WL_177 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=364400 $D=103
M178 1134 WL_178 1313 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=367310 $D=103
M179 1314 WL_179 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=367800 $D=103
M180 1134 WL_180 1315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=370710 $D=103
M181 1316 WL_181 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=371200 $D=103
M182 1134 WL_182 1317 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=374110 $D=103
M183 1318 WL_183 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=374600 $D=103
M184 1134 WL_184 1319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=377510 $D=103
M185 1320 WL_185 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=378000 $D=103
M186 1134 WL_186 1321 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=380910 $D=103
M187 1322 WL_187 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=381400 $D=103
M188 1134 WL_188 1323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=384310 $D=103
M189 1324 WL_189 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=384800 $D=103
M190 1134 WL_190 1325 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=387710 $D=103
M191 1326 WL_191 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=388200 $D=103
M192 1134 WL_192 1327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=391110 $D=103
M193 1328 WL_193 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=391600 $D=103
M194 1134 WL_194 1329 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=394510 $D=103
M195 1330 WL_195 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=395000 $D=103
M196 1134 WL_196 1331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=397910 $D=103
M197 1332 WL_197 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=398400 $D=103
M198 1134 WL_198 1333 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=401310 $D=103
M199 1334 WL_199 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=401800 $D=103
M200 1134 WL_200 1335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=404710 $D=103
M201 1336 WL_201 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=405200 $D=103
M202 1134 WL_202 1337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=408110 $D=103
M203 1338 WL_203 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=408600 $D=103
M204 1134 WL_204 1339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=411510 $D=103
M205 1340 WL_205 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=412000 $D=103
M206 1134 WL_206 1341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=414910 $D=103
M207 1342 WL_207 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=415400 $D=103
M208 1134 WL_208 1343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=418310 $D=103
M209 1344 WL_209 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=418800 $D=103
M210 1134 WL_210 1345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=421710 $D=103
M211 1346 WL_211 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=422200 $D=103
M212 1134 WL_212 1347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=425110 $D=103
M213 1348 WL_213 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=425600 $D=103
M214 1134 WL_214 1349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=428510 $D=103
M215 1350 WL_215 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=429000 $D=103
M216 1134 WL_216 1351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=431910 $D=103
M217 1352 WL_217 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=432400 $D=103
M218 1134 WL_218 1353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=435310 $D=103
M219 1354 WL_219 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=435800 $D=103
M220 1134 WL_220 1355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=438710 $D=103
M221 1356 WL_221 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=439200 $D=103
M222 1134 WL_222 1357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=442110 $D=103
M223 1358 WL_223 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=442600 $D=103
M224 1134 WL_224 1359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=445510 $D=103
M225 1360 WL_225 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=446000 $D=103
M226 1134 WL_226 1361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=448910 $D=103
M227 1362 WL_227 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=449400 $D=103
M228 1134 WL_228 1363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=452310 $D=103
M229 1364 WL_229 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=452800 $D=103
M230 1134 WL_230 1365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=455710 $D=103
M231 1366 WL_231 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=456200 $D=103
M232 1134 WL_232 1367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=459110 $D=103
M233 1368 WL_233 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=459600 $D=103
M234 1134 WL_234 1369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=462510 $D=103
M235 1370 WL_235 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=463000 $D=103
M236 1134 WL_236 1371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=465910 $D=103
M237 1372 WL_237 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=466400 $D=103
M238 1134 WL_238 1373 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=469310 $D=103
M239 1374 WL_239 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=469800 $D=103
M240 1134 WL_240 1375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=472710 $D=103
M241 1376 WL_241 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=473200 $D=103
M242 1134 WL_242 1377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=476110 $D=103
M243 1378 WL_243 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=476600 $D=103
M244 1134 WL_244 1379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=479510 $D=103
M245 1380 WL_245 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=480000 $D=103
M246 1134 WL_246 1381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=482910 $D=103
M247 1382 WL_247 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=483400 $D=103
M248 1134 WL_248 1383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=486310 $D=103
M249 1384 WL_249 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=486800 $D=103
M250 1134 WL_250 1385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=489710 $D=103
M251 1386 WL_251 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=490200 $D=103
M252 1134 WL_252 1387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=493110 $D=103
M253 1388 WL_253 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=493600 $D=103
M254 1134 WL_254 1389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=496510 $D=103
M255 1390 WL_255 1134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18950 $Y=497000 $D=103
M256 1391 WL_0 1393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=64710 $D=103
M257 1395 WL_1 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=65200 $D=103
M258 1391 WL_2 1397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=68110 $D=103
M259 1399 WL_3 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=68600 $D=103
M260 1391 WL_4 1401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=71510 $D=103
M261 1403 WL_5 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=72000 $D=103
M262 1391 WL_6 1405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=74910 $D=103
M263 1407 WL_7 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=75400 $D=103
M264 1391 WL_8 1409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=78310 $D=103
M265 1411 WL_9 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=78800 $D=103
M266 1391 WL_10 1413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=81710 $D=103
M267 1415 WL_11 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=82200 $D=103
M268 1391 WL_12 1417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=85110 $D=103
M269 1419 WL_13 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=85600 $D=103
M270 1391 WL_14 1421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=88510 $D=103
M271 1423 WL_15 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=89000 $D=103
M272 1391 WL_16 1425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=91910 $D=103
M273 1427 WL_17 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=92400 $D=103
M274 1391 WL_18 1429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=95310 $D=103
M275 1431 WL_19 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=95800 $D=103
M276 1391 WL_20 1433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=98710 $D=103
M277 1435 WL_21 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=99200 $D=103
M278 1391 WL_22 1437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=102110 $D=103
M279 1439 WL_23 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=102600 $D=103
M280 1391 WL_24 1441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=105510 $D=103
M281 1443 WL_25 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=106000 $D=103
M282 1391 WL_26 1445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=108910 $D=103
M283 1447 WL_27 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=109400 $D=103
M284 1391 WL_28 1449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=112310 $D=103
M285 1451 WL_29 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=112800 $D=103
M286 1391 WL_30 1453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=115710 $D=103
M287 1455 WL_31 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=116200 $D=103
M288 1391 WL_32 1457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=119110 $D=103
M289 1459 WL_33 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=119600 $D=103
M290 1391 WL_34 1461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=122510 $D=103
M291 1463 WL_35 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=123000 $D=103
M292 1391 WL_36 1465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=125910 $D=103
M293 1467 WL_37 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=126400 $D=103
M294 1391 WL_38 1469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=129310 $D=103
M295 1471 WL_39 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=129800 $D=103
M296 1391 WL_40 1473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=132710 $D=103
M297 1475 WL_41 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=133200 $D=103
M298 1391 WL_42 1477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=136110 $D=103
M299 1479 WL_43 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=136600 $D=103
M300 1391 WL_44 1481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=139510 $D=103
M301 1483 WL_45 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=140000 $D=103
M302 1391 WL_46 1485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=142910 $D=103
M303 1487 WL_47 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=143400 $D=103
M304 1391 WL_48 1489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=146310 $D=103
M305 1491 WL_49 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=146800 $D=103
M306 1391 WL_50 1493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=149710 $D=103
M307 1495 WL_51 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=150200 $D=103
M308 1391 WL_52 1497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=153110 $D=103
M309 1499 WL_53 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=153600 $D=103
M310 1391 WL_54 1501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=156510 $D=103
M311 1503 WL_55 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=157000 $D=103
M312 1391 WL_56 1505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=159910 $D=103
M313 1507 WL_57 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=160400 $D=103
M314 1391 WL_58 1509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=163310 $D=103
M315 1511 WL_59 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=163800 $D=103
M316 1391 WL_60 1513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=166710 $D=103
M317 1515 WL_61 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=167200 $D=103
M318 1391 WL_62 1517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=170110 $D=103
M319 1519 WL_63 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=170600 $D=103
M320 1391 WL_64 1521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=173510 $D=103
M321 1523 WL_65 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=174000 $D=103
M322 1391 WL_66 1525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=176910 $D=103
M323 1527 WL_67 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=177400 $D=103
M324 1391 WL_68 1529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=180310 $D=103
M325 1531 WL_69 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=180800 $D=103
M326 1391 WL_70 1533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=183710 $D=103
M327 1535 WL_71 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=184200 $D=103
M328 1391 WL_72 1537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=187110 $D=103
M329 1539 WL_73 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=187600 $D=103
M330 1391 WL_74 1541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=190510 $D=103
M331 1543 WL_75 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=191000 $D=103
M332 1391 WL_76 1545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=193910 $D=103
M333 1547 WL_77 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=194400 $D=103
M334 1391 WL_78 1549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=197310 $D=103
M335 1551 WL_79 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=197800 $D=103
M336 1391 WL_80 1553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=200710 $D=103
M337 1555 WL_81 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=201200 $D=103
M338 1391 WL_82 1557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=204110 $D=103
M339 1559 WL_83 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=204600 $D=103
M340 1391 WL_84 1561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=207510 $D=103
M341 1563 WL_85 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=208000 $D=103
M342 1391 WL_86 1565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=210910 $D=103
M343 1567 WL_87 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=211400 $D=103
M344 1391 WL_88 1569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=214310 $D=103
M345 1571 WL_89 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=214800 $D=103
M346 1391 WL_90 1573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=217710 $D=103
M347 1575 WL_91 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=218200 $D=103
M348 1391 WL_92 1577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=221110 $D=103
M349 1579 WL_93 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=221600 $D=103
M350 1391 WL_94 1581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=224510 $D=103
M351 1583 WL_95 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=225000 $D=103
M352 1391 WL_96 1585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=227910 $D=103
M353 1587 WL_97 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=228400 $D=103
M354 1391 WL_98 1589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=231310 $D=103
M355 1591 WL_99 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=231800 $D=103
M356 1391 WL_100 1593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=234710 $D=103
M357 1595 WL_101 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=235200 $D=103
M358 1391 WL_102 1597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=238110 $D=103
M359 1599 WL_103 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=238600 $D=103
M360 1391 WL_104 1601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=241510 $D=103
M361 1603 WL_105 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=242000 $D=103
M362 1391 WL_106 1605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=244910 $D=103
M363 1607 WL_107 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=245400 $D=103
M364 1391 WL_108 1609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=248310 $D=103
M365 1611 WL_109 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=248800 $D=103
M366 1391 WL_110 1613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=251710 $D=103
M367 1615 WL_111 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=252200 $D=103
M368 1391 WL_112 1617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=255110 $D=103
M369 1619 WL_113 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=255600 $D=103
M370 1391 WL_114 1621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=258510 $D=103
M371 1623 WL_115 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=259000 $D=103
M372 1391 WL_116 1625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=261910 $D=103
M373 1627 WL_117 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=262400 $D=103
M374 1391 WL_118 1629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=265310 $D=103
M375 1631 WL_119 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=265800 $D=103
M376 1391 WL_120 1633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=268710 $D=103
M377 1635 WL_121 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=269200 $D=103
M378 1391 WL_122 1637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=272110 $D=103
M379 1639 WL_123 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=272600 $D=103
M380 1391 WL_124 1641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=275510 $D=103
M381 1643 WL_125 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=276000 $D=103
M382 1391 WL_126 1645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=278910 $D=103
M383 1647 WL_127 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=279400 $D=103
M384 1391 WL_128 1649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=282310 $D=103
M385 1651 WL_129 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=282800 $D=103
M386 1391 WL_130 1653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=285710 $D=103
M387 1655 WL_131 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=286200 $D=103
M388 1391 WL_132 1657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=289110 $D=103
M389 1659 WL_133 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=289600 $D=103
M390 1391 WL_134 1661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=292510 $D=103
M391 1663 WL_135 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=293000 $D=103
M392 1391 WL_136 1665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=295910 $D=103
M393 1667 WL_137 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=296400 $D=103
M394 1391 WL_138 1669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=299310 $D=103
M395 1671 WL_139 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=299800 $D=103
M396 1391 WL_140 1673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=302710 $D=103
M397 1675 WL_141 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=303200 $D=103
M398 1391 WL_142 1677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=306110 $D=103
M399 1679 WL_143 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=306600 $D=103
M400 1391 WL_144 1681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=309510 $D=103
M401 1683 WL_145 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=310000 $D=103
M402 1391 WL_146 1685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=312910 $D=103
M403 1687 WL_147 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=313400 $D=103
M404 1391 WL_148 1689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=316310 $D=103
M405 1691 WL_149 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=316800 $D=103
M406 1391 WL_150 1693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=319710 $D=103
M407 1695 WL_151 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=320200 $D=103
M408 1391 WL_152 1697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=323110 $D=103
M409 1699 WL_153 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=323600 $D=103
M410 1391 WL_154 1701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=326510 $D=103
M411 1703 WL_155 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=327000 $D=103
M412 1391 WL_156 1705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=329910 $D=103
M413 1707 WL_157 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=330400 $D=103
M414 1391 WL_158 1709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=333310 $D=103
M415 1711 WL_159 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=333800 $D=103
M416 1391 WL_160 1713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=336710 $D=103
M417 1715 WL_161 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=337200 $D=103
M418 1391 WL_162 1717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=340110 $D=103
M419 1719 WL_163 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=340600 $D=103
M420 1391 WL_164 1721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=343510 $D=103
M421 1723 WL_165 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=344000 $D=103
M422 1391 WL_166 1725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=346910 $D=103
M423 1727 WL_167 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=347400 $D=103
M424 1391 WL_168 1729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=350310 $D=103
M425 1731 WL_169 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=350800 $D=103
M426 1391 WL_170 1733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=353710 $D=103
M427 1735 WL_171 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=354200 $D=103
M428 1391 WL_172 1737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=357110 $D=103
M429 1739 WL_173 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=357600 $D=103
M430 1391 WL_174 1741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=360510 $D=103
M431 1743 WL_175 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=361000 $D=103
M432 1391 WL_176 1745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=363910 $D=103
M433 1747 WL_177 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=364400 $D=103
M434 1391 WL_178 1749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=367310 $D=103
M435 1751 WL_179 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=367800 $D=103
M436 1391 WL_180 1753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=370710 $D=103
M437 1755 WL_181 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=371200 $D=103
M438 1391 WL_182 1757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=374110 $D=103
M439 1759 WL_183 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=374600 $D=103
M440 1391 WL_184 1761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=377510 $D=103
M441 1763 WL_185 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=378000 $D=103
M442 1391 WL_186 1765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=380910 $D=103
M443 1767 WL_187 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=381400 $D=103
M444 1391 WL_188 1769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=384310 $D=103
M445 1771 WL_189 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=384800 $D=103
M446 1391 WL_190 1773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=387710 $D=103
M447 1775 WL_191 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=388200 $D=103
M448 1391 WL_192 1777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=391110 $D=103
M449 1779 WL_193 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=391600 $D=103
M450 1391 WL_194 1781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=394510 $D=103
M451 1783 WL_195 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=395000 $D=103
M452 1391 WL_196 1785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=397910 $D=103
M453 1787 WL_197 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=398400 $D=103
M454 1391 WL_198 1789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=401310 $D=103
M455 1791 WL_199 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=401800 $D=103
M456 1391 WL_200 1793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=404710 $D=103
M457 1795 WL_201 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=405200 $D=103
M458 1391 WL_202 1797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=408110 $D=103
M459 1799 WL_203 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=408600 $D=103
M460 1391 WL_204 1801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=411510 $D=103
M461 1803 WL_205 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=412000 $D=103
M462 1391 WL_206 1805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=414910 $D=103
M463 1807 WL_207 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=415400 $D=103
M464 1391 WL_208 1809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=418310 $D=103
M465 1811 WL_209 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=418800 $D=103
M466 1391 WL_210 1813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=421710 $D=103
M467 1815 WL_211 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=422200 $D=103
M468 1391 WL_212 1817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=425110 $D=103
M469 1819 WL_213 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=425600 $D=103
M470 1391 WL_214 1821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=428510 $D=103
M471 1823 WL_215 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=429000 $D=103
M472 1391 WL_216 1825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=431910 $D=103
M473 1827 WL_217 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=432400 $D=103
M474 1391 WL_218 1829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=435310 $D=103
M475 1831 WL_219 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=435800 $D=103
M476 1391 WL_220 1833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=438710 $D=103
M477 1835 WL_221 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=439200 $D=103
M478 1391 WL_222 1837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=442110 $D=103
M479 1839 WL_223 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=442600 $D=103
M480 1391 WL_224 1841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=445510 $D=103
M481 1843 WL_225 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=446000 $D=103
M482 1391 WL_226 1845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=448910 $D=103
M483 1847 WL_227 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=449400 $D=103
M484 1391 WL_228 1849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=452310 $D=103
M485 1851 WL_229 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=452800 $D=103
M486 1391 WL_230 1853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=455710 $D=103
M487 1855 WL_231 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=456200 $D=103
M488 1391 WL_232 1857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=459110 $D=103
M489 1859 WL_233 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=459600 $D=103
M490 1391 WL_234 1861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=462510 $D=103
M491 1863 WL_235 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=463000 $D=103
M492 1391 WL_236 1865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=465910 $D=103
M493 1867 WL_237 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=466400 $D=103
M494 1391 WL_238 1869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=469310 $D=103
M495 1871 WL_239 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=469800 $D=103
M496 1391 WL_240 1873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=472710 $D=103
M497 1875 WL_241 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=473200 $D=103
M498 1391 WL_242 1877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=476110 $D=103
M499 1879 WL_243 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=476600 $D=103
M500 1391 WL_244 1881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=479510 $D=103
M501 1883 WL_245 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=480000 $D=103
M502 1391 WL_246 1885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=482910 $D=103
M503 1887 WL_247 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=483400 $D=103
M504 1391 WL_248 1889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=486310 $D=103
M505 1891 WL_249 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=486800 $D=103
M506 1391 WL_250 1893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=489710 $D=103
M507 1895 WL_251 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=490200 $D=103
M508 1391 WL_252 1897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=493110 $D=103
M509 1899 WL_253 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=493600 $D=103
M510 1391 WL_254 1901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=496510 $D=103
M511 1903 WL_255 1391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19290 $Y=497000 $D=103
M512 1392 WL_0 1394 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=64710 $D=103
M513 1396 WL_1 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=65200 $D=103
M514 1392 WL_2 1398 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=68110 $D=103
M515 1400 WL_3 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=68600 $D=103
M516 1392 WL_4 1402 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=71510 $D=103
M517 1404 WL_5 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=72000 $D=103
M518 1392 WL_6 1406 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=74910 $D=103
M519 1408 WL_7 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=75400 $D=103
M520 1392 WL_8 1410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=78310 $D=103
M521 1412 WL_9 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=78800 $D=103
M522 1392 WL_10 1414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=81710 $D=103
M523 1416 WL_11 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=82200 $D=103
M524 1392 WL_12 1418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=85110 $D=103
M525 1420 WL_13 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=85600 $D=103
M526 1392 WL_14 1422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=88510 $D=103
M527 1424 WL_15 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=89000 $D=103
M528 1392 WL_16 1426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=91910 $D=103
M529 1428 WL_17 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=92400 $D=103
M530 1392 WL_18 1430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=95310 $D=103
M531 1432 WL_19 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=95800 $D=103
M532 1392 WL_20 1434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=98710 $D=103
M533 1436 WL_21 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=99200 $D=103
M534 1392 WL_22 1438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=102110 $D=103
M535 1440 WL_23 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=102600 $D=103
M536 1392 WL_24 1442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=105510 $D=103
M537 1444 WL_25 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=106000 $D=103
M538 1392 WL_26 1446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=108910 $D=103
M539 1448 WL_27 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=109400 $D=103
M540 1392 WL_28 1450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=112310 $D=103
M541 1452 WL_29 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=112800 $D=103
M542 1392 WL_30 1454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=115710 $D=103
M543 1456 WL_31 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=116200 $D=103
M544 1392 WL_32 1458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=119110 $D=103
M545 1460 WL_33 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=119600 $D=103
M546 1392 WL_34 1462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=122510 $D=103
M547 1464 WL_35 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=123000 $D=103
M548 1392 WL_36 1466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=125910 $D=103
M549 1468 WL_37 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=126400 $D=103
M550 1392 WL_38 1470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=129310 $D=103
M551 1472 WL_39 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=129800 $D=103
M552 1392 WL_40 1474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=132710 $D=103
M553 1476 WL_41 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=133200 $D=103
M554 1392 WL_42 1478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=136110 $D=103
M555 1480 WL_43 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=136600 $D=103
M556 1392 WL_44 1482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=139510 $D=103
M557 1484 WL_45 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=140000 $D=103
M558 1392 WL_46 1486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=142910 $D=103
M559 1488 WL_47 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=143400 $D=103
M560 1392 WL_48 1490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=146310 $D=103
M561 1492 WL_49 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=146800 $D=103
M562 1392 WL_50 1494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=149710 $D=103
M563 1496 WL_51 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=150200 $D=103
M564 1392 WL_52 1498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=153110 $D=103
M565 1500 WL_53 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=153600 $D=103
M566 1392 WL_54 1502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=156510 $D=103
M567 1504 WL_55 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=157000 $D=103
M568 1392 WL_56 1506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=159910 $D=103
M569 1508 WL_57 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=160400 $D=103
M570 1392 WL_58 1510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=163310 $D=103
M571 1512 WL_59 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=163800 $D=103
M572 1392 WL_60 1514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=166710 $D=103
M573 1516 WL_61 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=167200 $D=103
M574 1392 WL_62 1518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=170110 $D=103
M575 1520 WL_63 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=170600 $D=103
M576 1392 WL_64 1522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=173510 $D=103
M577 1524 WL_65 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=174000 $D=103
M578 1392 WL_66 1526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=176910 $D=103
M579 1528 WL_67 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=177400 $D=103
M580 1392 WL_68 1530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=180310 $D=103
M581 1532 WL_69 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=180800 $D=103
M582 1392 WL_70 1534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=183710 $D=103
M583 1536 WL_71 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=184200 $D=103
M584 1392 WL_72 1538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=187110 $D=103
M585 1540 WL_73 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=187600 $D=103
M586 1392 WL_74 1542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=190510 $D=103
M587 1544 WL_75 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=191000 $D=103
M588 1392 WL_76 1546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=193910 $D=103
M589 1548 WL_77 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=194400 $D=103
M590 1392 WL_78 1550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=197310 $D=103
M591 1552 WL_79 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=197800 $D=103
M592 1392 WL_80 1554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=200710 $D=103
M593 1556 WL_81 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=201200 $D=103
M594 1392 WL_82 1558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=204110 $D=103
M595 1560 WL_83 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=204600 $D=103
M596 1392 WL_84 1562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=207510 $D=103
M597 1564 WL_85 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=208000 $D=103
M598 1392 WL_86 1566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=210910 $D=103
M599 1568 WL_87 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=211400 $D=103
M600 1392 WL_88 1570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=214310 $D=103
M601 1572 WL_89 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=214800 $D=103
M602 1392 WL_90 1574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=217710 $D=103
M603 1576 WL_91 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=218200 $D=103
M604 1392 WL_92 1578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=221110 $D=103
M605 1580 WL_93 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=221600 $D=103
M606 1392 WL_94 1582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=224510 $D=103
M607 1584 WL_95 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=225000 $D=103
M608 1392 WL_96 1586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=227910 $D=103
M609 1588 WL_97 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=228400 $D=103
M610 1392 WL_98 1590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=231310 $D=103
M611 1592 WL_99 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=231800 $D=103
M612 1392 WL_100 1594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=234710 $D=103
M613 1596 WL_101 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=235200 $D=103
M614 1392 WL_102 1598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=238110 $D=103
M615 1600 WL_103 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=238600 $D=103
M616 1392 WL_104 1602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=241510 $D=103
M617 1604 WL_105 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=242000 $D=103
M618 1392 WL_106 1606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=244910 $D=103
M619 1608 WL_107 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=245400 $D=103
M620 1392 WL_108 1610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=248310 $D=103
M621 1612 WL_109 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=248800 $D=103
M622 1392 WL_110 1614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=251710 $D=103
M623 1616 WL_111 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=252200 $D=103
M624 1392 WL_112 1618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=255110 $D=103
M625 1620 WL_113 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=255600 $D=103
M626 1392 WL_114 1622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=258510 $D=103
M627 1624 WL_115 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=259000 $D=103
M628 1392 WL_116 1626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=261910 $D=103
M629 1628 WL_117 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=262400 $D=103
M630 1392 WL_118 1630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=265310 $D=103
M631 1632 WL_119 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=265800 $D=103
M632 1392 WL_120 1634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=268710 $D=103
M633 1636 WL_121 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=269200 $D=103
M634 1392 WL_122 1638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=272110 $D=103
M635 1640 WL_123 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=272600 $D=103
M636 1392 WL_124 1642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=275510 $D=103
M637 1644 WL_125 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=276000 $D=103
M638 1392 WL_126 1646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=278910 $D=103
M639 1648 WL_127 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=279400 $D=103
M640 1392 WL_128 1650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=282310 $D=103
M641 1652 WL_129 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=282800 $D=103
M642 1392 WL_130 1654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=285710 $D=103
M643 1656 WL_131 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=286200 $D=103
M644 1392 WL_132 1658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=289110 $D=103
M645 1660 WL_133 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=289600 $D=103
M646 1392 WL_134 1662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=292510 $D=103
M647 1664 WL_135 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=293000 $D=103
M648 1392 WL_136 1666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=295910 $D=103
M649 1668 WL_137 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=296400 $D=103
M650 1392 WL_138 1670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=299310 $D=103
M651 1672 WL_139 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=299800 $D=103
M652 1392 WL_140 1674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=302710 $D=103
M653 1676 WL_141 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=303200 $D=103
M654 1392 WL_142 1678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=306110 $D=103
M655 1680 WL_143 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=306600 $D=103
M656 1392 WL_144 1682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=309510 $D=103
M657 1684 WL_145 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=310000 $D=103
M658 1392 WL_146 1686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=312910 $D=103
M659 1688 WL_147 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=313400 $D=103
M660 1392 WL_148 1690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=316310 $D=103
M661 1692 WL_149 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=316800 $D=103
M662 1392 WL_150 1694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=319710 $D=103
M663 1696 WL_151 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=320200 $D=103
M664 1392 WL_152 1698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=323110 $D=103
M665 1700 WL_153 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=323600 $D=103
M666 1392 WL_154 1702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=326510 $D=103
M667 1704 WL_155 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=327000 $D=103
M668 1392 WL_156 1706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=329910 $D=103
M669 1708 WL_157 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=330400 $D=103
M670 1392 WL_158 1710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=333310 $D=103
M671 1712 WL_159 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=333800 $D=103
M672 1392 WL_160 1714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=336710 $D=103
M673 1716 WL_161 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=337200 $D=103
M674 1392 WL_162 1718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=340110 $D=103
M675 1720 WL_163 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=340600 $D=103
M676 1392 WL_164 1722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=343510 $D=103
M677 1724 WL_165 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=344000 $D=103
M678 1392 WL_166 1726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=346910 $D=103
M679 1728 WL_167 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=347400 $D=103
M680 1392 WL_168 1730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=350310 $D=103
M681 1732 WL_169 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=350800 $D=103
M682 1392 WL_170 1734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=353710 $D=103
M683 1736 WL_171 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=354200 $D=103
M684 1392 WL_172 1738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=357110 $D=103
M685 1740 WL_173 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=357600 $D=103
M686 1392 WL_174 1742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=360510 $D=103
M687 1744 WL_175 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=361000 $D=103
M688 1392 WL_176 1746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=363910 $D=103
M689 1748 WL_177 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=364400 $D=103
M690 1392 WL_178 1750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=367310 $D=103
M691 1752 WL_179 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=367800 $D=103
M692 1392 WL_180 1754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=370710 $D=103
M693 1756 WL_181 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=371200 $D=103
M694 1392 WL_182 1758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=374110 $D=103
M695 1760 WL_183 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=374600 $D=103
M696 1392 WL_184 1762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=377510 $D=103
M697 1764 WL_185 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=378000 $D=103
M698 1392 WL_186 1766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=380910 $D=103
M699 1768 WL_187 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=381400 $D=103
M700 1392 WL_188 1770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=384310 $D=103
M701 1772 WL_189 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=384800 $D=103
M702 1392 WL_190 1774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=387710 $D=103
M703 1776 WL_191 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=388200 $D=103
M704 1392 WL_192 1778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=391110 $D=103
M705 1780 WL_193 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=391600 $D=103
M706 1392 WL_194 1782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=394510 $D=103
M707 1784 WL_195 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=395000 $D=103
M708 1392 WL_196 1786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=397910 $D=103
M709 1788 WL_197 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=398400 $D=103
M710 1392 WL_198 1790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=401310 $D=103
M711 1792 WL_199 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=401800 $D=103
M712 1392 WL_200 1794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=404710 $D=103
M713 1796 WL_201 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=405200 $D=103
M714 1392 WL_202 1798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=408110 $D=103
M715 1800 WL_203 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=408600 $D=103
M716 1392 WL_204 1802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=411510 $D=103
M717 1804 WL_205 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=412000 $D=103
M718 1392 WL_206 1806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=414910 $D=103
M719 1808 WL_207 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=415400 $D=103
M720 1392 WL_208 1810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=418310 $D=103
M721 1812 WL_209 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=418800 $D=103
M722 1392 WL_210 1814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=421710 $D=103
M723 1816 WL_211 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=422200 $D=103
M724 1392 WL_212 1818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=425110 $D=103
M725 1820 WL_213 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=425600 $D=103
M726 1392 WL_214 1822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=428510 $D=103
M727 1824 WL_215 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=429000 $D=103
M728 1392 WL_216 1826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=431910 $D=103
M729 1828 WL_217 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=432400 $D=103
M730 1392 WL_218 1830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=435310 $D=103
M731 1832 WL_219 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=435800 $D=103
M732 1392 WL_220 1834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=438710 $D=103
M733 1836 WL_221 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=439200 $D=103
M734 1392 WL_222 1838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=442110 $D=103
M735 1840 WL_223 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=442600 $D=103
M736 1392 WL_224 1842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=445510 $D=103
M737 1844 WL_225 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=446000 $D=103
M738 1392 WL_226 1846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=448910 $D=103
M739 1848 WL_227 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=449400 $D=103
M740 1392 WL_228 1850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=452310 $D=103
M741 1852 WL_229 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=452800 $D=103
M742 1392 WL_230 1854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=455710 $D=103
M743 1856 WL_231 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=456200 $D=103
M744 1392 WL_232 1858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=459110 $D=103
M745 1860 WL_233 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=459600 $D=103
M746 1392 WL_234 1862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=462510 $D=103
M747 1864 WL_235 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=463000 $D=103
M748 1392 WL_236 1866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=465910 $D=103
M749 1868 WL_237 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=466400 $D=103
M750 1392 WL_238 1870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=469310 $D=103
M751 1872 WL_239 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=469800 $D=103
M752 1392 WL_240 1874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=472710 $D=103
M753 1876 WL_241 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=473200 $D=103
M754 1392 WL_242 1878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=476110 $D=103
M755 1880 WL_243 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=476600 $D=103
M756 1392 WL_244 1882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=479510 $D=103
M757 1884 WL_245 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=480000 $D=103
M758 1392 WL_246 1886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=482910 $D=103
M759 1888 WL_247 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=483400 $D=103
M760 1392 WL_248 1890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=486310 $D=103
M761 1892 WL_249 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=486800 $D=103
M762 1392 WL_250 1894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=489710 $D=103
M763 1896 WL_251 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=490200 $D=103
M764 1392 WL_252 1898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=493110 $D=103
M765 1900 WL_253 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=493600 $D=103
M766 1392 WL_254 1902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=496510 $D=103
M767 1904 WL_255 1392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38150 $Y=497000 $D=103
M768 1906 WL_0 1907 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=64710 $D=103
M769 1909 WL_1 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=65200 $D=103
M770 1906 WL_2 1911 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=68110 $D=103
M771 1913 WL_3 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=68600 $D=103
M772 1906 WL_4 1915 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=71510 $D=103
M773 1917 WL_5 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=72000 $D=103
M774 1906 WL_6 1919 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=74910 $D=103
M775 1921 WL_7 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=75400 $D=103
M776 1906 WL_8 1923 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=78310 $D=103
M777 1925 WL_9 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=78800 $D=103
M778 1906 WL_10 1927 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=81710 $D=103
M779 1929 WL_11 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=82200 $D=103
M780 1906 WL_12 1931 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=85110 $D=103
M781 1933 WL_13 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=85600 $D=103
M782 1906 WL_14 1935 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=88510 $D=103
M783 1937 WL_15 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=89000 $D=103
M784 1906 WL_16 1939 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=91910 $D=103
M785 1941 WL_17 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=92400 $D=103
M786 1906 WL_18 1943 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=95310 $D=103
M787 1945 WL_19 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=95800 $D=103
M788 1906 WL_20 1947 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=98710 $D=103
M789 1949 WL_21 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=99200 $D=103
M790 1906 WL_22 1951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=102110 $D=103
M791 1953 WL_23 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=102600 $D=103
M792 1906 WL_24 1955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=105510 $D=103
M793 1957 WL_25 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=106000 $D=103
M794 1906 WL_26 1959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=108910 $D=103
M795 1961 WL_27 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=109400 $D=103
M796 1906 WL_28 1963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=112310 $D=103
M797 1965 WL_29 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=112800 $D=103
M798 1906 WL_30 1967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=115710 $D=103
M799 1969 WL_31 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=116200 $D=103
M800 1906 WL_32 1971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=119110 $D=103
M801 1973 WL_33 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=119600 $D=103
M802 1906 WL_34 1975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=122510 $D=103
M803 1977 WL_35 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=123000 $D=103
M804 1906 WL_36 1979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=125910 $D=103
M805 1981 WL_37 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=126400 $D=103
M806 1906 WL_38 1983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=129310 $D=103
M807 1985 WL_39 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=129800 $D=103
M808 1906 WL_40 1987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=132710 $D=103
M809 1989 WL_41 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=133200 $D=103
M810 1906 WL_42 1991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=136110 $D=103
M811 1993 WL_43 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=136600 $D=103
M812 1906 WL_44 1995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=139510 $D=103
M813 1997 WL_45 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=140000 $D=103
M814 1906 WL_46 1999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=142910 $D=103
M815 2001 WL_47 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=143400 $D=103
M816 1906 WL_48 2003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=146310 $D=103
M817 2005 WL_49 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=146800 $D=103
M818 1906 WL_50 2007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=149710 $D=103
M819 2009 WL_51 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=150200 $D=103
M820 1906 WL_52 2011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=153110 $D=103
M821 2013 WL_53 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=153600 $D=103
M822 1906 WL_54 2015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=156510 $D=103
M823 2017 WL_55 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=157000 $D=103
M824 1906 WL_56 2019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=159910 $D=103
M825 2021 WL_57 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=160400 $D=103
M826 1906 WL_58 2023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=163310 $D=103
M827 2025 WL_59 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=163800 $D=103
M828 1906 WL_60 2027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=166710 $D=103
M829 2029 WL_61 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=167200 $D=103
M830 1906 WL_62 2031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=170110 $D=103
M831 2033 WL_63 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=170600 $D=103
M832 1906 WL_64 2035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=173510 $D=103
M833 2037 WL_65 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=174000 $D=103
M834 1906 WL_66 2039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=176910 $D=103
M835 2041 WL_67 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=177400 $D=103
M836 1906 WL_68 2043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=180310 $D=103
M837 2045 WL_69 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=180800 $D=103
M838 1906 WL_70 2047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=183710 $D=103
M839 2049 WL_71 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=184200 $D=103
M840 1906 WL_72 2051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=187110 $D=103
M841 2053 WL_73 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=187600 $D=103
M842 1906 WL_74 2055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=190510 $D=103
M843 2057 WL_75 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=191000 $D=103
M844 1906 WL_76 2059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=193910 $D=103
M845 2061 WL_77 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=194400 $D=103
M846 1906 WL_78 2063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=197310 $D=103
M847 2065 WL_79 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=197800 $D=103
M848 1906 WL_80 2067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=200710 $D=103
M849 2069 WL_81 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=201200 $D=103
M850 1906 WL_82 2071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=204110 $D=103
M851 2073 WL_83 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=204600 $D=103
M852 1906 WL_84 2075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=207510 $D=103
M853 2077 WL_85 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=208000 $D=103
M854 1906 WL_86 2079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=210910 $D=103
M855 2081 WL_87 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=211400 $D=103
M856 1906 WL_88 2083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=214310 $D=103
M857 2085 WL_89 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=214800 $D=103
M858 1906 WL_90 2087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=217710 $D=103
M859 2089 WL_91 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=218200 $D=103
M860 1906 WL_92 2091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=221110 $D=103
M861 2093 WL_93 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=221600 $D=103
M862 1906 WL_94 2095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=224510 $D=103
M863 2097 WL_95 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=225000 $D=103
M864 1906 WL_96 2099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=227910 $D=103
M865 2101 WL_97 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=228400 $D=103
M866 1906 WL_98 2103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=231310 $D=103
M867 2105 WL_99 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=231800 $D=103
M868 1906 WL_100 2107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=234710 $D=103
M869 2109 WL_101 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=235200 $D=103
M870 1906 WL_102 2111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=238110 $D=103
M871 2113 WL_103 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=238600 $D=103
M872 1906 WL_104 2115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=241510 $D=103
M873 2117 WL_105 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=242000 $D=103
M874 1906 WL_106 2119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=244910 $D=103
M875 2121 WL_107 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=245400 $D=103
M876 1906 WL_108 2123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=248310 $D=103
M877 2125 WL_109 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=248800 $D=103
M878 1906 WL_110 2127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=251710 $D=103
M879 2129 WL_111 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=252200 $D=103
M880 1906 WL_112 2131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=255110 $D=103
M881 2133 WL_113 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=255600 $D=103
M882 1906 WL_114 2135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=258510 $D=103
M883 2137 WL_115 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=259000 $D=103
M884 1906 WL_116 2139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=261910 $D=103
M885 2141 WL_117 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=262400 $D=103
M886 1906 WL_118 2143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=265310 $D=103
M887 2145 WL_119 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=265800 $D=103
M888 1906 WL_120 2147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=268710 $D=103
M889 2149 WL_121 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=269200 $D=103
M890 1906 WL_122 2151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=272110 $D=103
M891 2153 WL_123 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=272600 $D=103
M892 1906 WL_124 2155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=275510 $D=103
M893 2157 WL_125 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=276000 $D=103
M894 1906 WL_126 2159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=278910 $D=103
M895 2161 WL_127 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=279400 $D=103
M896 1906 WL_128 2163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=282310 $D=103
M897 2165 WL_129 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=282800 $D=103
M898 1906 WL_130 2167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=285710 $D=103
M899 2169 WL_131 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=286200 $D=103
M900 1906 WL_132 2171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=289110 $D=103
M901 2173 WL_133 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=289600 $D=103
M902 1906 WL_134 2175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=292510 $D=103
M903 2177 WL_135 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=293000 $D=103
M904 1906 WL_136 2179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=295910 $D=103
M905 2181 WL_137 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=296400 $D=103
M906 1906 WL_138 2183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=299310 $D=103
M907 2185 WL_139 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=299800 $D=103
M908 1906 WL_140 2187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=302710 $D=103
M909 2189 WL_141 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=303200 $D=103
M910 1906 WL_142 2191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=306110 $D=103
M911 2193 WL_143 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=306600 $D=103
M912 1906 WL_144 2195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=309510 $D=103
M913 2197 WL_145 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=310000 $D=103
M914 1906 WL_146 2199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=312910 $D=103
M915 2201 WL_147 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=313400 $D=103
M916 1906 WL_148 2203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=316310 $D=103
M917 2205 WL_149 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=316800 $D=103
M918 1906 WL_150 2207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=319710 $D=103
M919 2209 WL_151 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=320200 $D=103
M920 1906 WL_152 2211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=323110 $D=103
M921 2213 WL_153 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=323600 $D=103
M922 1906 WL_154 2215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=326510 $D=103
M923 2217 WL_155 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=327000 $D=103
M924 1906 WL_156 2219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=329910 $D=103
M925 2221 WL_157 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=330400 $D=103
M926 1906 WL_158 2223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=333310 $D=103
M927 2225 WL_159 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=333800 $D=103
M928 1906 WL_160 2227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=336710 $D=103
M929 2229 WL_161 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=337200 $D=103
M930 1906 WL_162 2231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=340110 $D=103
M931 2233 WL_163 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=340600 $D=103
M932 1906 WL_164 2235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=343510 $D=103
M933 2237 WL_165 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=344000 $D=103
M934 1906 WL_166 2239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=346910 $D=103
M935 2241 WL_167 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=347400 $D=103
M936 1906 WL_168 2243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=350310 $D=103
M937 2245 WL_169 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=350800 $D=103
M938 1906 WL_170 2247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=353710 $D=103
M939 2249 WL_171 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=354200 $D=103
M940 1906 WL_172 2251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=357110 $D=103
M941 2253 WL_173 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=357600 $D=103
M942 1906 WL_174 2255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=360510 $D=103
M943 2257 WL_175 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=361000 $D=103
M944 1906 WL_176 2259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=363910 $D=103
M945 2261 WL_177 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=364400 $D=103
M946 1906 WL_178 2263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=367310 $D=103
M947 2265 WL_179 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=367800 $D=103
M948 1906 WL_180 2267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=370710 $D=103
M949 2269 WL_181 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=371200 $D=103
M950 1906 WL_182 2271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=374110 $D=103
M951 2273 WL_183 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=374600 $D=103
M952 1906 WL_184 2275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=377510 $D=103
M953 2277 WL_185 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=378000 $D=103
M954 1906 WL_186 2279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=380910 $D=103
M955 2281 WL_187 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=381400 $D=103
M956 1906 WL_188 2283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=384310 $D=103
M957 2285 WL_189 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=384800 $D=103
M958 1906 WL_190 2287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=387710 $D=103
M959 2289 WL_191 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=388200 $D=103
M960 1906 WL_192 2291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=391110 $D=103
M961 2293 WL_193 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=391600 $D=103
M962 1906 WL_194 2295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=394510 $D=103
M963 2297 WL_195 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=395000 $D=103
M964 1906 WL_196 2299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=397910 $D=103
M965 2301 WL_197 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=398400 $D=103
M966 1906 WL_198 2303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=401310 $D=103
M967 2305 WL_199 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=401800 $D=103
M968 1906 WL_200 2307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=404710 $D=103
M969 2309 WL_201 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=405200 $D=103
M970 1906 WL_202 2311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=408110 $D=103
M971 2313 WL_203 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=408600 $D=103
M972 1906 WL_204 2315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=411510 $D=103
M973 2317 WL_205 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=412000 $D=103
M974 1906 WL_206 2319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=414910 $D=103
M975 2321 WL_207 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=415400 $D=103
M976 1906 WL_208 2323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=418310 $D=103
M977 2325 WL_209 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=418800 $D=103
M978 1906 WL_210 2327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=421710 $D=103
M979 2329 WL_211 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=422200 $D=103
M980 1906 WL_212 2331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=425110 $D=103
M981 2333 WL_213 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=425600 $D=103
M982 1906 WL_214 2335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=428510 $D=103
M983 2337 WL_215 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=429000 $D=103
M984 1906 WL_216 2339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=431910 $D=103
M985 2341 WL_217 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=432400 $D=103
M986 1906 WL_218 2343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=435310 $D=103
M987 2345 WL_219 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=435800 $D=103
M988 1906 WL_220 2347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=438710 $D=103
M989 2349 WL_221 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=439200 $D=103
M990 1906 WL_222 2351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=442110 $D=103
M991 2353 WL_223 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=442600 $D=103
M992 1906 WL_224 2355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=445510 $D=103
M993 2357 WL_225 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=446000 $D=103
M994 1906 WL_226 2359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=448910 $D=103
M995 2361 WL_227 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=449400 $D=103
M996 1906 WL_228 2363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=452310 $D=103
M997 2365 WL_229 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=452800 $D=103
M998 1906 WL_230 2367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=455710 $D=103
M999 2369 WL_231 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=456200 $D=103
M1000 1906 WL_232 2371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=459110 $D=103
M1001 2373 WL_233 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=459600 $D=103
M1002 1906 WL_234 2375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=462510 $D=103
M1003 2377 WL_235 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=463000 $D=103
M1004 1906 WL_236 2379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=465910 $D=103
M1005 2381 WL_237 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=466400 $D=103
M1006 1906 WL_238 2383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=469310 $D=103
M1007 2385 WL_239 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=469800 $D=103
M1008 1906 WL_240 2387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=472710 $D=103
M1009 2389 WL_241 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=473200 $D=103
M1010 1906 WL_242 2391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=476110 $D=103
M1011 2393 WL_243 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=476600 $D=103
M1012 1906 WL_244 2395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=479510 $D=103
M1013 2397 WL_245 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=480000 $D=103
M1014 1906 WL_246 2399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=482910 $D=103
M1015 2401 WL_247 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=483400 $D=103
M1016 1906 WL_248 2403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=486310 $D=103
M1017 2405 WL_249 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=486800 $D=103
M1018 1906 WL_250 2407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=489710 $D=103
M1019 2409 WL_251 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=490200 $D=103
M1020 1906 WL_252 2411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=493110 $D=103
M1021 2413 WL_253 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=493600 $D=103
M1022 1906 WL_254 2415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=496510 $D=103
M1023 2417 WL_255 1906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39690 $Y=497000 $D=103
M1024 1905 WL_0 1908 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=64710 $D=103
M1025 1910 WL_1 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=65200 $D=103
M1026 1905 WL_2 1912 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=68110 $D=103
M1027 1914 WL_3 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=68600 $D=103
M1028 1905 WL_4 1916 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=71510 $D=103
M1029 1918 WL_5 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=72000 $D=103
M1030 1905 WL_6 1920 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=74910 $D=103
M1031 1922 WL_7 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=75400 $D=103
M1032 1905 WL_8 1924 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=78310 $D=103
M1033 1926 WL_9 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=78800 $D=103
M1034 1905 WL_10 1928 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=81710 $D=103
M1035 1930 WL_11 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=82200 $D=103
M1036 1905 WL_12 1932 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=85110 $D=103
M1037 1934 WL_13 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=85600 $D=103
M1038 1905 WL_14 1936 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=88510 $D=103
M1039 1938 WL_15 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=89000 $D=103
M1040 1905 WL_16 1940 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=91910 $D=103
M1041 1942 WL_17 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=92400 $D=103
M1042 1905 WL_18 1944 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=95310 $D=103
M1043 1946 WL_19 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=95800 $D=103
M1044 1905 WL_20 1948 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=98710 $D=103
M1045 1950 WL_21 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=99200 $D=103
M1046 1905 WL_22 1952 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=102110 $D=103
M1047 1954 WL_23 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=102600 $D=103
M1048 1905 WL_24 1956 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=105510 $D=103
M1049 1958 WL_25 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=106000 $D=103
M1050 1905 WL_26 1960 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=108910 $D=103
M1051 1962 WL_27 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=109400 $D=103
M1052 1905 WL_28 1964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=112310 $D=103
M1053 1966 WL_29 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=112800 $D=103
M1054 1905 WL_30 1968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=115710 $D=103
M1055 1970 WL_31 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=116200 $D=103
M1056 1905 WL_32 1972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=119110 $D=103
M1057 1974 WL_33 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=119600 $D=103
M1058 1905 WL_34 1976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=122510 $D=103
M1059 1978 WL_35 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=123000 $D=103
M1060 1905 WL_36 1980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=125910 $D=103
M1061 1982 WL_37 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=126400 $D=103
M1062 1905 WL_38 1984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=129310 $D=103
M1063 1986 WL_39 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=129800 $D=103
M1064 1905 WL_40 1988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=132710 $D=103
M1065 1990 WL_41 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=133200 $D=103
M1066 1905 WL_42 1992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=136110 $D=103
M1067 1994 WL_43 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=136600 $D=103
M1068 1905 WL_44 1996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=139510 $D=103
M1069 1998 WL_45 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=140000 $D=103
M1070 1905 WL_46 2000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=142910 $D=103
M1071 2002 WL_47 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=143400 $D=103
M1072 1905 WL_48 2004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=146310 $D=103
M1073 2006 WL_49 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=146800 $D=103
M1074 1905 WL_50 2008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=149710 $D=103
M1075 2010 WL_51 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=150200 $D=103
M1076 1905 WL_52 2012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=153110 $D=103
M1077 2014 WL_53 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=153600 $D=103
M1078 1905 WL_54 2016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=156510 $D=103
M1079 2018 WL_55 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=157000 $D=103
M1080 1905 WL_56 2020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=159910 $D=103
M1081 2022 WL_57 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=160400 $D=103
M1082 1905 WL_58 2024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=163310 $D=103
M1083 2026 WL_59 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=163800 $D=103
M1084 1905 WL_60 2028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=166710 $D=103
M1085 2030 WL_61 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=167200 $D=103
M1086 1905 WL_62 2032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=170110 $D=103
M1087 2034 WL_63 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=170600 $D=103
M1088 1905 WL_64 2036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=173510 $D=103
M1089 2038 WL_65 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=174000 $D=103
M1090 1905 WL_66 2040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=176910 $D=103
M1091 2042 WL_67 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=177400 $D=103
M1092 1905 WL_68 2044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=180310 $D=103
M1093 2046 WL_69 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=180800 $D=103
M1094 1905 WL_70 2048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=183710 $D=103
M1095 2050 WL_71 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=184200 $D=103
M1096 1905 WL_72 2052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=187110 $D=103
M1097 2054 WL_73 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=187600 $D=103
M1098 1905 WL_74 2056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=190510 $D=103
M1099 2058 WL_75 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=191000 $D=103
M1100 1905 WL_76 2060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=193910 $D=103
M1101 2062 WL_77 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=194400 $D=103
M1102 1905 WL_78 2064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=197310 $D=103
M1103 2066 WL_79 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=197800 $D=103
M1104 1905 WL_80 2068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=200710 $D=103
M1105 2070 WL_81 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=201200 $D=103
M1106 1905 WL_82 2072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=204110 $D=103
M1107 2074 WL_83 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=204600 $D=103
M1108 1905 WL_84 2076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=207510 $D=103
M1109 2078 WL_85 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=208000 $D=103
M1110 1905 WL_86 2080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=210910 $D=103
M1111 2082 WL_87 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=211400 $D=103
M1112 1905 WL_88 2084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=214310 $D=103
M1113 2086 WL_89 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=214800 $D=103
M1114 1905 WL_90 2088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=217710 $D=103
M1115 2090 WL_91 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=218200 $D=103
M1116 1905 WL_92 2092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=221110 $D=103
M1117 2094 WL_93 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=221600 $D=103
M1118 1905 WL_94 2096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=224510 $D=103
M1119 2098 WL_95 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=225000 $D=103
M1120 1905 WL_96 2100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=227910 $D=103
M1121 2102 WL_97 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=228400 $D=103
M1122 1905 WL_98 2104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=231310 $D=103
M1123 2106 WL_99 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=231800 $D=103
M1124 1905 WL_100 2108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=234710 $D=103
M1125 2110 WL_101 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=235200 $D=103
M1126 1905 WL_102 2112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=238110 $D=103
M1127 2114 WL_103 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=238600 $D=103
M1128 1905 WL_104 2116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=241510 $D=103
M1129 2118 WL_105 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=242000 $D=103
M1130 1905 WL_106 2120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=244910 $D=103
M1131 2122 WL_107 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=245400 $D=103
M1132 1905 WL_108 2124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=248310 $D=103
M1133 2126 WL_109 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=248800 $D=103
M1134 1905 WL_110 2128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=251710 $D=103
M1135 2130 WL_111 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=252200 $D=103
M1136 1905 WL_112 2132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=255110 $D=103
M1137 2134 WL_113 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=255600 $D=103
M1138 1905 WL_114 2136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=258510 $D=103
M1139 2138 WL_115 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=259000 $D=103
M1140 1905 WL_116 2140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=261910 $D=103
M1141 2142 WL_117 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=262400 $D=103
M1142 1905 WL_118 2144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=265310 $D=103
M1143 2146 WL_119 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=265800 $D=103
M1144 1905 WL_120 2148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=268710 $D=103
M1145 2150 WL_121 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=269200 $D=103
M1146 1905 WL_122 2152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=272110 $D=103
M1147 2154 WL_123 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=272600 $D=103
M1148 1905 WL_124 2156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=275510 $D=103
M1149 2158 WL_125 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=276000 $D=103
M1150 1905 WL_126 2160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=278910 $D=103
M1151 2162 WL_127 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=279400 $D=103
M1152 1905 WL_128 2164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=282310 $D=103
M1153 2166 WL_129 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=282800 $D=103
M1154 1905 WL_130 2168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=285710 $D=103
M1155 2170 WL_131 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=286200 $D=103
M1156 1905 WL_132 2172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=289110 $D=103
M1157 2174 WL_133 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=289600 $D=103
M1158 1905 WL_134 2176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=292510 $D=103
M1159 2178 WL_135 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=293000 $D=103
M1160 1905 WL_136 2180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=295910 $D=103
M1161 2182 WL_137 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=296400 $D=103
M1162 1905 WL_138 2184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=299310 $D=103
M1163 2186 WL_139 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=299800 $D=103
M1164 1905 WL_140 2188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=302710 $D=103
M1165 2190 WL_141 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=303200 $D=103
M1166 1905 WL_142 2192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=306110 $D=103
M1167 2194 WL_143 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=306600 $D=103
M1168 1905 WL_144 2196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=309510 $D=103
M1169 2198 WL_145 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=310000 $D=103
M1170 1905 WL_146 2200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=312910 $D=103
M1171 2202 WL_147 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=313400 $D=103
M1172 1905 WL_148 2204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=316310 $D=103
M1173 2206 WL_149 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=316800 $D=103
M1174 1905 WL_150 2208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=319710 $D=103
M1175 2210 WL_151 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=320200 $D=103
M1176 1905 WL_152 2212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=323110 $D=103
M1177 2214 WL_153 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=323600 $D=103
M1178 1905 WL_154 2216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=326510 $D=103
M1179 2218 WL_155 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=327000 $D=103
M1180 1905 WL_156 2220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=329910 $D=103
M1181 2222 WL_157 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=330400 $D=103
M1182 1905 WL_158 2224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=333310 $D=103
M1183 2226 WL_159 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=333800 $D=103
M1184 1905 WL_160 2228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=336710 $D=103
M1185 2230 WL_161 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=337200 $D=103
M1186 1905 WL_162 2232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=340110 $D=103
M1187 2234 WL_163 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=340600 $D=103
M1188 1905 WL_164 2236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=343510 $D=103
M1189 2238 WL_165 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=344000 $D=103
M1190 1905 WL_166 2240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=346910 $D=103
M1191 2242 WL_167 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=347400 $D=103
M1192 1905 WL_168 2244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=350310 $D=103
M1193 2246 WL_169 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=350800 $D=103
M1194 1905 WL_170 2248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=353710 $D=103
M1195 2250 WL_171 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=354200 $D=103
M1196 1905 WL_172 2252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=357110 $D=103
M1197 2254 WL_173 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=357600 $D=103
M1198 1905 WL_174 2256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=360510 $D=103
M1199 2258 WL_175 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=361000 $D=103
M1200 1905 WL_176 2260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=363910 $D=103
M1201 2262 WL_177 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=364400 $D=103
M1202 1905 WL_178 2264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=367310 $D=103
M1203 2266 WL_179 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=367800 $D=103
M1204 1905 WL_180 2268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=370710 $D=103
M1205 2270 WL_181 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=371200 $D=103
M1206 1905 WL_182 2272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=374110 $D=103
M1207 2274 WL_183 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=374600 $D=103
M1208 1905 WL_184 2276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=377510 $D=103
M1209 2278 WL_185 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=378000 $D=103
M1210 1905 WL_186 2280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=380910 $D=103
M1211 2282 WL_187 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=381400 $D=103
M1212 1905 WL_188 2284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=384310 $D=103
M1213 2286 WL_189 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=384800 $D=103
M1214 1905 WL_190 2288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=387710 $D=103
M1215 2290 WL_191 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=388200 $D=103
M1216 1905 WL_192 2292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=391110 $D=103
M1217 2294 WL_193 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=391600 $D=103
M1218 1905 WL_194 2296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=394510 $D=103
M1219 2298 WL_195 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=395000 $D=103
M1220 1905 WL_196 2300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=397910 $D=103
M1221 2302 WL_197 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=398400 $D=103
M1222 1905 WL_198 2304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=401310 $D=103
M1223 2306 WL_199 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=401800 $D=103
M1224 1905 WL_200 2308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=404710 $D=103
M1225 2310 WL_201 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=405200 $D=103
M1226 1905 WL_202 2312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=408110 $D=103
M1227 2314 WL_203 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=408600 $D=103
M1228 1905 WL_204 2316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=411510 $D=103
M1229 2318 WL_205 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=412000 $D=103
M1230 1905 WL_206 2320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=414910 $D=103
M1231 2322 WL_207 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=415400 $D=103
M1232 1905 WL_208 2324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=418310 $D=103
M1233 2326 WL_209 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=418800 $D=103
M1234 1905 WL_210 2328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=421710 $D=103
M1235 2330 WL_211 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=422200 $D=103
M1236 1905 WL_212 2332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=425110 $D=103
M1237 2334 WL_213 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=425600 $D=103
M1238 1905 WL_214 2336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=428510 $D=103
M1239 2338 WL_215 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=429000 $D=103
M1240 1905 WL_216 2340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=431910 $D=103
M1241 2342 WL_217 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=432400 $D=103
M1242 1905 WL_218 2344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=435310 $D=103
M1243 2346 WL_219 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=435800 $D=103
M1244 1905 WL_220 2348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=438710 $D=103
M1245 2350 WL_221 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=439200 $D=103
M1246 1905 WL_222 2352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=442110 $D=103
M1247 2354 WL_223 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=442600 $D=103
M1248 1905 WL_224 2356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=445510 $D=103
M1249 2358 WL_225 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=446000 $D=103
M1250 1905 WL_226 2360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=448910 $D=103
M1251 2362 WL_227 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=449400 $D=103
M1252 1905 WL_228 2364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=452310 $D=103
M1253 2366 WL_229 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=452800 $D=103
M1254 1905 WL_230 2368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=455710 $D=103
M1255 2370 WL_231 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=456200 $D=103
M1256 1905 WL_232 2372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=459110 $D=103
M1257 2374 WL_233 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=459600 $D=103
M1258 1905 WL_234 2376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=462510 $D=103
M1259 2378 WL_235 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=463000 $D=103
M1260 1905 WL_236 2380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=465910 $D=103
M1261 2382 WL_237 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=466400 $D=103
M1262 1905 WL_238 2384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=469310 $D=103
M1263 2386 WL_239 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=469800 $D=103
M1264 1905 WL_240 2388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=472710 $D=103
M1265 2390 WL_241 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=473200 $D=103
M1266 1905 WL_242 2392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=476110 $D=103
M1267 2394 WL_243 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=476600 $D=103
M1268 1905 WL_244 2396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=479510 $D=103
M1269 2398 WL_245 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=480000 $D=103
M1270 1905 WL_246 2400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=482910 $D=103
M1271 2402 WL_247 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=483400 $D=103
M1272 1905 WL_248 2404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=486310 $D=103
M1273 2406 WL_249 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=486800 $D=103
M1274 1905 WL_250 2408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=489710 $D=103
M1275 2410 WL_251 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=490200 $D=103
M1276 1905 WL_252 2412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=493110 $D=103
M1277 2414 WL_253 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=493600 $D=103
M1278 1905 WL_254 2416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=496510 $D=103
M1279 2418 WL_255 1905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58550 $Y=497000 $D=103
M1280 2419 WL_0 2421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=64710 $D=103
M1281 2423 WL_1 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=65200 $D=103
M1282 2419 WL_2 2425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=68110 $D=103
M1283 2427 WL_3 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=68600 $D=103
M1284 2419 WL_4 2429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=71510 $D=103
M1285 2431 WL_5 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=72000 $D=103
M1286 2419 WL_6 2433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=74910 $D=103
M1287 2435 WL_7 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=75400 $D=103
M1288 2419 WL_8 2437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=78310 $D=103
M1289 2439 WL_9 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=78800 $D=103
M1290 2419 WL_10 2441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=81710 $D=103
M1291 2443 WL_11 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=82200 $D=103
M1292 2419 WL_12 2445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=85110 $D=103
M1293 2447 WL_13 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=85600 $D=103
M1294 2419 WL_14 2449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=88510 $D=103
M1295 2451 WL_15 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=89000 $D=103
M1296 2419 WL_16 2453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=91910 $D=103
M1297 2455 WL_17 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=92400 $D=103
M1298 2419 WL_18 2457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=95310 $D=103
M1299 2459 WL_19 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=95800 $D=103
M1300 2419 WL_20 2461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=98710 $D=103
M1301 2463 WL_21 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=99200 $D=103
M1302 2419 WL_22 2465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=102110 $D=103
M1303 2467 WL_23 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=102600 $D=103
M1304 2419 WL_24 2469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=105510 $D=103
M1305 2471 WL_25 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=106000 $D=103
M1306 2419 WL_26 2473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=108910 $D=103
M1307 2475 WL_27 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=109400 $D=103
M1308 2419 WL_28 2477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=112310 $D=103
M1309 2479 WL_29 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=112800 $D=103
M1310 2419 WL_30 2481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=115710 $D=103
M1311 2483 WL_31 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=116200 $D=103
M1312 2419 WL_32 2485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=119110 $D=103
M1313 2487 WL_33 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=119600 $D=103
M1314 2419 WL_34 2489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=122510 $D=103
M1315 2491 WL_35 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=123000 $D=103
M1316 2419 WL_36 2493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=125910 $D=103
M1317 2495 WL_37 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=126400 $D=103
M1318 2419 WL_38 2497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=129310 $D=103
M1319 2499 WL_39 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=129800 $D=103
M1320 2419 WL_40 2501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=132710 $D=103
M1321 2503 WL_41 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=133200 $D=103
M1322 2419 WL_42 2505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=136110 $D=103
M1323 2507 WL_43 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=136600 $D=103
M1324 2419 WL_44 2509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=139510 $D=103
M1325 2511 WL_45 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=140000 $D=103
M1326 2419 WL_46 2513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=142910 $D=103
M1327 2515 WL_47 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=143400 $D=103
M1328 2419 WL_48 2517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=146310 $D=103
M1329 2519 WL_49 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=146800 $D=103
M1330 2419 WL_50 2521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=149710 $D=103
M1331 2523 WL_51 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=150200 $D=103
M1332 2419 WL_52 2525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=153110 $D=103
M1333 2527 WL_53 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=153600 $D=103
M1334 2419 WL_54 2529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=156510 $D=103
M1335 2531 WL_55 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=157000 $D=103
M1336 2419 WL_56 2533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=159910 $D=103
M1337 2535 WL_57 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=160400 $D=103
M1338 2419 WL_58 2537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=163310 $D=103
M1339 2539 WL_59 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=163800 $D=103
M1340 2419 WL_60 2541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=166710 $D=103
M1341 2543 WL_61 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=167200 $D=103
M1342 2419 WL_62 2545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=170110 $D=103
M1343 2547 WL_63 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=170600 $D=103
M1344 2419 WL_64 2549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=173510 $D=103
M1345 2551 WL_65 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=174000 $D=103
M1346 2419 WL_66 2553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=176910 $D=103
M1347 2555 WL_67 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=177400 $D=103
M1348 2419 WL_68 2557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=180310 $D=103
M1349 2559 WL_69 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=180800 $D=103
M1350 2419 WL_70 2561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=183710 $D=103
M1351 2563 WL_71 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=184200 $D=103
M1352 2419 WL_72 2565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=187110 $D=103
M1353 2567 WL_73 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=187600 $D=103
M1354 2419 WL_74 2569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=190510 $D=103
M1355 2571 WL_75 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=191000 $D=103
M1356 2419 WL_76 2573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=193910 $D=103
M1357 2575 WL_77 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=194400 $D=103
M1358 2419 WL_78 2577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=197310 $D=103
M1359 2579 WL_79 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=197800 $D=103
M1360 2419 WL_80 2581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=200710 $D=103
M1361 2583 WL_81 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=201200 $D=103
M1362 2419 WL_82 2585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=204110 $D=103
M1363 2587 WL_83 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=204600 $D=103
M1364 2419 WL_84 2589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=207510 $D=103
M1365 2591 WL_85 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=208000 $D=103
M1366 2419 WL_86 2593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=210910 $D=103
M1367 2595 WL_87 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=211400 $D=103
M1368 2419 WL_88 2597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=214310 $D=103
M1369 2599 WL_89 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=214800 $D=103
M1370 2419 WL_90 2601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=217710 $D=103
M1371 2603 WL_91 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=218200 $D=103
M1372 2419 WL_92 2605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=221110 $D=103
M1373 2607 WL_93 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=221600 $D=103
M1374 2419 WL_94 2609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=224510 $D=103
M1375 2611 WL_95 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=225000 $D=103
M1376 2419 WL_96 2613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=227910 $D=103
M1377 2615 WL_97 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=228400 $D=103
M1378 2419 WL_98 2617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=231310 $D=103
M1379 2619 WL_99 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=231800 $D=103
M1380 2419 WL_100 2621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=234710 $D=103
M1381 2623 WL_101 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=235200 $D=103
M1382 2419 WL_102 2625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=238110 $D=103
M1383 2627 WL_103 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=238600 $D=103
M1384 2419 WL_104 2629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=241510 $D=103
M1385 2631 WL_105 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=242000 $D=103
M1386 2419 WL_106 2633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=244910 $D=103
M1387 2635 WL_107 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=245400 $D=103
M1388 2419 WL_108 2637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=248310 $D=103
M1389 2639 WL_109 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=248800 $D=103
M1390 2419 WL_110 2641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=251710 $D=103
M1391 2643 WL_111 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=252200 $D=103
M1392 2419 WL_112 2645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=255110 $D=103
M1393 2647 WL_113 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=255600 $D=103
M1394 2419 WL_114 2649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=258510 $D=103
M1395 2651 WL_115 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=259000 $D=103
M1396 2419 WL_116 2653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=261910 $D=103
M1397 2655 WL_117 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=262400 $D=103
M1398 2419 WL_118 2657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=265310 $D=103
M1399 2659 WL_119 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=265800 $D=103
M1400 2419 WL_120 2661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=268710 $D=103
M1401 2663 WL_121 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=269200 $D=103
M1402 2419 WL_122 2665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=272110 $D=103
M1403 2667 WL_123 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=272600 $D=103
M1404 2419 WL_124 2669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=275510 $D=103
M1405 2671 WL_125 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=276000 $D=103
M1406 2419 WL_126 2673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=278910 $D=103
M1407 2675 WL_127 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=279400 $D=103
M1408 2419 WL_128 2677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=282310 $D=103
M1409 2679 WL_129 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=282800 $D=103
M1410 2419 WL_130 2681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=285710 $D=103
M1411 2683 WL_131 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=286200 $D=103
M1412 2419 WL_132 2685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=289110 $D=103
M1413 2687 WL_133 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=289600 $D=103
M1414 2419 WL_134 2689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=292510 $D=103
M1415 2691 WL_135 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=293000 $D=103
M1416 2419 WL_136 2693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=295910 $D=103
M1417 2695 WL_137 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=296400 $D=103
M1418 2419 WL_138 2697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=299310 $D=103
M1419 2699 WL_139 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=299800 $D=103
M1420 2419 WL_140 2701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=302710 $D=103
M1421 2703 WL_141 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=303200 $D=103
M1422 2419 WL_142 2705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=306110 $D=103
M1423 2707 WL_143 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=306600 $D=103
M1424 2419 WL_144 2709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=309510 $D=103
M1425 2711 WL_145 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=310000 $D=103
M1426 2419 WL_146 2713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=312910 $D=103
M1427 2715 WL_147 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=313400 $D=103
M1428 2419 WL_148 2717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=316310 $D=103
M1429 2719 WL_149 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=316800 $D=103
M1430 2419 WL_150 2721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=319710 $D=103
M1431 2723 WL_151 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=320200 $D=103
M1432 2419 WL_152 2725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=323110 $D=103
M1433 2727 WL_153 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=323600 $D=103
M1434 2419 WL_154 2729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=326510 $D=103
M1435 2731 WL_155 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=327000 $D=103
M1436 2419 WL_156 2733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=329910 $D=103
M1437 2735 WL_157 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=330400 $D=103
M1438 2419 WL_158 2737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=333310 $D=103
M1439 2739 WL_159 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=333800 $D=103
M1440 2419 WL_160 2741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=336710 $D=103
M1441 2743 WL_161 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=337200 $D=103
M1442 2419 WL_162 2745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=340110 $D=103
M1443 2747 WL_163 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=340600 $D=103
M1444 2419 WL_164 2749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=343510 $D=103
M1445 2751 WL_165 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=344000 $D=103
M1446 2419 WL_166 2753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=346910 $D=103
M1447 2755 WL_167 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=347400 $D=103
M1448 2419 WL_168 2757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=350310 $D=103
M1449 2759 WL_169 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=350800 $D=103
M1450 2419 WL_170 2761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=353710 $D=103
M1451 2763 WL_171 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=354200 $D=103
M1452 2419 WL_172 2765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=357110 $D=103
M1453 2767 WL_173 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=357600 $D=103
M1454 2419 WL_174 2769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=360510 $D=103
M1455 2771 WL_175 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=361000 $D=103
M1456 2419 WL_176 2773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=363910 $D=103
M1457 2775 WL_177 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=364400 $D=103
M1458 2419 WL_178 2777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=367310 $D=103
M1459 2779 WL_179 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=367800 $D=103
M1460 2419 WL_180 2781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=370710 $D=103
M1461 2783 WL_181 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=371200 $D=103
M1462 2419 WL_182 2785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=374110 $D=103
M1463 2787 WL_183 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=374600 $D=103
M1464 2419 WL_184 2789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=377510 $D=103
M1465 2791 WL_185 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=378000 $D=103
M1466 2419 WL_186 2793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=380910 $D=103
M1467 2795 WL_187 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=381400 $D=103
M1468 2419 WL_188 2797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=384310 $D=103
M1469 2799 WL_189 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=384800 $D=103
M1470 2419 WL_190 2801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=387710 $D=103
M1471 2803 WL_191 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=388200 $D=103
M1472 2419 WL_192 2805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=391110 $D=103
M1473 2807 WL_193 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=391600 $D=103
M1474 2419 WL_194 2809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=394510 $D=103
M1475 2811 WL_195 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=395000 $D=103
M1476 2419 WL_196 2813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=397910 $D=103
M1477 2815 WL_197 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=398400 $D=103
M1478 2419 WL_198 2817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=401310 $D=103
M1479 2819 WL_199 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=401800 $D=103
M1480 2419 WL_200 2821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=404710 $D=103
M1481 2823 WL_201 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=405200 $D=103
M1482 2419 WL_202 2825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=408110 $D=103
M1483 2827 WL_203 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=408600 $D=103
M1484 2419 WL_204 2829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=411510 $D=103
M1485 2831 WL_205 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=412000 $D=103
M1486 2419 WL_206 2833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=414910 $D=103
M1487 2835 WL_207 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=415400 $D=103
M1488 2419 WL_208 2837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=418310 $D=103
M1489 2839 WL_209 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=418800 $D=103
M1490 2419 WL_210 2841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=421710 $D=103
M1491 2843 WL_211 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=422200 $D=103
M1492 2419 WL_212 2845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=425110 $D=103
M1493 2847 WL_213 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=425600 $D=103
M1494 2419 WL_214 2849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=428510 $D=103
M1495 2851 WL_215 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=429000 $D=103
M1496 2419 WL_216 2853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=431910 $D=103
M1497 2855 WL_217 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=432400 $D=103
M1498 2419 WL_218 2857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=435310 $D=103
M1499 2859 WL_219 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=435800 $D=103
M1500 2419 WL_220 2861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=438710 $D=103
M1501 2863 WL_221 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=439200 $D=103
M1502 2419 WL_222 2865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=442110 $D=103
M1503 2867 WL_223 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=442600 $D=103
M1504 2419 WL_224 2869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=445510 $D=103
M1505 2871 WL_225 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=446000 $D=103
M1506 2419 WL_226 2873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=448910 $D=103
M1507 2875 WL_227 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=449400 $D=103
M1508 2419 WL_228 2877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=452310 $D=103
M1509 2879 WL_229 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=452800 $D=103
M1510 2419 WL_230 2881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=455710 $D=103
M1511 2883 WL_231 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=456200 $D=103
M1512 2419 WL_232 2885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=459110 $D=103
M1513 2887 WL_233 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=459600 $D=103
M1514 2419 WL_234 2889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=462510 $D=103
M1515 2891 WL_235 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=463000 $D=103
M1516 2419 WL_236 2893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=465910 $D=103
M1517 2895 WL_237 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=466400 $D=103
M1518 2419 WL_238 2897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=469310 $D=103
M1519 2899 WL_239 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=469800 $D=103
M1520 2419 WL_240 2901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=472710 $D=103
M1521 2903 WL_241 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=473200 $D=103
M1522 2419 WL_242 2905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=476110 $D=103
M1523 2907 WL_243 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=476600 $D=103
M1524 2419 WL_244 2909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=479510 $D=103
M1525 2911 WL_245 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=480000 $D=103
M1526 2419 WL_246 2913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=482910 $D=103
M1527 2915 WL_247 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=483400 $D=103
M1528 2419 WL_248 2917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=486310 $D=103
M1529 2919 WL_249 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=486800 $D=103
M1530 2419 WL_250 2921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=489710 $D=103
M1531 2923 WL_251 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=490200 $D=103
M1532 2419 WL_252 2925 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=493110 $D=103
M1533 2927 WL_253 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=493600 $D=103
M1534 2419 WL_254 2929 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=496510 $D=103
M1535 2931 WL_255 2419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58890 $Y=497000 $D=103
M1536 2420 WL_0 2422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=64710 $D=103
M1537 2424 WL_1 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=65200 $D=103
M1538 2420 WL_2 2426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=68110 $D=103
M1539 2428 WL_3 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=68600 $D=103
M1540 2420 WL_4 2430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=71510 $D=103
M1541 2432 WL_5 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=72000 $D=103
M1542 2420 WL_6 2434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=74910 $D=103
M1543 2436 WL_7 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=75400 $D=103
M1544 2420 WL_8 2438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=78310 $D=103
M1545 2440 WL_9 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=78800 $D=103
M1546 2420 WL_10 2442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=81710 $D=103
M1547 2444 WL_11 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=82200 $D=103
M1548 2420 WL_12 2446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=85110 $D=103
M1549 2448 WL_13 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=85600 $D=103
M1550 2420 WL_14 2450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=88510 $D=103
M1551 2452 WL_15 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=89000 $D=103
M1552 2420 WL_16 2454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=91910 $D=103
M1553 2456 WL_17 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=92400 $D=103
M1554 2420 WL_18 2458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=95310 $D=103
M1555 2460 WL_19 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=95800 $D=103
M1556 2420 WL_20 2462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=98710 $D=103
M1557 2464 WL_21 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=99200 $D=103
M1558 2420 WL_22 2466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=102110 $D=103
M1559 2468 WL_23 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=102600 $D=103
M1560 2420 WL_24 2470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=105510 $D=103
M1561 2472 WL_25 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=106000 $D=103
M1562 2420 WL_26 2474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=108910 $D=103
M1563 2476 WL_27 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=109400 $D=103
M1564 2420 WL_28 2478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=112310 $D=103
M1565 2480 WL_29 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=112800 $D=103
M1566 2420 WL_30 2482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=115710 $D=103
M1567 2484 WL_31 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=116200 $D=103
M1568 2420 WL_32 2486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=119110 $D=103
M1569 2488 WL_33 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=119600 $D=103
M1570 2420 WL_34 2490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=122510 $D=103
M1571 2492 WL_35 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=123000 $D=103
M1572 2420 WL_36 2494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=125910 $D=103
M1573 2496 WL_37 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=126400 $D=103
M1574 2420 WL_38 2498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=129310 $D=103
M1575 2500 WL_39 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=129800 $D=103
M1576 2420 WL_40 2502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=132710 $D=103
M1577 2504 WL_41 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=133200 $D=103
M1578 2420 WL_42 2506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=136110 $D=103
M1579 2508 WL_43 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=136600 $D=103
M1580 2420 WL_44 2510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=139510 $D=103
M1581 2512 WL_45 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=140000 $D=103
M1582 2420 WL_46 2514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=142910 $D=103
M1583 2516 WL_47 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=143400 $D=103
M1584 2420 WL_48 2518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=146310 $D=103
M1585 2520 WL_49 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=146800 $D=103
M1586 2420 WL_50 2522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=149710 $D=103
M1587 2524 WL_51 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=150200 $D=103
M1588 2420 WL_52 2526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=153110 $D=103
M1589 2528 WL_53 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=153600 $D=103
M1590 2420 WL_54 2530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=156510 $D=103
M1591 2532 WL_55 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=157000 $D=103
M1592 2420 WL_56 2534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=159910 $D=103
M1593 2536 WL_57 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=160400 $D=103
M1594 2420 WL_58 2538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=163310 $D=103
M1595 2540 WL_59 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=163800 $D=103
M1596 2420 WL_60 2542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=166710 $D=103
M1597 2544 WL_61 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=167200 $D=103
M1598 2420 WL_62 2546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=170110 $D=103
M1599 2548 WL_63 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=170600 $D=103
M1600 2420 WL_64 2550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=173510 $D=103
M1601 2552 WL_65 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=174000 $D=103
M1602 2420 WL_66 2554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=176910 $D=103
M1603 2556 WL_67 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=177400 $D=103
M1604 2420 WL_68 2558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=180310 $D=103
M1605 2560 WL_69 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=180800 $D=103
M1606 2420 WL_70 2562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=183710 $D=103
M1607 2564 WL_71 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=184200 $D=103
M1608 2420 WL_72 2566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=187110 $D=103
M1609 2568 WL_73 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=187600 $D=103
M1610 2420 WL_74 2570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=190510 $D=103
M1611 2572 WL_75 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=191000 $D=103
M1612 2420 WL_76 2574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=193910 $D=103
M1613 2576 WL_77 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=194400 $D=103
M1614 2420 WL_78 2578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=197310 $D=103
M1615 2580 WL_79 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=197800 $D=103
M1616 2420 WL_80 2582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=200710 $D=103
M1617 2584 WL_81 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=201200 $D=103
M1618 2420 WL_82 2586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=204110 $D=103
M1619 2588 WL_83 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=204600 $D=103
M1620 2420 WL_84 2590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=207510 $D=103
M1621 2592 WL_85 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=208000 $D=103
M1622 2420 WL_86 2594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=210910 $D=103
M1623 2596 WL_87 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=211400 $D=103
M1624 2420 WL_88 2598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=214310 $D=103
M1625 2600 WL_89 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=214800 $D=103
M1626 2420 WL_90 2602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=217710 $D=103
M1627 2604 WL_91 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=218200 $D=103
M1628 2420 WL_92 2606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=221110 $D=103
M1629 2608 WL_93 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=221600 $D=103
M1630 2420 WL_94 2610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=224510 $D=103
M1631 2612 WL_95 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=225000 $D=103
M1632 2420 WL_96 2614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=227910 $D=103
M1633 2616 WL_97 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=228400 $D=103
M1634 2420 WL_98 2618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=231310 $D=103
M1635 2620 WL_99 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=231800 $D=103
M1636 2420 WL_100 2622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=234710 $D=103
M1637 2624 WL_101 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=235200 $D=103
M1638 2420 WL_102 2626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=238110 $D=103
M1639 2628 WL_103 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=238600 $D=103
M1640 2420 WL_104 2630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=241510 $D=103
M1641 2632 WL_105 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=242000 $D=103
M1642 2420 WL_106 2634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=244910 $D=103
M1643 2636 WL_107 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=245400 $D=103
M1644 2420 WL_108 2638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=248310 $D=103
M1645 2640 WL_109 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=248800 $D=103
M1646 2420 WL_110 2642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=251710 $D=103
M1647 2644 WL_111 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=252200 $D=103
M1648 2420 WL_112 2646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=255110 $D=103
M1649 2648 WL_113 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=255600 $D=103
M1650 2420 WL_114 2650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=258510 $D=103
M1651 2652 WL_115 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=259000 $D=103
M1652 2420 WL_116 2654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=261910 $D=103
M1653 2656 WL_117 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=262400 $D=103
M1654 2420 WL_118 2658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=265310 $D=103
M1655 2660 WL_119 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=265800 $D=103
M1656 2420 WL_120 2662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=268710 $D=103
M1657 2664 WL_121 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=269200 $D=103
M1658 2420 WL_122 2666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=272110 $D=103
M1659 2668 WL_123 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=272600 $D=103
M1660 2420 WL_124 2670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=275510 $D=103
M1661 2672 WL_125 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=276000 $D=103
M1662 2420 WL_126 2674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=278910 $D=103
M1663 2676 WL_127 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=279400 $D=103
M1664 2420 WL_128 2678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=282310 $D=103
M1665 2680 WL_129 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=282800 $D=103
M1666 2420 WL_130 2682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=285710 $D=103
M1667 2684 WL_131 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=286200 $D=103
M1668 2420 WL_132 2686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=289110 $D=103
M1669 2688 WL_133 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=289600 $D=103
M1670 2420 WL_134 2690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=292510 $D=103
M1671 2692 WL_135 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=293000 $D=103
M1672 2420 WL_136 2694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=295910 $D=103
M1673 2696 WL_137 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=296400 $D=103
M1674 2420 WL_138 2698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=299310 $D=103
M1675 2700 WL_139 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=299800 $D=103
M1676 2420 WL_140 2702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=302710 $D=103
M1677 2704 WL_141 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=303200 $D=103
M1678 2420 WL_142 2706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=306110 $D=103
M1679 2708 WL_143 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=306600 $D=103
M1680 2420 WL_144 2710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=309510 $D=103
M1681 2712 WL_145 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=310000 $D=103
M1682 2420 WL_146 2714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=312910 $D=103
M1683 2716 WL_147 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=313400 $D=103
M1684 2420 WL_148 2718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=316310 $D=103
M1685 2720 WL_149 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=316800 $D=103
M1686 2420 WL_150 2722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=319710 $D=103
M1687 2724 WL_151 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=320200 $D=103
M1688 2420 WL_152 2726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=323110 $D=103
M1689 2728 WL_153 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=323600 $D=103
M1690 2420 WL_154 2730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=326510 $D=103
M1691 2732 WL_155 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=327000 $D=103
M1692 2420 WL_156 2734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=329910 $D=103
M1693 2736 WL_157 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=330400 $D=103
M1694 2420 WL_158 2738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=333310 $D=103
M1695 2740 WL_159 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=333800 $D=103
M1696 2420 WL_160 2742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=336710 $D=103
M1697 2744 WL_161 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=337200 $D=103
M1698 2420 WL_162 2746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=340110 $D=103
M1699 2748 WL_163 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=340600 $D=103
M1700 2420 WL_164 2750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=343510 $D=103
M1701 2752 WL_165 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=344000 $D=103
M1702 2420 WL_166 2754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=346910 $D=103
M1703 2756 WL_167 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=347400 $D=103
M1704 2420 WL_168 2758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=350310 $D=103
M1705 2760 WL_169 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=350800 $D=103
M1706 2420 WL_170 2762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=353710 $D=103
M1707 2764 WL_171 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=354200 $D=103
M1708 2420 WL_172 2766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=357110 $D=103
M1709 2768 WL_173 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=357600 $D=103
M1710 2420 WL_174 2770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=360510 $D=103
M1711 2772 WL_175 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=361000 $D=103
M1712 2420 WL_176 2774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=363910 $D=103
M1713 2776 WL_177 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=364400 $D=103
M1714 2420 WL_178 2778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=367310 $D=103
M1715 2780 WL_179 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=367800 $D=103
M1716 2420 WL_180 2782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=370710 $D=103
M1717 2784 WL_181 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=371200 $D=103
M1718 2420 WL_182 2786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=374110 $D=103
M1719 2788 WL_183 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=374600 $D=103
M1720 2420 WL_184 2790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=377510 $D=103
M1721 2792 WL_185 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=378000 $D=103
M1722 2420 WL_186 2794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=380910 $D=103
M1723 2796 WL_187 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=381400 $D=103
M1724 2420 WL_188 2798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=384310 $D=103
M1725 2800 WL_189 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=384800 $D=103
M1726 2420 WL_190 2802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=387710 $D=103
M1727 2804 WL_191 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=388200 $D=103
M1728 2420 WL_192 2806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=391110 $D=103
M1729 2808 WL_193 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=391600 $D=103
M1730 2420 WL_194 2810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=394510 $D=103
M1731 2812 WL_195 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=395000 $D=103
M1732 2420 WL_196 2814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=397910 $D=103
M1733 2816 WL_197 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=398400 $D=103
M1734 2420 WL_198 2818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=401310 $D=103
M1735 2820 WL_199 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=401800 $D=103
M1736 2420 WL_200 2822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=404710 $D=103
M1737 2824 WL_201 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=405200 $D=103
M1738 2420 WL_202 2826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=408110 $D=103
M1739 2828 WL_203 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=408600 $D=103
M1740 2420 WL_204 2830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=411510 $D=103
M1741 2832 WL_205 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=412000 $D=103
M1742 2420 WL_206 2834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=414910 $D=103
M1743 2836 WL_207 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=415400 $D=103
M1744 2420 WL_208 2838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=418310 $D=103
M1745 2840 WL_209 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=418800 $D=103
M1746 2420 WL_210 2842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=421710 $D=103
M1747 2844 WL_211 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=422200 $D=103
M1748 2420 WL_212 2846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=425110 $D=103
M1749 2848 WL_213 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=425600 $D=103
M1750 2420 WL_214 2850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=428510 $D=103
M1751 2852 WL_215 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=429000 $D=103
M1752 2420 WL_216 2854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=431910 $D=103
M1753 2856 WL_217 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=432400 $D=103
M1754 2420 WL_218 2858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=435310 $D=103
M1755 2860 WL_219 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=435800 $D=103
M1756 2420 WL_220 2862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=438710 $D=103
M1757 2864 WL_221 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=439200 $D=103
M1758 2420 WL_222 2866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=442110 $D=103
M1759 2868 WL_223 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=442600 $D=103
M1760 2420 WL_224 2870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=445510 $D=103
M1761 2872 WL_225 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=446000 $D=103
M1762 2420 WL_226 2874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=448910 $D=103
M1763 2876 WL_227 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=449400 $D=103
M1764 2420 WL_228 2878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=452310 $D=103
M1765 2880 WL_229 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=452800 $D=103
M1766 2420 WL_230 2882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=455710 $D=103
M1767 2884 WL_231 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=456200 $D=103
M1768 2420 WL_232 2886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=459110 $D=103
M1769 2888 WL_233 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=459600 $D=103
M1770 2420 WL_234 2890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=462510 $D=103
M1771 2892 WL_235 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=463000 $D=103
M1772 2420 WL_236 2894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=465910 $D=103
M1773 2896 WL_237 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=466400 $D=103
M1774 2420 WL_238 2898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=469310 $D=103
M1775 2900 WL_239 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=469800 $D=103
M1776 2420 WL_240 2902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=472710 $D=103
M1777 2904 WL_241 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=473200 $D=103
M1778 2420 WL_242 2906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=476110 $D=103
M1779 2908 WL_243 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=476600 $D=103
M1780 2420 WL_244 2910 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=479510 $D=103
M1781 2912 WL_245 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=480000 $D=103
M1782 2420 WL_246 2914 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=482910 $D=103
M1783 2916 WL_247 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=483400 $D=103
M1784 2420 WL_248 2918 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=486310 $D=103
M1785 2920 WL_249 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=486800 $D=103
M1786 2420 WL_250 2922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=489710 $D=103
M1787 2924 WL_251 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=490200 $D=103
M1788 2420 WL_252 2926 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=493110 $D=103
M1789 2928 WL_253 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=493600 $D=103
M1790 2420 WL_254 2930 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=496510 $D=103
M1791 2932 WL_255 2420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77750 $Y=497000 $D=103
M1792 2934 WL_0 2935 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=64710 $D=103
M1793 2937 WL_1 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=65200 $D=103
M1794 2934 WL_2 2939 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=68110 $D=103
M1795 2941 WL_3 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=68600 $D=103
M1796 2934 WL_4 2943 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=71510 $D=103
M1797 2945 WL_5 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=72000 $D=103
M1798 2934 WL_6 2947 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=74910 $D=103
M1799 2949 WL_7 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=75400 $D=103
M1800 2934 WL_8 2951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=78310 $D=103
M1801 2953 WL_9 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=78800 $D=103
M1802 2934 WL_10 2955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=81710 $D=103
M1803 2957 WL_11 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=82200 $D=103
M1804 2934 WL_12 2959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=85110 $D=103
M1805 2961 WL_13 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=85600 $D=103
M1806 2934 WL_14 2963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=88510 $D=103
M1807 2965 WL_15 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=89000 $D=103
M1808 2934 WL_16 2967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=91910 $D=103
M1809 2969 WL_17 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=92400 $D=103
M1810 2934 WL_18 2971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=95310 $D=103
M1811 2973 WL_19 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=95800 $D=103
M1812 2934 WL_20 2975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=98710 $D=103
M1813 2977 WL_21 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=99200 $D=103
M1814 2934 WL_22 2979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=102110 $D=103
M1815 2981 WL_23 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=102600 $D=103
M1816 2934 WL_24 2983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=105510 $D=103
M1817 2985 WL_25 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=106000 $D=103
M1818 2934 WL_26 2987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=108910 $D=103
M1819 2989 WL_27 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=109400 $D=103
M1820 2934 WL_28 2991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=112310 $D=103
M1821 2993 WL_29 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=112800 $D=103
M1822 2934 WL_30 2995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=115710 $D=103
M1823 2997 WL_31 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=116200 $D=103
M1824 2934 WL_32 2999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=119110 $D=103
M1825 3001 WL_33 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=119600 $D=103
M1826 2934 WL_34 3003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=122510 $D=103
M1827 3005 WL_35 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=123000 $D=103
M1828 2934 WL_36 3007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=125910 $D=103
M1829 3009 WL_37 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=126400 $D=103
M1830 2934 WL_38 3011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=129310 $D=103
M1831 3013 WL_39 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=129800 $D=103
M1832 2934 WL_40 3015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=132710 $D=103
M1833 3017 WL_41 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=133200 $D=103
M1834 2934 WL_42 3019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=136110 $D=103
M1835 3021 WL_43 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=136600 $D=103
M1836 2934 WL_44 3023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=139510 $D=103
M1837 3025 WL_45 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=140000 $D=103
M1838 2934 WL_46 3027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=142910 $D=103
M1839 3029 WL_47 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=143400 $D=103
M1840 2934 WL_48 3031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=146310 $D=103
M1841 3033 WL_49 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=146800 $D=103
M1842 2934 WL_50 3035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=149710 $D=103
M1843 3037 WL_51 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=150200 $D=103
M1844 2934 WL_52 3039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=153110 $D=103
M1845 3041 WL_53 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=153600 $D=103
M1846 2934 WL_54 3043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=156510 $D=103
M1847 3045 WL_55 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=157000 $D=103
M1848 2934 WL_56 3047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=159910 $D=103
M1849 3049 WL_57 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=160400 $D=103
M1850 2934 WL_58 3051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=163310 $D=103
M1851 3053 WL_59 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=163800 $D=103
M1852 2934 WL_60 3055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=166710 $D=103
M1853 3057 WL_61 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=167200 $D=103
M1854 2934 WL_62 3059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=170110 $D=103
M1855 3061 WL_63 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=170600 $D=103
M1856 2934 WL_64 3063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=173510 $D=103
M1857 3065 WL_65 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=174000 $D=103
M1858 2934 WL_66 3067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=176910 $D=103
M1859 3069 WL_67 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=177400 $D=103
M1860 2934 WL_68 3071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=180310 $D=103
M1861 3073 WL_69 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=180800 $D=103
M1862 2934 WL_70 3075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=183710 $D=103
M1863 3077 WL_71 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=184200 $D=103
M1864 2934 WL_72 3079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=187110 $D=103
M1865 3081 WL_73 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=187600 $D=103
M1866 2934 WL_74 3083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=190510 $D=103
M1867 3085 WL_75 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=191000 $D=103
M1868 2934 WL_76 3087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=193910 $D=103
M1869 3089 WL_77 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=194400 $D=103
M1870 2934 WL_78 3091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=197310 $D=103
M1871 3093 WL_79 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=197800 $D=103
M1872 2934 WL_80 3095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=200710 $D=103
M1873 3097 WL_81 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=201200 $D=103
M1874 2934 WL_82 3099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=204110 $D=103
M1875 3101 WL_83 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=204600 $D=103
M1876 2934 WL_84 3103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=207510 $D=103
M1877 3105 WL_85 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=208000 $D=103
M1878 2934 WL_86 3107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=210910 $D=103
M1879 3109 WL_87 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=211400 $D=103
M1880 2934 WL_88 3111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=214310 $D=103
M1881 3113 WL_89 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=214800 $D=103
M1882 2934 WL_90 3115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=217710 $D=103
M1883 3117 WL_91 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=218200 $D=103
M1884 2934 WL_92 3119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=221110 $D=103
M1885 3121 WL_93 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=221600 $D=103
M1886 2934 WL_94 3123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=224510 $D=103
M1887 3125 WL_95 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=225000 $D=103
M1888 2934 WL_96 3127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=227910 $D=103
M1889 3129 WL_97 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=228400 $D=103
M1890 2934 WL_98 3131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=231310 $D=103
M1891 3133 WL_99 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=231800 $D=103
M1892 2934 WL_100 3135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=234710 $D=103
M1893 3137 WL_101 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=235200 $D=103
M1894 2934 WL_102 3139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=238110 $D=103
M1895 3141 WL_103 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=238600 $D=103
M1896 2934 WL_104 3143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=241510 $D=103
M1897 3145 WL_105 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=242000 $D=103
M1898 2934 WL_106 3147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=244910 $D=103
M1899 3149 WL_107 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=245400 $D=103
M1900 2934 WL_108 3151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=248310 $D=103
M1901 3153 WL_109 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=248800 $D=103
M1902 2934 WL_110 3155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=251710 $D=103
M1903 3157 WL_111 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=252200 $D=103
M1904 2934 WL_112 3159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=255110 $D=103
M1905 3161 WL_113 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=255600 $D=103
M1906 2934 WL_114 3163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=258510 $D=103
M1907 3165 WL_115 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=259000 $D=103
M1908 2934 WL_116 3167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=261910 $D=103
M1909 3169 WL_117 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=262400 $D=103
M1910 2934 WL_118 3171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=265310 $D=103
M1911 3173 WL_119 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=265800 $D=103
M1912 2934 WL_120 3175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=268710 $D=103
M1913 3177 WL_121 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=269200 $D=103
M1914 2934 WL_122 3179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=272110 $D=103
M1915 3181 WL_123 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=272600 $D=103
M1916 2934 WL_124 3183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=275510 $D=103
M1917 3185 WL_125 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=276000 $D=103
M1918 2934 WL_126 3187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=278910 $D=103
M1919 3189 WL_127 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=279400 $D=103
M1920 2934 WL_128 3191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=282310 $D=103
M1921 3193 WL_129 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=282800 $D=103
M1922 2934 WL_130 3195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=285710 $D=103
M1923 3197 WL_131 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=286200 $D=103
M1924 2934 WL_132 3199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=289110 $D=103
M1925 3201 WL_133 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=289600 $D=103
M1926 2934 WL_134 3203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=292510 $D=103
M1927 3205 WL_135 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=293000 $D=103
M1928 2934 WL_136 3207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=295910 $D=103
M1929 3209 WL_137 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=296400 $D=103
M1930 2934 WL_138 3211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=299310 $D=103
M1931 3213 WL_139 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=299800 $D=103
M1932 2934 WL_140 3215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=302710 $D=103
M1933 3217 WL_141 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=303200 $D=103
M1934 2934 WL_142 3219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=306110 $D=103
M1935 3221 WL_143 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=306600 $D=103
M1936 2934 WL_144 3223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=309510 $D=103
M1937 3225 WL_145 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=310000 $D=103
M1938 2934 WL_146 3227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=312910 $D=103
M1939 3229 WL_147 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=313400 $D=103
M1940 2934 WL_148 3231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=316310 $D=103
M1941 3233 WL_149 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=316800 $D=103
M1942 2934 WL_150 3235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=319710 $D=103
M1943 3237 WL_151 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=320200 $D=103
M1944 2934 WL_152 3239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=323110 $D=103
M1945 3241 WL_153 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=323600 $D=103
M1946 2934 WL_154 3243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=326510 $D=103
M1947 3245 WL_155 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=327000 $D=103
M1948 2934 WL_156 3247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=329910 $D=103
M1949 3249 WL_157 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=330400 $D=103
M1950 2934 WL_158 3251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=333310 $D=103
M1951 3253 WL_159 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=333800 $D=103
M1952 2934 WL_160 3255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=336710 $D=103
M1953 3257 WL_161 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=337200 $D=103
M1954 2934 WL_162 3259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=340110 $D=103
M1955 3261 WL_163 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=340600 $D=103
M1956 2934 WL_164 3263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=343510 $D=103
M1957 3265 WL_165 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=344000 $D=103
M1958 2934 WL_166 3267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=346910 $D=103
M1959 3269 WL_167 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=347400 $D=103
M1960 2934 WL_168 3271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=350310 $D=103
M1961 3273 WL_169 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=350800 $D=103
M1962 2934 WL_170 3275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=353710 $D=103
M1963 3277 WL_171 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=354200 $D=103
M1964 2934 WL_172 3279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=357110 $D=103
M1965 3281 WL_173 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=357600 $D=103
M1966 2934 WL_174 3283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=360510 $D=103
M1967 3285 WL_175 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=361000 $D=103
M1968 2934 WL_176 3287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=363910 $D=103
M1969 3289 WL_177 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=364400 $D=103
M1970 2934 WL_178 3291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=367310 $D=103
M1971 3293 WL_179 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=367800 $D=103
M1972 2934 WL_180 3295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=370710 $D=103
M1973 3297 WL_181 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=371200 $D=103
M1974 2934 WL_182 3299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=374110 $D=103
M1975 3301 WL_183 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=374600 $D=103
M1976 2934 WL_184 3303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=377510 $D=103
M1977 3305 WL_185 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=378000 $D=103
M1978 2934 WL_186 3307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=380910 $D=103
M1979 3309 WL_187 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=381400 $D=103
M1980 2934 WL_188 3311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=384310 $D=103
M1981 3313 WL_189 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=384800 $D=103
M1982 2934 WL_190 3315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=387710 $D=103
M1983 3317 WL_191 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=388200 $D=103
M1984 2934 WL_192 3319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=391110 $D=103
M1985 3321 WL_193 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=391600 $D=103
M1986 2934 WL_194 3323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=394510 $D=103
M1987 3325 WL_195 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=395000 $D=103
M1988 2934 WL_196 3327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=397910 $D=103
M1989 3329 WL_197 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=398400 $D=103
M1990 2934 WL_198 3331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=401310 $D=103
M1991 3333 WL_199 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=401800 $D=103
M1992 2934 WL_200 3335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=404710 $D=103
M1993 3337 WL_201 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=405200 $D=103
M1994 2934 WL_202 3339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=408110 $D=103
M1995 3341 WL_203 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=408600 $D=103
M1996 2934 WL_204 3343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=411510 $D=103
M1997 3345 WL_205 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=412000 $D=103
M1998 2934 WL_206 3347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=414910 $D=103
M1999 3349 WL_207 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=415400 $D=103
M2000 2934 WL_208 3351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=418310 $D=103
M2001 3353 WL_209 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=418800 $D=103
M2002 2934 WL_210 3355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=421710 $D=103
M2003 3357 WL_211 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=422200 $D=103
M2004 2934 WL_212 3359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=425110 $D=103
M2005 3361 WL_213 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=425600 $D=103
M2006 2934 WL_214 3363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=428510 $D=103
M2007 3365 WL_215 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=429000 $D=103
M2008 2934 WL_216 3367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=431910 $D=103
M2009 3369 WL_217 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=432400 $D=103
M2010 2934 WL_218 3371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=435310 $D=103
M2011 3373 WL_219 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=435800 $D=103
M2012 2934 WL_220 3375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=438710 $D=103
M2013 3377 WL_221 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=439200 $D=103
M2014 2934 WL_222 3379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=442110 $D=103
M2015 3381 WL_223 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=442600 $D=103
M2016 2934 WL_224 3383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=445510 $D=103
M2017 3385 WL_225 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=446000 $D=103
M2018 2934 WL_226 3387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=448910 $D=103
M2019 3389 WL_227 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=449400 $D=103
M2020 2934 WL_228 3391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=452310 $D=103
M2021 3393 WL_229 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=452800 $D=103
M2022 2934 WL_230 3395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=455710 $D=103
M2023 3397 WL_231 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=456200 $D=103
M2024 2934 WL_232 3399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=459110 $D=103
M2025 3401 WL_233 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=459600 $D=103
M2026 2934 WL_234 3403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=462510 $D=103
M2027 3405 WL_235 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=463000 $D=103
M2028 2934 WL_236 3407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=465910 $D=103
M2029 3409 WL_237 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=466400 $D=103
M2030 2934 WL_238 3411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=469310 $D=103
M2031 3413 WL_239 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=469800 $D=103
M2032 2934 WL_240 3415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=472710 $D=103
M2033 3417 WL_241 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=473200 $D=103
M2034 2934 WL_242 3419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=476110 $D=103
M2035 3421 WL_243 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=476600 $D=103
M2036 2934 WL_244 3423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=479510 $D=103
M2037 3425 WL_245 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=480000 $D=103
M2038 2934 WL_246 3427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=482910 $D=103
M2039 3429 WL_247 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=483400 $D=103
M2040 2934 WL_248 3431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=486310 $D=103
M2041 3433 WL_249 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=486800 $D=103
M2042 2934 WL_250 3435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=489710 $D=103
M2043 3437 WL_251 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=490200 $D=103
M2044 2934 WL_252 3439 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=493110 $D=103
M2045 3441 WL_253 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=493600 $D=103
M2046 2934 WL_254 3443 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=496510 $D=103
M2047 3445 WL_255 2934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79290 $Y=497000 $D=103
M2048 2933 WL_0 2936 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=64710 $D=103
M2049 2938 WL_1 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=65200 $D=103
M2050 2933 WL_2 2940 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=68110 $D=103
M2051 2942 WL_3 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=68600 $D=103
M2052 2933 WL_4 2944 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=71510 $D=103
M2053 2946 WL_5 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=72000 $D=103
M2054 2933 WL_6 2948 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=74910 $D=103
M2055 2950 WL_7 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=75400 $D=103
M2056 2933 WL_8 2952 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=78310 $D=103
M2057 2954 WL_9 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=78800 $D=103
M2058 2933 WL_10 2956 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=81710 $D=103
M2059 2958 WL_11 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=82200 $D=103
M2060 2933 WL_12 2960 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=85110 $D=103
M2061 2962 WL_13 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=85600 $D=103
M2062 2933 WL_14 2964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=88510 $D=103
M2063 2966 WL_15 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=89000 $D=103
M2064 2933 WL_16 2968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=91910 $D=103
M2065 2970 WL_17 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=92400 $D=103
M2066 2933 WL_18 2972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=95310 $D=103
M2067 2974 WL_19 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=95800 $D=103
M2068 2933 WL_20 2976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=98710 $D=103
M2069 2978 WL_21 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=99200 $D=103
M2070 2933 WL_22 2980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=102110 $D=103
M2071 2982 WL_23 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=102600 $D=103
M2072 2933 WL_24 2984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=105510 $D=103
M2073 2986 WL_25 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=106000 $D=103
M2074 2933 WL_26 2988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=108910 $D=103
M2075 2990 WL_27 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=109400 $D=103
M2076 2933 WL_28 2992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=112310 $D=103
M2077 2994 WL_29 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=112800 $D=103
M2078 2933 WL_30 2996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=115710 $D=103
M2079 2998 WL_31 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=116200 $D=103
M2080 2933 WL_32 3000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=119110 $D=103
M2081 3002 WL_33 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=119600 $D=103
M2082 2933 WL_34 3004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=122510 $D=103
M2083 3006 WL_35 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=123000 $D=103
M2084 2933 WL_36 3008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=125910 $D=103
M2085 3010 WL_37 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=126400 $D=103
M2086 2933 WL_38 3012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=129310 $D=103
M2087 3014 WL_39 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=129800 $D=103
M2088 2933 WL_40 3016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=132710 $D=103
M2089 3018 WL_41 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=133200 $D=103
M2090 2933 WL_42 3020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=136110 $D=103
M2091 3022 WL_43 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=136600 $D=103
M2092 2933 WL_44 3024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=139510 $D=103
M2093 3026 WL_45 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=140000 $D=103
M2094 2933 WL_46 3028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=142910 $D=103
M2095 3030 WL_47 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=143400 $D=103
M2096 2933 WL_48 3032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=146310 $D=103
M2097 3034 WL_49 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=146800 $D=103
M2098 2933 WL_50 3036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=149710 $D=103
M2099 3038 WL_51 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=150200 $D=103
M2100 2933 WL_52 3040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=153110 $D=103
M2101 3042 WL_53 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=153600 $D=103
M2102 2933 WL_54 3044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=156510 $D=103
M2103 3046 WL_55 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=157000 $D=103
M2104 2933 WL_56 3048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=159910 $D=103
M2105 3050 WL_57 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=160400 $D=103
M2106 2933 WL_58 3052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=163310 $D=103
M2107 3054 WL_59 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=163800 $D=103
M2108 2933 WL_60 3056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=166710 $D=103
M2109 3058 WL_61 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=167200 $D=103
M2110 2933 WL_62 3060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=170110 $D=103
M2111 3062 WL_63 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=170600 $D=103
M2112 2933 WL_64 3064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=173510 $D=103
M2113 3066 WL_65 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=174000 $D=103
M2114 2933 WL_66 3068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=176910 $D=103
M2115 3070 WL_67 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=177400 $D=103
M2116 2933 WL_68 3072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=180310 $D=103
M2117 3074 WL_69 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=180800 $D=103
M2118 2933 WL_70 3076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=183710 $D=103
M2119 3078 WL_71 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=184200 $D=103
M2120 2933 WL_72 3080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=187110 $D=103
M2121 3082 WL_73 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=187600 $D=103
M2122 2933 WL_74 3084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=190510 $D=103
M2123 3086 WL_75 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=191000 $D=103
M2124 2933 WL_76 3088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=193910 $D=103
M2125 3090 WL_77 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=194400 $D=103
M2126 2933 WL_78 3092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=197310 $D=103
M2127 3094 WL_79 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=197800 $D=103
M2128 2933 WL_80 3096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=200710 $D=103
M2129 3098 WL_81 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=201200 $D=103
M2130 2933 WL_82 3100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=204110 $D=103
M2131 3102 WL_83 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=204600 $D=103
M2132 2933 WL_84 3104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=207510 $D=103
M2133 3106 WL_85 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=208000 $D=103
M2134 2933 WL_86 3108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=210910 $D=103
M2135 3110 WL_87 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=211400 $D=103
M2136 2933 WL_88 3112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=214310 $D=103
M2137 3114 WL_89 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=214800 $D=103
M2138 2933 WL_90 3116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=217710 $D=103
M2139 3118 WL_91 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=218200 $D=103
M2140 2933 WL_92 3120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=221110 $D=103
M2141 3122 WL_93 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=221600 $D=103
M2142 2933 WL_94 3124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=224510 $D=103
M2143 3126 WL_95 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=225000 $D=103
M2144 2933 WL_96 3128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=227910 $D=103
M2145 3130 WL_97 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=228400 $D=103
M2146 2933 WL_98 3132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=231310 $D=103
M2147 3134 WL_99 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=231800 $D=103
M2148 2933 WL_100 3136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=234710 $D=103
M2149 3138 WL_101 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=235200 $D=103
M2150 2933 WL_102 3140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=238110 $D=103
M2151 3142 WL_103 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=238600 $D=103
M2152 2933 WL_104 3144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=241510 $D=103
M2153 3146 WL_105 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=242000 $D=103
M2154 2933 WL_106 3148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=244910 $D=103
M2155 3150 WL_107 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=245400 $D=103
M2156 2933 WL_108 3152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=248310 $D=103
M2157 3154 WL_109 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=248800 $D=103
M2158 2933 WL_110 3156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=251710 $D=103
M2159 3158 WL_111 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=252200 $D=103
M2160 2933 WL_112 3160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=255110 $D=103
M2161 3162 WL_113 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=255600 $D=103
M2162 2933 WL_114 3164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=258510 $D=103
M2163 3166 WL_115 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=259000 $D=103
M2164 2933 WL_116 3168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=261910 $D=103
M2165 3170 WL_117 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=262400 $D=103
M2166 2933 WL_118 3172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=265310 $D=103
M2167 3174 WL_119 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=265800 $D=103
M2168 2933 WL_120 3176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=268710 $D=103
M2169 3178 WL_121 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=269200 $D=103
M2170 2933 WL_122 3180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=272110 $D=103
M2171 3182 WL_123 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=272600 $D=103
M2172 2933 WL_124 3184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=275510 $D=103
M2173 3186 WL_125 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=276000 $D=103
M2174 2933 WL_126 3188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=278910 $D=103
M2175 3190 WL_127 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=279400 $D=103
M2176 2933 WL_128 3192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=282310 $D=103
M2177 3194 WL_129 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=282800 $D=103
M2178 2933 WL_130 3196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=285710 $D=103
M2179 3198 WL_131 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=286200 $D=103
M2180 2933 WL_132 3200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=289110 $D=103
M2181 3202 WL_133 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=289600 $D=103
M2182 2933 WL_134 3204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=292510 $D=103
M2183 3206 WL_135 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=293000 $D=103
M2184 2933 WL_136 3208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=295910 $D=103
M2185 3210 WL_137 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=296400 $D=103
M2186 2933 WL_138 3212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=299310 $D=103
M2187 3214 WL_139 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=299800 $D=103
M2188 2933 WL_140 3216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=302710 $D=103
M2189 3218 WL_141 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=303200 $D=103
M2190 2933 WL_142 3220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=306110 $D=103
M2191 3222 WL_143 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=306600 $D=103
M2192 2933 WL_144 3224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=309510 $D=103
M2193 3226 WL_145 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=310000 $D=103
M2194 2933 WL_146 3228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=312910 $D=103
M2195 3230 WL_147 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=313400 $D=103
M2196 2933 WL_148 3232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=316310 $D=103
M2197 3234 WL_149 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=316800 $D=103
M2198 2933 WL_150 3236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=319710 $D=103
M2199 3238 WL_151 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=320200 $D=103
M2200 2933 WL_152 3240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=323110 $D=103
M2201 3242 WL_153 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=323600 $D=103
M2202 2933 WL_154 3244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=326510 $D=103
M2203 3246 WL_155 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=327000 $D=103
M2204 2933 WL_156 3248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=329910 $D=103
M2205 3250 WL_157 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=330400 $D=103
M2206 2933 WL_158 3252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=333310 $D=103
M2207 3254 WL_159 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=333800 $D=103
M2208 2933 WL_160 3256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=336710 $D=103
M2209 3258 WL_161 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=337200 $D=103
M2210 2933 WL_162 3260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=340110 $D=103
M2211 3262 WL_163 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=340600 $D=103
M2212 2933 WL_164 3264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=343510 $D=103
M2213 3266 WL_165 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=344000 $D=103
M2214 2933 WL_166 3268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=346910 $D=103
M2215 3270 WL_167 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=347400 $D=103
M2216 2933 WL_168 3272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=350310 $D=103
M2217 3274 WL_169 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=350800 $D=103
M2218 2933 WL_170 3276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=353710 $D=103
M2219 3278 WL_171 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=354200 $D=103
M2220 2933 WL_172 3280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=357110 $D=103
M2221 3282 WL_173 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=357600 $D=103
M2222 2933 WL_174 3284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=360510 $D=103
M2223 3286 WL_175 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=361000 $D=103
M2224 2933 WL_176 3288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=363910 $D=103
M2225 3290 WL_177 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=364400 $D=103
M2226 2933 WL_178 3292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=367310 $D=103
M2227 3294 WL_179 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=367800 $D=103
M2228 2933 WL_180 3296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=370710 $D=103
M2229 3298 WL_181 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=371200 $D=103
M2230 2933 WL_182 3300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=374110 $D=103
M2231 3302 WL_183 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=374600 $D=103
M2232 2933 WL_184 3304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=377510 $D=103
M2233 3306 WL_185 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=378000 $D=103
M2234 2933 WL_186 3308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=380910 $D=103
M2235 3310 WL_187 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=381400 $D=103
M2236 2933 WL_188 3312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=384310 $D=103
M2237 3314 WL_189 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=384800 $D=103
M2238 2933 WL_190 3316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=387710 $D=103
M2239 3318 WL_191 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=388200 $D=103
M2240 2933 WL_192 3320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=391110 $D=103
M2241 3322 WL_193 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=391600 $D=103
M2242 2933 WL_194 3324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=394510 $D=103
M2243 3326 WL_195 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=395000 $D=103
M2244 2933 WL_196 3328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=397910 $D=103
M2245 3330 WL_197 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=398400 $D=103
M2246 2933 WL_198 3332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=401310 $D=103
M2247 3334 WL_199 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=401800 $D=103
M2248 2933 WL_200 3336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=404710 $D=103
M2249 3338 WL_201 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=405200 $D=103
M2250 2933 WL_202 3340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=408110 $D=103
M2251 3342 WL_203 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=408600 $D=103
M2252 2933 WL_204 3344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=411510 $D=103
M2253 3346 WL_205 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=412000 $D=103
M2254 2933 WL_206 3348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=414910 $D=103
M2255 3350 WL_207 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=415400 $D=103
M2256 2933 WL_208 3352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=418310 $D=103
M2257 3354 WL_209 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=418800 $D=103
M2258 2933 WL_210 3356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=421710 $D=103
M2259 3358 WL_211 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=422200 $D=103
M2260 2933 WL_212 3360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=425110 $D=103
M2261 3362 WL_213 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=425600 $D=103
M2262 2933 WL_214 3364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=428510 $D=103
M2263 3366 WL_215 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=429000 $D=103
M2264 2933 WL_216 3368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=431910 $D=103
M2265 3370 WL_217 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=432400 $D=103
M2266 2933 WL_218 3372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=435310 $D=103
M2267 3374 WL_219 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=435800 $D=103
M2268 2933 WL_220 3376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=438710 $D=103
M2269 3378 WL_221 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=439200 $D=103
M2270 2933 WL_222 3380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=442110 $D=103
M2271 3382 WL_223 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=442600 $D=103
M2272 2933 WL_224 3384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=445510 $D=103
M2273 3386 WL_225 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=446000 $D=103
M2274 2933 WL_226 3388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=448910 $D=103
M2275 3390 WL_227 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=449400 $D=103
M2276 2933 WL_228 3392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=452310 $D=103
M2277 3394 WL_229 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=452800 $D=103
M2278 2933 WL_230 3396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=455710 $D=103
M2279 3398 WL_231 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=456200 $D=103
M2280 2933 WL_232 3400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=459110 $D=103
M2281 3402 WL_233 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=459600 $D=103
M2282 2933 WL_234 3404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=462510 $D=103
M2283 3406 WL_235 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=463000 $D=103
M2284 2933 WL_236 3408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=465910 $D=103
M2285 3410 WL_237 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=466400 $D=103
M2286 2933 WL_238 3412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=469310 $D=103
M2287 3414 WL_239 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=469800 $D=103
M2288 2933 WL_240 3416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=472710 $D=103
M2289 3418 WL_241 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=473200 $D=103
M2290 2933 WL_242 3420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=476110 $D=103
M2291 3422 WL_243 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=476600 $D=103
M2292 2933 WL_244 3424 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=479510 $D=103
M2293 3426 WL_245 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=480000 $D=103
M2294 2933 WL_246 3428 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=482910 $D=103
M2295 3430 WL_247 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=483400 $D=103
M2296 2933 WL_248 3432 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=486310 $D=103
M2297 3434 WL_249 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=486800 $D=103
M2298 2933 WL_250 3436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=489710 $D=103
M2299 3438 WL_251 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=490200 $D=103
M2300 2933 WL_252 3440 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=493110 $D=103
M2301 3442 WL_253 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=493600 $D=103
M2302 2933 WL_254 3444 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=496510 $D=103
M2303 3446 WL_255 2933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98150 $Y=497000 $D=103
M2304 3447 WL_0 3449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=64710 $D=103
M2305 3451 WL_1 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=65200 $D=103
M2306 3447 WL_2 3453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=68110 $D=103
M2307 3455 WL_3 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=68600 $D=103
M2308 3447 WL_4 3457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=71510 $D=103
M2309 3459 WL_5 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=72000 $D=103
M2310 3447 WL_6 3461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=74910 $D=103
M2311 3463 WL_7 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=75400 $D=103
M2312 3447 WL_8 3465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=78310 $D=103
M2313 3467 WL_9 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=78800 $D=103
M2314 3447 WL_10 3469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=81710 $D=103
M2315 3471 WL_11 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=82200 $D=103
M2316 3447 WL_12 3473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=85110 $D=103
M2317 3475 WL_13 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=85600 $D=103
M2318 3447 WL_14 3477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=88510 $D=103
M2319 3479 WL_15 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=89000 $D=103
M2320 3447 WL_16 3481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=91910 $D=103
M2321 3483 WL_17 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=92400 $D=103
M2322 3447 WL_18 3485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=95310 $D=103
M2323 3487 WL_19 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=95800 $D=103
M2324 3447 WL_20 3489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=98710 $D=103
M2325 3491 WL_21 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=99200 $D=103
M2326 3447 WL_22 3493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=102110 $D=103
M2327 3495 WL_23 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=102600 $D=103
M2328 3447 WL_24 3497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=105510 $D=103
M2329 3499 WL_25 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=106000 $D=103
M2330 3447 WL_26 3501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=108910 $D=103
M2331 3503 WL_27 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=109400 $D=103
M2332 3447 WL_28 3505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=112310 $D=103
M2333 3507 WL_29 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=112800 $D=103
M2334 3447 WL_30 3509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=115710 $D=103
M2335 3511 WL_31 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=116200 $D=103
M2336 3447 WL_32 3513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=119110 $D=103
M2337 3515 WL_33 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=119600 $D=103
M2338 3447 WL_34 3517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=122510 $D=103
M2339 3519 WL_35 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=123000 $D=103
M2340 3447 WL_36 3521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=125910 $D=103
M2341 3523 WL_37 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=126400 $D=103
M2342 3447 WL_38 3525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=129310 $D=103
M2343 3527 WL_39 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=129800 $D=103
M2344 3447 WL_40 3529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=132710 $D=103
M2345 3531 WL_41 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=133200 $D=103
M2346 3447 WL_42 3533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=136110 $D=103
M2347 3535 WL_43 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=136600 $D=103
M2348 3447 WL_44 3537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=139510 $D=103
M2349 3539 WL_45 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=140000 $D=103
M2350 3447 WL_46 3541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=142910 $D=103
M2351 3543 WL_47 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=143400 $D=103
M2352 3447 WL_48 3545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=146310 $D=103
M2353 3547 WL_49 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=146800 $D=103
M2354 3447 WL_50 3549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=149710 $D=103
M2355 3551 WL_51 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=150200 $D=103
M2356 3447 WL_52 3553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=153110 $D=103
M2357 3555 WL_53 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=153600 $D=103
M2358 3447 WL_54 3557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=156510 $D=103
M2359 3559 WL_55 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=157000 $D=103
M2360 3447 WL_56 3561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=159910 $D=103
M2361 3563 WL_57 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=160400 $D=103
M2362 3447 WL_58 3565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=163310 $D=103
M2363 3567 WL_59 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=163800 $D=103
M2364 3447 WL_60 3569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=166710 $D=103
M2365 3571 WL_61 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=167200 $D=103
M2366 3447 WL_62 3573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=170110 $D=103
M2367 3575 WL_63 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=170600 $D=103
M2368 3447 WL_64 3577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=173510 $D=103
M2369 3579 WL_65 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=174000 $D=103
M2370 3447 WL_66 3581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=176910 $D=103
M2371 3583 WL_67 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=177400 $D=103
M2372 3447 WL_68 3585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=180310 $D=103
M2373 3587 WL_69 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=180800 $D=103
M2374 3447 WL_70 3589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=183710 $D=103
M2375 3591 WL_71 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=184200 $D=103
M2376 3447 WL_72 3593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=187110 $D=103
M2377 3595 WL_73 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=187600 $D=103
M2378 3447 WL_74 3597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=190510 $D=103
M2379 3599 WL_75 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=191000 $D=103
M2380 3447 WL_76 3601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=193910 $D=103
M2381 3603 WL_77 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=194400 $D=103
M2382 3447 WL_78 3605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=197310 $D=103
M2383 3607 WL_79 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=197800 $D=103
M2384 3447 WL_80 3609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=200710 $D=103
M2385 3611 WL_81 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=201200 $D=103
M2386 3447 WL_82 3613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=204110 $D=103
M2387 3615 WL_83 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=204600 $D=103
M2388 3447 WL_84 3617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=207510 $D=103
M2389 3619 WL_85 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=208000 $D=103
M2390 3447 WL_86 3621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=210910 $D=103
M2391 3623 WL_87 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=211400 $D=103
M2392 3447 WL_88 3625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=214310 $D=103
M2393 3627 WL_89 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=214800 $D=103
M2394 3447 WL_90 3629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=217710 $D=103
M2395 3631 WL_91 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=218200 $D=103
M2396 3447 WL_92 3633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=221110 $D=103
M2397 3635 WL_93 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=221600 $D=103
M2398 3447 WL_94 3637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=224510 $D=103
M2399 3639 WL_95 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=225000 $D=103
M2400 3447 WL_96 3641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=227910 $D=103
M2401 3643 WL_97 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=228400 $D=103
M2402 3447 WL_98 3645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=231310 $D=103
M2403 3647 WL_99 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=231800 $D=103
M2404 3447 WL_100 3649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=234710 $D=103
M2405 3651 WL_101 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=235200 $D=103
M2406 3447 WL_102 3653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=238110 $D=103
M2407 3655 WL_103 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=238600 $D=103
M2408 3447 WL_104 3657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=241510 $D=103
M2409 3659 WL_105 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=242000 $D=103
M2410 3447 WL_106 3661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=244910 $D=103
M2411 3663 WL_107 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=245400 $D=103
M2412 3447 WL_108 3665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=248310 $D=103
M2413 3667 WL_109 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=248800 $D=103
M2414 3447 WL_110 3669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=251710 $D=103
M2415 3671 WL_111 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=252200 $D=103
M2416 3447 WL_112 3673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=255110 $D=103
M2417 3675 WL_113 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=255600 $D=103
M2418 3447 WL_114 3677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=258510 $D=103
M2419 3679 WL_115 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=259000 $D=103
M2420 3447 WL_116 3681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=261910 $D=103
M2421 3683 WL_117 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=262400 $D=103
M2422 3447 WL_118 3685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=265310 $D=103
M2423 3687 WL_119 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=265800 $D=103
M2424 3447 WL_120 3689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=268710 $D=103
M2425 3691 WL_121 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=269200 $D=103
M2426 3447 WL_122 3693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=272110 $D=103
M2427 3695 WL_123 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=272600 $D=103
M2428 3447 WL_124 3697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=275510 $D=103
M2429 3699 WL_125 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=276000 $D=103
M2430 3447 WL_126 3701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=278910 $D=103
M2431 3703 WL_127 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=279400 $D=103
M2432 3447 WL_128 3705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=282310 $D=103
M2433 3707 WL_129 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=282800 $D=103
M2434 3447 WL_130 3709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=285710 $D=103
M2435 3711 WL_131 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=286200 $D=103
M2436 3447 WL_132 3713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=289110 $D=103
M2437 3715 WL_133 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=289600 $D=103
M2438 3447 WL_134 3717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=292510 $D=103
M2439 3719 WL_135 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=293000 $D=103
M2440 3447 WL_136 3721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=295910 $D=103
M2441 3723 WL_137 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=296400 $D=103
M2442 3447 WL_138 3725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=299310 $D=103
M2443 3727 WL_139 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=299800 $D=103
M2444 3447 WL_140 3729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=302710 $D=103
M2445 3731 WL_141 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=303200 $D=103
M2446 3447 WL_142 3733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=306110 $D=103
M2447 3735 WL_143 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=306600 $D=103
M2448 3447 WL_144 3737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=309510 $D=103
M2449 3739 WL_145 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=310000 $D=103
M2450 3447 WL_146 3741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=312910 $D=103
M2451 3743 WL_147 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=313400 $D=103
M2452 3447 WL_148 3745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=316310 $D=103
M2453 3747 WL_149 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=316800 $D=103
M2454 3447 WL_150 3749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=319710 $D=103
M2455 3751 WL_151 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=320200 $D=103
M2456 3447 WL_152 3753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=323110 $D=103
M2457 3755 WL_153 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=323600 $D=103
M2458 3447 WL_154 3757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=326510 $D=103
M2459 3759 WL_155 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=327000 $D=103
M2460 3447 WL_156 3761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=329910 $D=103
M2461 3763 WL_157 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=330400 $D=103
M2462 3447 WL_158 3765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=333310 $D=103
M2463 3767 WL_159 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=333800 $D=103
M2464 3447 WL_160 3769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=336710 $D=103
M2465 3771 WL_161 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=337200 $D=103
M2466 3447 WL_162 3773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=340110 $D=103
M2467 3775 WL_163 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=340600 $D=103
M2468 3447 WL_164 3777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=343510 $D=103
M2469 3779 WL_165 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=344000 $D=103
M2470 3447 WL_166 3781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=346910 $D=103
M2471 3783 WL_167 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=347400 $D=103
M2472 3447 WL_168 3785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=350310 $D=103
M2473 3787 WL_169 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=350800 $D=103
M2474 3447 WL_170 3789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=353710 $D=103
M2475 3791 WL_171 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=354200 $D=103
M2476 3447 WL_172 3793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=357110 $D=103
M2477 3795 WL_173 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=357600 $D=103
M2478 3447 WL_174 3797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=360510 $D=103
M2479 3799 WL_175 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=361000 $D=103
M2480 3447 WL_176 3801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=363910 $D=103
M2481 3803 WL_177 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=364400 $D=103
M2482 3447 WL_178 3805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=367310 $D=103
M2483 3807 WL_179 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=367800 $D=103
M2484 3447 WL_180 3809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=370710 $D=103
M2485 3811 WL_181 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=371200 $D=103
M2486 3447 WL_182 3813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=374110 $D=103
M2487 3815 WL_183 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=374600 $D=103
M2488 3447 WL_184 3817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=377510 $D=103
M2489 3819 WL_185 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=378000 $D=103
M2490 3447 WL_186 3821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=380910 $D=103
M2491 3823 WL_187 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=381400 $D=103
M2492 3447 WL_188 3825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=384310 $D=103
M2493 3827 WL_189 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=384800 $D=103
M2494 3447 WL_190 3829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=387710 $D=103
M2495 3831 WL_191 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=388200 $D=103
M2496 3447 WL_192 3833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=391110 $D=103
M2497 3835 WL_193 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=391600 $D=103
M2498 3447 WL_194 3837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=394510 $D=103
M2499 3839 WL_195 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=395000 $D=103
M2500 3447 WL_196 3841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=397910 $D=103
M2501 3843 WL_197 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=398400 $D=103
M2502 3447 WL_198 3845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=401310 $D=103
M2503 3847 WL_199 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=401800 $D=103
M2504 3447 WL_200 3849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=404710 $D=103
M2505 3851 WL_201 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=405200 $D=103
M2506 3447 WL_202 3853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=408110 $D=103
M2507 3855 WL_203 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=408600 $D=103
M2508 3447 WL_204 3857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=411510 $D=103
M2509 3859 WL_205 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=412000 $D=103
M2510 3447 WL_206 3861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=414910 $D=103
M2511 3863 WL_207 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=415400 $D=103
M2512 3447 WL_208 3865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=418310 $D=103
M2513 3867 WL_209 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=418800 $D=103
M2514 3447 WL_210 3869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=421710 $D=103
M2515 3871 WL_211 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=422200 $D=103
M2516 3447 WL_212 3873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=425110 $D=103
M2517 3875 WL_213 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=425600 $D=103
M2518 3447 WL_214 3877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=428510 $D=103
M2519 3879 WL_215 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=429000 $D=103
M2520 3447 WL_216 3881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=431910 $D=103
M2521 3883 WL_217 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=432400 $D=103
M2522 3447 WL_218 3885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=435310 $D=103
M2523 3887 WL_219 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=435800 $D=103
M2524 3447 WL_220 3889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=438710 $D=103
M2525 3891 WL_221 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=439200 $D=103
M2526 3447 WL_222 3893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=442110 $D=103
M2527 3895 WL_223 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=442600 $D=103
M2528 3447 WL_224 3897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=445510 $D=103
M2529 3899 WL_225 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=446000 $D=103
M2530 3447 WL_226 3901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=448910 $D=103
M2531 3903 WL_227 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=449400 $D=103
M2532 3447 WL_228 3905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=452310 $D=103
M2533 3907 WL_229 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=452800 $D=103
M2534 3447 WL_230 3909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=455710 $D=103
M2535 3911 WL_231 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=456200 $D=103
M2536 3447 WL_232 3913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=459110 $D=103
M2537 3915 WL_233 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=459600 $D=103
M2538 3447 WL_234 3917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=462510 $D=103
M2539 3919 WL_235 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=463000 $D=103
M2540 3447 WL_236 3921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=465910 $D=103
M2541 3923 WL_237 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=466400 $D=103
M2542 3447 WL_238 3925 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=469310 $D=103
M2543 3927 WL_239 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=469800 $D=103
M2544 3447 WL_240 3929 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=472710 $D=103
M2545 3931 WL_241 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=473200 $D=103
M2546 3447 WL_242 3933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=476110 $D=103
M2547 3935 WL_243 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=476600 $D=103
M2548 3447 WL_244 3937 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=479510 $D=103
M2549 3939 WL_245 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=480000 $D=103
M2550 3447 WL_246 3941 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=482910 $D=103
M2551 3943 WL_247 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=483400 $D=103
M2552 3447 WL_248 3945 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=486310 $D=103
M2553 3947 WL_249 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=486800 $D=103
M2554 3447 WL_250 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=489710 $D=103
M2555 3951 WL_251 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=490200 $D=103
M2556 3447 WL_252 3953 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=493110 $D=103
M2557 3955 WL_253 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=493600 $D=103
M2558 3447 WL_254 3957 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=496510 $D=103
M2559 3959 WL_255 3447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98490 $Y=497000 $D=103
M2560 3448 WL_0 3450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=64710 $D=103
M2561 3452 WL_1 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=65200 $D=103
M2562 3448 WL_2 3454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=68110 $D=103
M2563 3456 WL_3 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=68600 $D=103
M2564 3448 WL_4 3458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=71510 $D=103
M2565 3460 WL_5 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=72000 $D=103
M2566 3448 WL_6 3462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=74910 $D=103
M2567 3464 WL_7 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=75400 $D=103
M2568 3448 WL_8 3466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=78310 $D=103
M2569 3468 WL_9 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=78800 $D=103
M2570 3448 WL_10 3470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=81710 $D=103
M2571 3472 WL_11 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=82200 $D=103
M2572 3448 WL_12 3474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=85110 $D=103
M2573 3476 WL_13 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=85600 $D=103
M2574 3448 WL_14 3478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=88510 $D=103
M2575 3480 WL_15 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=89000 $D=103
M2576 3448 WL_16 3482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=91910 $D=103
M2577 3484 WL_17 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=92400 $D=103
M2578 3448 WL_18 3486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=95310 $D=103
M2579 3488 WL_19 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=95800 $D=103
M2580 3448 WL_20 3490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=98710 $D=103
M2581 3492 WL_21 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=99200 $D=103
M2582 3448 WL_22 3494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=102110 $D=103
M2583 3496 WL_23 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=102600 $D=103
M2584 3448 WL_24 3498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=105510 $D=103
M2585 3500 WL_25 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=106000 $D=103
M2586 3448 WL_26 3502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=108910 $D=103
M2587 3504 WL_27 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=109400 $D=103
M2588 3448 WL_28 3506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=112310 $D=103
M2589 3508 WL_29 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=112800 $D=103
M2590 3448 WL_30 3510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=115710 $D=103
M2591 3512 WL_31 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=116200 $D=103
M2592 3448 WL_32 3514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=119110 $D=103
M2593 3516 WL_33 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=119600 $D=103
M2594 3448 WL_34 3518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=122510 $D=103
M2595 3520 WL_35 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=123000 $D=103
M2596 3448 WL_36 3522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=125910 $D=103
M2597 3524 WL_37 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=126400 $D=103
M2598 3448 WL_38 3526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=129310 $D=103
M2599 3528 WL_39 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=129800 $D=103
M2600 3448 WL_40 3530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=132710 $D=103
M2601 3532 WL_41 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=133200 $D=103
M2602 3448 WL_42 3534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=136110 $D=103
M2603 3536 WL_43 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=136600 $D=103
M2604 3448 WL_44 3538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=139510 $D=103
M2605 3540 WL_45 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=140000 $D=103
M2606 3448 WL_46 3542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=142910 $D=103
M2607 3544 WL_47 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=143400 $D=103
M2608 3448 WL_48 3546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=146310 $D=103
M2609 3548 WL_49 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=146800 $D=103
M2610 3448 WL_50 3550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=149710 $D=103
M2611 3552 WL_51 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=150200 $D=103
M2612 3448 WL_52 3554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=153110 $D=103
M2613 3556 WL_53 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=153600 $D=103
M2614 3448 WL_54 3558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=156510 $D=103
M2615 3560 WL_55 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=157000 $D=103
M2616 3448 WL_56 3562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=159910 $D=103
M2617 3564 WL_57 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=160400 $D=103
M2618 3448 WL_58 3566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=163310 $D=103
M2619 3568 WL_59 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=163800 $D=103
M2620 3448 WL_60 3570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=166710 $D=103
M2621 3572 WL_61 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=167200 $D=103
M2622 3448 WL_62 3574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=170110 $D=103
M2623 3576 WL_63 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=170600 $D=103
M2624 3448 WL_64 3578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=173510 $D=103
M2625 3580 WL_65 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=174000 $D=103
M2626 3448 WL_66 3582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=176910 $D=103
M2627 3584 WL_67 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=177400 $D=103
M2628 3448 WL_68 3586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=180310 $D=103
M2629 3588 WL_69 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=180800 $D=103
M2630 3448 WL_70 3590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=183710 $D=103
M2631 3592 WL_71 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=184200 $D=103
M2632 3448 WL_72 3594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=187110 $D=103
M2633 3596 WL_73 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=187600 $D=103
M2634 3448 WL_74 3598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=190510 $D=103
M2635 3600 WL_75 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=191000 $D=103
M2636 3448 WL_76 3602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=193910 $D=103
M2637 3604 WL_77 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=194400 $D=103
M2638 3448 WL_78 3606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=197310 $D=103
M2639 3608 WL_79 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=197800 $D=103
M2640 3448 WL_80 3610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=200710 $D=103
M2641 3612 WL_81 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=201200 $D=103
M2642 3448 WL_82 3614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=204110 $D=103
M2643 3616 WL_83 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=204600 $D=103
M2644 3448 WL_84 3618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=207510 $D=103
M2645 3620 WL_85 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=208000 $D=103
M2646 3448 WL_86 3622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=210910 $D=103
M2647 3624 WL_87 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=211400 $D=103
M2648 3448 WL_88 3626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=214310 $D=103
M2649 3628 WL_89 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=214800 $D=103
M2650 3448 WL_90 3630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=217710 $D=103
M2651 3632 WL_91 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=218200 $D=103
M2652 3448 WL_92 3634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=221110 $D=103
M2653 3636 WL_93 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=221600 $D=103
M2654 3448 WL_94 3638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=224510 $D=103
M2655 3640 WL_95 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=225000 $D=103
M2656 3448 WL_96 3642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=227910 $D=103
M2657 3644 WL_97 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=228400 $D=103
M2658 3448 WL_98 3646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=231310 $D=103
M2659 3648 WL_99 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=231800 $D=103
M2660 3448 WL_100 3650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=234710 $D=103
M2661 3652 WL_101 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=235200 $D=103
M2662 3448 WL_102 3654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=238110 $D=103
M2663 3656 WL_103 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=238600 $D=103
M2664 3448 WL_104 3658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=241510 $D=103
M2665 3660 WL_105 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=242000 $D=103
M2666 3448 WL_106 3662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=244910 $D=103
M2667 3664 WL_107 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=245400 $D=103
M2668 3448 WL_108 3666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=248310 $D=103
M2669 3668 WL_109 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=248800 $D=103
M2670 3448 WL_110 3670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=251710 $D=103
M2671 3672 WL_111 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=252200 $D=103
M2672 3448 WL_112 3674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=255110 $D=103
M2673 3676 WL_113 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=255600 $D=103
M2674 3448 WL_114 3678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=258510 $D=103
M2675 3680 WL_115 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=259000 $D=103
M2676 3448 WL_116 3682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=261910 $D=103
M2677 3684 WL_117 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=262400 $D=103
M2678 3448 WL_118 3686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=265310 $D=103
M2679 3688 WL_119 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=265800 $D=103
M2680 3448 WL_120 3690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=268710 $D=103
M2681 3692 WL_121 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=269200 $D=103
M2682 3448 WL_122 3694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=272110 $D=103
M2683 3696 WL_123 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=272600 $D=103
M2684 3448 WL_124 3698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=275510 $D=103
M2685 3700 WL_125 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=276000 $D=103
M2686 3448 WL_126 3702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=278910 $D=103
M2687 3704 WL_127 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=279400 $D=103
M2688 3448 WL_128 3706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=282310 $D=103
M2689 3708 WL_129 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=282800 $D=103
M2690 3448 WL_130 3710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=285710 $D=103
M2691 3712 WL_131 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=286200 $D=103
M2692 3448 WL_132 3714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=289110 $D=103
M2693 3716 WL_133 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=289600 $D=103
M2694 3448 WL_134 3718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=292510 $D=103
M2695 3720 WL_135 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=293000 $D=103
M2696 3448 WL_136 3722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=295910 $D=103
M2697 3724 WL_137 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=296400 $D=103
M2698 3448 WL_138 3726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=299310 $D=103
M2699 3728 WL_139 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=299800 $D=103
M2700 3448 WL_140 3730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=302710 $D=103
M2701 3732 WL_141 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=303200 $D=103
M2702 3448 WL_142 3734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=306110 $D=103
M2703 3736 WL_143 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=306600 $D=103
M2704 3448 WL_144 3738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=309510 $D=103
M2705 3740 WL_145 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=310000 $D=103
M2706 3448 WL_146 3742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=312910 $D=103
M2707 3744 WL_147 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=313400 $D=103
M2708 3448 WL_148 3746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=316310 $D=103
M2709 3748 WL_149 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=316800 $D=103
M2710 3448 WL_150 3750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=319710 $D=103
M2711 3752 WL_151 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=320200 $D=103
M2712 3448 WL_152 3754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=323110 $D=103
M2713 3756 WL_153 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=323600 $D=103
M2714 3448 WL_154 3758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=326510 $D=103
M2715 3760 WL_155 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=327000 $D=103
M2716 3448 WL_156 3762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=329910 $D=103
M2717 3764 WL_157 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=330400 $D=103
M2718 3448 WL_158 3766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=333310 $D=103
M2719 3768 WL_159 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=333800 $D=103
M2720 3448 WL_160 3770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=336710 $D=103
M2721 3772 WL_161 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=337200 $D=103
M2722 3448 WL_162 3774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=340110 $D=103
M2723 3776 WL_163 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=340600 $D=103
M2724 3448 WL_164 3778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=343510 $D=103
M2725 3780 WL_165 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=344000 $D=103
M2726 3448 WL_166 3782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=346910 $D=103
M2727 3784 WL_167 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=347400 $D=103
M2728 3448 WL_168 3786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=350310 $D=103
M2729 3788 WL_169 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=350800 $D=103
M2730 3448 WL_170 3790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=353710 $D=103
M2731 3792 WL_171 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=354200 $D=103
M2732 3448 WL_172 3794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=357110 $D=103
M2733 3796 WL_173 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=357600 $D=103
M2734 3448 WL_174 3798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=360510 $D=103
M2735 3800 WL_175 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=361000 $D=103
M2736 3448 WL_176 3802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=363910 $D=103
M2737 3804 WL_177 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=364400 $D=103
M2738 3448 WL_178 3806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=367310 $D=103
M2739 3808 WL_179 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=367800 $D=103
M2740 3448 WL_180 3810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=370710 $D=103
M2741 3812 WL_181 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=371200 $D=103
M2742 3448 WL_182 3814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=374110 $D=103
M2743 3816 WL_183 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=374600 $D=103
M2744 3448 WL_184 3818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=377510 $D=103
M2745 3820 WL_185 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=378000 $D=103
M2746 3448 WL_186 3822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=380910 $D=103
M2747 3824 WL_187 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=381400 $D=103
M2748 3448 WL_188 3826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=384310 $D=103
M2749 3828 WL_189 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=384800 $D=103
M2750 3448 WL_190 3830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=387710 $D=103
M2751 3832 WL_191 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=388200 $D=103
M2752 3448 WL_192 3834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=391110 $D=103
M2753 3836 WL_193 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=391600 $D=103
M2754 3448 WL_194 3838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=394510 $D=103
M2755 3840 WL_195 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=395000 $D=103
M2756 3448 WL_196 3842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=397910 $D=103
M2757 3844 WL_197 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=398400 $D=103
M2758 3448 WL_198 3846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=401310 $D=103
M2759 3848 WL_199 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=401800 $D=103
M2760 3448 WL_200 3850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=404710 $D=103
M2761 3852 WL_201 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=405200 $D=103
M2762 3448 WL_202 3854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=408110 $D=103
M2763 3856 WL_203 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=408600 $D=103
M2764 3448 WL_204 3858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=411510 $D=103
M2765 3860 WL_205 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=412000 $D=103
M2766 3448 WL_206 3862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=414910 $D=103
M2767 3864 WL_207 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=415400 $D=103
M2768 3448 WL_208 3866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=418310 $D=103
M2769 3868 WL_209 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=418800 $D=103
M2770 3448 WL_210 3870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=421710 $D=103
M2771 3872 WL_211 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=422200 $D=103
M2772 3448 WL_212 3874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=425110 $D=103
M2773 3876 WL_213 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=425600 $D=103
M2774 3448 WL_214 3878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=428510 $D=103
M2775 3880 WL_215 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=429000 $D=103
M2776 3448 WL_216 3882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=431910 $D=103
M2777 3884 WL_217 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=432400 $D=103
M2778 3448 WL_218 3886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=435310 $D=103
M2779 3888 WL_219 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=435800 $D=103
M2780 3448 WL_220 3890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=438710 $D=103
M2781 3892 WL_221 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=439200 $D=103
M2782 3448 WL_222 3894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=442110 $D=103
M2783 3896 WL_223 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=442600 $D=103
M2784 3448 WL_224 3898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=445510 $D=103
M2785 3900 WL_225 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=446000 $D=103
M2786 3448 WL_226 3902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=448910 $D=103
M2787 3904 WL_227 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=449400 $D=103
M2788 3448 WL_228 3906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=452310 $D=103
M2789 3908 WL_229 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=452800 $D=103
M2790 3448 WL_230 3910 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=455710 $D=103
M2791 3912 WL_231 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=456200 $D=103
M2792 3448 WL_232 3914 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=459110 $D=103
M2793 3916 WL_233 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=459600 $D=103
M2794 3448 WL_234 3918 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=462510 $D=103
M2795 3920 WL_235 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=463000 $D=103
M2796 3448 WL_236 3922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=465910 $D=103
M2797 3924 WL_237 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=466400 $D=103
M2798 3448 WL_238 3926 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=469310 $D=103
M2799 3928 WL_239 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=469800 $D=103
M2800 3448 WL_240 3930 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=472710 $D=103
M2801 3932 WL_241 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=473200 $D=103
M2802 3448 WL_242 3934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=476110 $D=103
M2803 3936 WL_243 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=476600 $D=103
M2804 3448 WL_244 3938 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=479510 $D=103
M2805 3940 WL_245 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=480000 $D=103
M2806 3448 WL_246 3942 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=482910 $D=103
M2807 3944 WL_247 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=483400 $D=103
M2808 3448 WL_248 3946 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=486310 $D=103
M2809 3948 WL_249 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=486800 $D=103
M2810 3448 WL_250 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=489710 $D=103
M2811 3952 WL_251 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=490200 $D=103
M2812 3448 WL_252 3954 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=493110 $D=103
M2813 3956 WL_253 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=493600 $D=103
M2814 3448 WL_254 3958 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=496510 $D=103
M2815 3960 WL_255 3448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117350 $Y=497000 $D=103
M2816 3962 WL_0 3963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=64710 $D=103
M2817 3965 WL_1 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=65200 $D=103
M2818 3962 WL_2 3967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=68110 $D=103
M2819 3969 WL_3 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=68600 $D=103
M2820 3962 WL_4 3971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=71510 $D=103
M2821 3973 WL_5 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=72000 $D=103
M2822 3962 WL_6 3975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=74910 $D=103
M2823 3977 WL_7 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=75400 $D=103
M2824 3962 WL_8 3979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=78310 $D=103
M2825 3981 WL_9 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=78800 $D=103
M2826 3962 WL_10 3983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=81710 $D=103
M2827 3985 WL_11 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=82200 $D=103
M2828 3962 WL_12 3987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=85110 $D=103
M2829 3989 WL_13 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=85600 $D=103
M2830 3962 WL_14 3991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=88510 $D=103
M2831 3993 WL_15 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=89000 $D=103
M2832 3962 WL_16 3995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=91910 $D=103
M2833 3997 WL_17 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=92400 $D=103
M2834 3962 WL_18 3999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=95310 $D=103
M2835 4001 WL_19 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=95800 $D=103
M2836 3962 WL_20 4003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=98710 $D=103
M2837 4005 WL_21 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=99200 $D=103
M2838 3962 WL_22 4007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=102110 $D=103
M2839 4009 WL_23 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=102600 $D=103
M2840 3962 WL_24 4011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=105510 $D=103
M2841 4013 WL_25 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=106000 $D=103
M2842 3962 WL_26 4015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=108910 $D=103
M2843 4017 WL_27 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=109400 $D=103
M2844 3962 WL_28 4019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=112310 $D=103
M2845 4021 WL_29 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=112800 $D=103
M2846 3962 WL_30 4023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=115710 $D=103
M2847 4025 WL_31 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=116200 $D=103
M2848 3962 WL_32 4027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=119110 $D=103
M2849 4029 WL_33 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=119600 $D=103
M2850 3962 WL_34 4031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=122510 $D=103
M2851 4033 WL_35 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=123000 $D=103
M2852 3962 WL_36 4035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=125910 $D=103
M2853 4037 WL_37 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=126400 $D=103
M2854 3962 WL_38 4039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=129310 $D=103
M2855 4041 WL_39 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=129800 $D=103
M2856 3962 WL_40 4043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=132710 $D=103
M2857 4045 WL_41 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=133200 $D=103
M2858 3962 WL_42 4047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=136110 $D=103
M2859 4049 WL_43 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=136600 $D=103
M2860 3962 WL_44 4051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=139510 $D=103
M2861 4053 WL_45 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=140000 $D=103
M2862 3962 WL_46 4055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=142910 $D=103
M2863 4057 WL_47 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=143400 $D=103
M2864 3962 WL_48 4059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=146310 $D=103
M2865 4061 WL_49 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=146800 $D=103
M2866 3962 WL_50 4063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=149710 $D=103
M2867 4065 WL_51 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=150200 $D=103
M2868 3962 WL_52 4067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=153110 $D=103
M2869 4069 WL_53 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=153600 $D=103
M2870 3962 WL_54 4071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=156510 $D=103
M2871 4073 WL_55 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=157000 $D=103
M2872 3962 WL_56 4075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=159910 $D=103
M2873 4077 WL_57 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=160400 $D=103
M2874 3962 WL_58 4079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=163310 $D=103
M2875 4081 WL_59 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=163800 $D=103
M2876 3962 WL_60 4083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=166710 $D=103
M2877 4085 WL_61 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=167200 $D=103
M2878 3962 WL_62 4087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=170110 $D=103
M2879 4089 WL_63 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=170600 $D=103
M2880 3962 WL_64 4091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=173510 $D=103
M2881 4093 WL_65 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=174000 $D=103
M2882 3962 WL_66 4095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=176910 $D=103
M2883 4097 WL_67 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=177400 $D=103
M2884 3962 WL_68 4099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=180310 $D=103
M2885 4101 WL_69 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=180800 $D=103
M2886 3962 WL_70 4103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=183710 $D=103
M2887 4105 WL_71 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=184200 $D=103
M2888 3962 WL_72 4107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=187110 $D=103
M2889 4109 WL_73 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=187600 $D=103
M2890 3962 WL_74 4111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=190510 $D=103
M2891 4113 WL_75 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=191000 $D=103
M2892 3962 WL_76 4115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=193910 $D=103
M2893 4117 WL_77 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=194400 $D=103
M2894 3962 WL_78 4119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=197310 $D=103
M2895 4121 WL_79 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=197800 $D=103
M2896 3962 WL_80 4123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=200710 $D=103
M2897 4125 WL_81 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=201200 $D=103
M2898 3962 WL_82 4127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=204110 $D=103
M2899 4129 WL_83 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=204600 $D=103
M2900 3962 WL_84 4131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=207510 $D=103
M2901 4133 WL_85 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=208000 $D=103
M2902 3962 WL_86 4135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=210910 $D=103
M2903 4137 WL_87 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=211400 $D=103
M2904 3962 WL_88 4139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=214310 $D=103
M2905 4141 WL_89 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=214800 $D=103
M2906 3962 WL_90 4143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=217710 $D=103
M2907 4145 WL_91 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=218200 $D=103
M2908 3962 WL_92 4147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=221110 $D=103
M2909 4149 WL_93 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=221600 $D=103
M2910 3962 WL_94 4151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=224510 $D=103
M2911 4153 WL_95 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=225000 $D=103
M2912 3962 WL_96 4155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=227910 $D=103
M2913 4157 WL_97 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=228400 $D=103
M2914 3962 WL_98 4159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=231310 $D=103
M2915 4161 WL_99 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=231800 $D=103
M2916 3962 WL_100 4163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=234710 $D=103
M2917 4165 WL_101 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=235200 $D=103
M2918 3962 WL_102 4167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=238110 $D=103
M2919 4169 WL_103 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=238600 $D=103
M2920 3962 WL_104 4171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=241510 $D=103
M2921 4173 WL_105 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=242000 $D=103
M2922 3962 WL_106 4175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=244910 $D=103
M2923 4177 WL_107 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=245400 $D=103
M2924 3962 WL_108 4179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=248310 $D=103
M2925 4181 WL_109 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=248800 $D=103
M2926 3962 WL_110 4183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=251710 $D=103
M2927 4185 WL_111 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=252200 $D=103
M2928 3962 WL_112 4187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=255110 $D=103
M2929 4189 WL_113 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=255600 $D=103
M2930 3962 WL_114 4191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=258510 $D=103
M2931 4193 WL_115 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=259000 $D=103
M2932 3962 WL_116 4195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=261910 $D=103
M2933 4197 WL_117 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=262400 $D=103
M2934 3962 WL_118 4199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=265310 $D=103
M2935 4201 WL_119 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=265800 $D=103
M2936 3962 WL_120 4203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=268710 $D=103
M2937 4205 WL_121 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=269200 $D=103
M2938 3962 WL_122 4207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=272110 $D=103
M2939 4209 WL_123 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=272600 $D=103
M2940 3962 WL_124 4211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=275510 $D=103
M2941 4213 WL_125 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=276000 $D=103
M2942 3962 WL_126 4215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=278910 $D=103
M2943 4217 WL_127 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=279400 $D=103
M2944 3962 WL_128 4219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=282310 $D=103
M2945 4221 WL_129 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=282800 $D=103
M2946 3962 WL_130 4223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=285710 $D=103
M2947 4225 WL_131 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=286200 $D=103
M2948 3962 WL_132 4227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=289110 $D=103
M2949 4229 WL_133 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=289600 $D=103
M2950 3962 WL_134 4231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=292510 $D=103
M2951 4233 WL_135 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=293000 $D=103
M2952 3962 WL_136 4235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=295910 $D=103
M2953 4237 WL_137 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=296400 $D=103
M2954 3962 WL_138 4239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=299310 $D=103
M2955 4241 WL_139 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=299800 $D=103
M2956 3962 WL_140 4243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=302710 $D=103
M2957 4245 WL_141 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=303200 $D=103
M2958 3962 WL_142 4247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=306110 $D=103
M2959 4249 WL_143 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=306600 $D=103
M2960 3962 WL_144 4251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=309510 $D=103
M2961 4253 WL_145 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=310000 $D=103
M2962 3962 WL_146 4255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=312910 $D=103
M2963 4257 WL_147 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=313400 $D=103
M2964 3962 WL_148 4259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=316310 $D=103
M2965 4261 WL_149 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=316800 $D=103
M2966 3962 WL_150 4263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=319710 $D=103
M2967 4265 WL_151 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=320200 $D=103
M2968 3962 WL_152 4267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=323110 $D=103
M2969 4269 WL_153 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=323600 $D=103
M2970 3962 WL_154 4271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=326510 $D=103
M2971 4273 WL_155 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=327000 $D=103
M2972 3962 WL_156 4275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=329910 $D=103
M2973 4277 WL_157 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=330400 $D=103
M2974 3962 WL_158 4279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=333310 $D=103
M2975 4281 WL_159 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=333800 $D=103
M2976 3962 WL_160 4283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=336710 $D=103
M2977 4285 WL_161 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=337200 $D=103
M2978 3962 WL_162 4287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=340110 $D=103
M2979 4289 WL_163 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=340600 $D=103
M2980 3962 WL_164 4291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=343510 $D=103
M2981 4293 WL_165 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=344000 $D=103
M2982 3962 WL_166 4295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=346910 $D=103
M2983 4297 WL_167 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=347400 $D=103
M2984 3962 WL_168 4299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=350310 $D=103
M2985 4301 WL_169 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=350800 $D=103
M2986 3962 WL_170 4303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=353710 $D=103
M2987 4305 WL_171 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=354200 $D=103
M2988 3962 WL_172 4307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=357110 $D=103
M2989 4309 WL_173 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=357600 $D=103
M2990 3962 WL_174 4311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=360510 $D=103
M2991 4313 WL_175 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=361000 $D=103
M2992 3962 WL_176 4315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=363910 $D=103
M2993 4317 WL_177 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=364400 $D=103
M2994 3962 WL_178 4319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=367310 $D=103
M2995 4321 WL_179 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=367800 $D=103
M2996 3962 WL_180 4323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=370710 $D=103
M2997 4325 WL_181 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=371200 $D=103
M2998 3962 WL_182 4327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=374110 $D=103
M2999 4329 WL_183 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=374600 $D=103
M3000 3962 WL_184 4331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=377510 $D=103
M3001 4333 WL_185 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=378000 $D=103
M3002 3962 WL_186 4335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=380910 $D=103
M3003 4337 WL_187 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=381400 $D=103
M3004 3962 WL_188 4339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=384310 $D=103
M3005 4341 WL_189 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=384800 $D=103
M3006 3962 WL_190 4343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=387710 $D=103
M3007 4345 WL_191 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=388200 $D=103
M3008 3962 WL_192 4347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=391110 $D=103
M3009 4349 WL_193 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=391600 $D=103
M3010 3962 WL_194 4351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=394510 $D=103
M3011 4353 WL_195 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=395000 $D=103
M3012 3962 WL_196 4355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=397910 $D=103
M3013 4357 WL_197 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=398400 $D=103
M3014 3962 WL_198 4359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=401310 $D=103
M3015 4361 WL_199 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=401800 $D=103
M3016 3962 WL_200 4363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=404710 $D=103
M3017 4365 WL_201 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=405200 $D=103
M3018 3962 WL_202 4367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=408110 $D=103
M3019 4369 WL_203 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=408600 $D=103
M3020 3962 WL_204 4371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=411510 $D=103
M3021 4373 WL_205 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=412000 $D=103
M3022 3962 WL_206 4375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=414910 $D=103
M3023 4377 WL_207 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=415400 $D=103
M3024 3962 WL_208 4379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=418310 $D=103
M3025 4381 WL_209 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=418800 $D=103
M3026 3962 WL_210 4383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=421710 $D=103
M3027 4385 WL_211 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=422200 $D=103
M3028 3962 WL_212 4387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=425110 $D=103
M3029 4389 WL_213 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=425600 $D=103
M3030 3962 WL_214 4391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=428510 $D=103
M3031 4393 WL_215 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=429000 $D=103
M3032 3962 WL_216 4395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=431910 $D=103
M3033 4397 WL_217 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=432400 $D=103
M3034 3962 WL_218 4399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=435310 $D=103
M3035 4401 WL_219 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=435800 $D=103
M3036 3962 WL_220 4403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=438710 $D=103
M3037 4405 WL_221 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=439200 $D=103
M3038 3962 WL_222 4407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=442110 $D=103
M3039 4409 WL_223 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=442600 $D=103
M3040 3962 WL_224 4411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=445510 $D=103
M3041 4413 WL_225 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=446000 $D=103
M3042 3962 WL_226 4415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=448910 $D=103
M3043 4417 WL_227 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=449400 $D=103
M3044 3962 WL_228 4419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=452310 $D=103
M3045 4421 WL_229 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=452800 $D=103
M3046 3962 WL_230 4423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=455710 $D=103
M3047 4425 WL_231 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=456200 $D=103
M3048 3962 WL_232 4427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=459110 $D=103
M3049 4429 WL_233 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=459600 $D=103
M3050 3962 WL_234 4431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=462510 $D=103
M3051 4433 WL_235 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=463000 $D=103
M3052 3962 WL_236 4435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=465910 $D=103
M3053 4437 WL_237 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=466400 $D=103
M3054 3962 WL_238 4439 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=469310 $D=103
M3055 4441 WL_239 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=469800 $D=103
M3056 3962 WL_240 4443 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=472710 $D=103
M3057 4445 WL_241 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=473200 $D=103
M3058 3962 WL_242 4447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=476110 $D=103
M3059 4449 WL_243 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=476600 $D=103
M3060 3962 WL_244 4451 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=479510 $D=103
M3061 4453 WL_245 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=480000 $D=103
M3062 3962 WL_246 4455 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=482910 $D=103
M3063 4457 WL_247 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=483400 $D=103
M3064 3962 WL_248 4459 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=486310 $D=103
M3065 4461 WL_249 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=486800 $D=103
M3066 3962 WL_250 4463 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=489710 $D=103
M3067 4465 WL_251 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=490200 $D=103
M3068 3962 WL_252 4467 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=493110 $D=103
M3069 4469 WL_253 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=493600 $D=103
M3070 3962 WL_254 4471 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=496510 $D=103
M3071 4473 WL_255 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118890 $Y=497000 $D=103
M3072 3961 WL_0 3964 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=64710 $D=103
M3073 3966 WL_1 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=65200 $D=103
M3074 3961 WL_2 3968 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=68110 $D=103
M3075 3970 WL_3 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=68600 $D=103
M3076 3961 WL_4 3972 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=71510 $D=103
M3077 3974 WL_5 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=72000 $D=103
M3078 3961 WL_6 3976 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=74910 $D=103
M3079 3978 WL_7 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=75400 $D=103
M3080 3961 WL_8 3980 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=78310 $D=103
M3081 3982 WL_9 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=78800 $D=103
M3082 3961 WL_10 3984 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=81710 $D=103
M3083 3986 WL_11 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=82200 $D=103
M3084 3961 WL_12 3988 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=85110 $D=103
M3085 3990 WL_13 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=85600 $D=103
M3086 3961 WL_14 3992 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=88510 $D=103
M3087 3994 WL_15 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=89000 $D=103
M3088 3961 WL_16 3996 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=91910 $D=103
M3089 3998 WL_17 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=92400 $D=103
M3090 3961 WL_18 4000 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=95310 $D=103
M3091 4002 WL_19 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=95800 $D=103
M3092 3961 WL_20 4004 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=98710 $D=103
M3093 4006 WL_21 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=99200 $D=103
M3094 3961 WL_22 4008 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=102110 $D=103
M3095 4010 WL_23 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=102600 $D=103
M3096 3961 WL_24 4012 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=105510 $D=103
M3097 4014 WL_25 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=106000 $D=103
M3098 3961 WL_26 4016 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=108910 $D=103
M3099 4018 WL_27 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=109400 $D=103
M3100 3961 WL_28 4020 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=112310 $D=103
M3101 4022 WL_29 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=112800 $D=103
M3102 3961 WL_30 4024 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=115710 $D=103
M3103 4026 WL_31 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=116200 $D=103
M3104 3961 WL_32 4028 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=119110 $D=103
M3105 4030 WL_33 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=119600 $D=103
M3106 3961 WL_34 4032 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=122510 $D=103
M3107 4034 WL_35 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=123000 $D=103
M3108 3961 WL_36 4036 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=125910 $D=103
M3109 4038 WL_37 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=126400 $D=103
M3110 3961 WL_38 4040 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=129310 $D=103
M3111 4042 WL_39 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=129800 $D=103
M3112 3961 WL_40 4044 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=132710 $D=103
M3113 4046 WL_41 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=133200 $D=103
M3114 3961 WL_42 4048 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=136110 $D=103
M3115 4050 WL_43 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=136600 $D=103
M3116 3961 WL_44 4052 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=139510 $D=103
M3117 4054 WL_45 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=140000 $D=103
M3118 3961 WL_46 4056 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=142910 $D=103
M3119 4058 WL_47 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=143400 $D=103
M3120 3961 WL_48 4060 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=146310 $D=103
M3121 4062 WL_49 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=146800 $D=103
M3122 3961 WL_50 4064 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=149710 $D=103
M3123 4066 WL_51 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=150200 $D=103
M3124 3961 WL_52 4068 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=153110 $D=103
M3125 4070 WL_53 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=153600 $D=103
M3126 3961 WL_54 4072 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=156510 $D=103
M3127 4074 WL_55 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=157000 $D=103
M3128 3961 WL_56 4076 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=159910 $D=103
M3129 4078 WL_57 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=160400 $D=103
M3130 3961 WL_58 4080 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=163310 $D=103
M3131 4082 WL_59 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=163800 $D=103
M3132 3961 WL_60 4084 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=166710 $D=103
M3133 4086 WL_61 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=167200 $D=103
M3134 3961 WL_62 4088 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=170110 $D=103
M3135 4090 WL_63 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=170600 $D=103
M3136 3961 WL_64 4092 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=173510 $D=103
M3137 4094 WL_65 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=174000 $D=103
M3138 3961 WL_66 4096 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=176910 $D=103
M3139 4098 WL_67 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=177400 $D=103
M3140 3961 WL_68 4100 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=180310 $D=103
M3141 4102 WL_69 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=180800 $D=103
M3142 3961 WL_70 4104 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=183710 $D=103
M3143 4106 WL_71 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=184200 $D=103
M3144 3961 WL_72 4108 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=187110 $D=103
M3145 4110 WL_73 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=187600 $D=103
M3146 3961 WL_74 4112 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=190510 $D=103
M3147 4114 WL_75 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=191000 $D=103
M3148 3961 WL_76 4116 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=193910 $D=103
M3149 4118 WL_77 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=194400 $D=103
M3150 3961 WL_78 4120 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=197310 $D=103
M3151 4122 WL_79 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=197800 $D=103
M3152 3961 WL_80 4124 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=200710 $D=103
M3153 4126 WL_81 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=201200 $D=103
M3154 3961 WL_82 4128 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=204110 $D=103
M3155 4130 WL_83 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=204600 $D=103
M3156 3961 WL_84 4132 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=207510 $D=103
M3157 4134 WL_85 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=208000 $D=103
M3158 3961 WL_86 4136 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=210910 $D=103
M3159 4138 WL_87 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=211400 $D=103
M3160 3961 WL_88 4140 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=214310 $D=103
M3161 4142 WL_89 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=214800 $D=103
M3162 3961 WL_90 4144 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=217710 $D=103
M3163 4146 WL_91 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=218200 $D=103
M3164 3961 WL_92 4148 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=221110 $D=103
M3165 4150 WL_93 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=221600 $D=103
M3166 3961 WL_94 4152 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=224510 $D=103
M3167 4154 WL_95 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=225000 $D=103
M3168 3961 WL_96 4156 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=227910 $D=103
M3169 4158 WL_97 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=228400 $D=103
M3170 3961 WL_98 4160 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=231310 $D=103
M3171 4162 WL_99 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=231800 $D=103
M3172 3961 WL_100 4164 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=234710 $D=103
M3173 4166 WL_101 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=235200 $D=103
M3174 3961 WL_102 4168 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=238110 $D=103
M3175 4170 WL_103 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=238600 $D=103
M3176 3961 WL_104 4172 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=241510 $D=103
M3177 4174 WL_105 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=242000 $D=103
M3178 3961 WL_106 4176 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=244910 $D=103
M3179 4178 WL_107 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=245400 $D=103
M3180 3961 WL_108 4180 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=248310 $D=103
M3181 4182 WL_109 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=248800 $D=103
M3182 3961 WL_110 4184 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=251710 $D=103
M3183 4186 WL_111 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=252200 $D=103
M3184 3961 WL_112 4188 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=255110 $D=103
M3185 4190 WL_113 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=255600 $D=103
M3186 3961 WL_114 4192 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=258510 $D=103
M3187 4194 WL_115 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=259000 $D=103
M3188 3961 WL_116 4196 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=261910 $D=103
M3189 4198 WL_117 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=262400 $D=103
M3190 3961 WL_118 4200 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=265310 $D=103
M3191 4202 WL_119 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=265800 $D=103
M3192 3961 WL_120 4204 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=268710 $D=103
M3193 4206 WL_121 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=269200 $D=103
M3194 3961 WL_122 4208 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=272110 $D=103
M3195 4210 WL_123 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=272600 $D=103
M3196 3961 WL_124 4212 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=275510 $D=103
M3197 4214 WL_125 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=276000 $D=103
M3198 3961 WL_126 4216 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=278910 $D=103
M3199 4218 WL_127 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=279400 $D=103
M3200 3961 WL_128 4220 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=282310 $D=103
M3201 4222 WL_129 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=282800 $D=103
M3202 3961 WL_130 4224 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=285710 $D=103
M3203 4226 WL_131 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=286200 $D=103
M3204 3961 WL_132 4228 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=289110 $D=103
M3205 4230 WL_133 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=289600 $D=103
M3206 3961 WL_134 4232 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=292510 $D=103
M3207 4234 WL_135 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=293000 $D=103
M3208 3961 WL_136 4236 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=295910 $D=103
M3209 4238 WL_137 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=296400 $D=103
M3210 3961 WL_138 4240 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=299310 $D=103
M3211 4242 WL_139 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=299800 $D=103
M3212 3961 WL_140 4244 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=302710 $D=103
M3213 4246 WL_141 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=303200 $D=103
M3214 3961 WL_142 4248 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=306110 $D=103
M3215 4250 WL_143 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=306600 $D=103
M3216 3961 WL_144 4252 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=309510 $D=103
M3217 4254 WL_145 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=310000 $D=103
M3218 3961 WL_146 4256 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=312910 $D=103
M3219 4258 WL_147 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=313400 $D=103
M3220 3961 WL_148 4260 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=316310 $D=103
M3221 4262 WL_149 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=316800 $D=103
M3222 3961 WL_150 4264 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=319710 $D=103
M3223 4266 WL_151 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=320200 $D=103
M3224 3961 WL_152 4268 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=323110 $D=103
M3225 4270 WL_153 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=323600 $D=103
M3226 3961 WL_154 4272 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=326510 $D=103
M3227 4274 WL_155 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=327000 $D=103
M3228 3961 WL_156 4276 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=329910 $D=103
M3229 4278 WL_157 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=330400 $D=103
M3230 3961 WL_158 4280 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=333310 $D=103
M3231 4282 WL_159 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=333800 $D=103
M3232 3961 WL_160 4284 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=336710 $D=103
M3233 4286 WL_161 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=337200 $D=103
M3234 3961 WL_162 4288 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=340110 $D=103
M3235 4290 WL_163 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=340600 $D=103
M3236 3961 WL_164 4292 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=343510 $D=103
M3237 4294 WL_165 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=344000 $D=103
M3238 3961 WL_166 4296 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=346910 $D=103
M3239 4298 WL_167 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=347400 $D=103
M3240 3961 WL_168 4300 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=350310 $D=103
M3241 4302 WL_169 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=350800 $D=103
M3242 3961 WL_170 4304 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=353710 $D=103
M3243 4306 WL_171 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=354200 $D=103
M3244 3961 WL_172 4308 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=357110 $D=103
M3245 4310 WL_173 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=357600 $D=103
M3246 3961 WL_174 4312 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=360510 $D=103
M3247 4314 WL_175 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=361000 $D=103
M3248 3961 WL_176 4316 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=363910 $D=103
M3249 4318 WL_177 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=364400 $D=103
M3250 3961 WL_178 4320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=367310 $D=103
M3251 4322 WL_179 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=367800 $D=103
M3252 3961 WL_180 4324 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=370710 $D=103
M3253 4326 WL_181 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=371200 $D=103
M3254 3961 WL_182 4328 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=374110 $D=103
M3255 4330 WL_183 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=374600 $D=103
M3256 3961 WL_184 4332 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=377510 $D=103
M3257 4334 WL_185 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=378000 $D=103
M3258 3961 WL_186 4336 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=380910 $D=103
M3259 4338 WL_187 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=381400 $D=103
M3260 3961 WL_188 4340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=384310 $D=103
M3261 4342 WL_189 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=384800 $D=103
M3262 3961 WL_190 4344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=387710 $D=103
M3263 4346 WL_191 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=388200 $D=103
M3264 3961 WL_192 4348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=391110 $D=103
M3265 4350 WL_193 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=391600 $D=103
M3266 3961 WL_194 4352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=394510 $D=103
M3267 4354 WL_195 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=395000 $D=103
M3268 3961 WL_196 4356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=397910 $D=103
M3269 4358 WL_197 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=398400 $D=103
M3270 3961 WL_198 4360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=401310 $D=103
M3271 4362 WL_199 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=401800 $D=103
M3272 3961 WL_200 4364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=404710 $D=103
M3273 4366 WL_201 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=405200 $D=103
M3274 3961 WL_202 4368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=408110 $D=103
M3275 4370 WL_203 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=408600 $D=103
M3276 3961 WL_204 4372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=411510 $D=103
M3277 4374 WL_205 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=412000 $D=103
M3278 3961 WL_206 4376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=414910 $D=103
M3279 4378 WL_207 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=415400 $D=103
M3280 3961 WL_208 4380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=418310 $D=103
M3281 4382 WL_209 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=418800 $D=103
M3282 3961 WL_210 4384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=421710 $D=103
M3283 4386 WL_211 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=422200 $D=103
M3284 3961 WL_212 4388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=425110 $D=103
M3285 4390 WL_213 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=425600 $D=103
M3286 3961 WL_214 4392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=428510 $D=103
M3287 4394 WL_215 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=429000 $D=103
M3288 3961 WL_216 4396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=431910 $D=103
M3289 4398 WL_217 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=432400 $D=103
M3290 3961 WL_218 4400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=435310 $D=103
M3291 4402 WL_219 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=435800 $D=103
M3292 3961 WL_220 4404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=438710 $D=103
M3293 4406 WL_221 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=439200 $D=103
M3294 3961 WL_222 4408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=442110 $D=103
M3295 4410 WL_223 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=442600 $D=103
M3296 3961 WL_224 4412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=445510 $D=103
M3297 4414 WL_225 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=446000 $D=103
M3298 3961 WL_226 4416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=448910 $D=103
M3299 4418 WL_227 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=449400 $D=103
M3300 3961 WL_228 4420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=452310 $D=103
M3301 4422 WL_229 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=452800 $D=103
M3302 3961 WL_230 4424 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=455710 $D=103
M3303 4426 WL_231 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=456200 $D=103
M3304 3961 WL_232 4428 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=459110 $D=103
M3305 4430 WL_233 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=459600 $D=103
M3306 3961 WL_234 4432 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=462510 $D=103
M3307 4434 WL_235 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=463000 $D=103
M3308 3961 WL_236 4436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=465910 $D=103
M3309 4438 WL_237 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=466400 $D=103
M3310 3961 WL_238 4440 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=469310 $D=103
M3311 4442 WL_239 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=469800 $D=103
M3312 3961 WL_240 4444 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=472710 $D=103
M3313 4446 WL_241 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=473200 $D=103
M3314 3961 WL_242 4448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=476110 $D=103
M3315 4450 WL_243 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=476600 $D=103
M3316 3961 WL_244 4452 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=479510 $D=103
M3317 4454 WL_245 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=480000 $D=103
M3318 3961 WL_246 4456 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=482910 $D=103
M3319 4458 WL_247 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=483400 $D=103
M3320 3961 WL_248 4460 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=486310 $D=103
M3321 4462 WL_249 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=486800 $D=103
M3322 3961 WL_250 4464 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=489710 $D=103
M3323 4466 WL_251 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=490200 $D=103
M3324 3961 WL_252 4468 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=493110 $D=103
M3325 4470 WL_253 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=493600 $D=103
M3326 3961 WL_254 4472 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=496510 $D=103
M3327 4474 WL_255 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137750 $Y=497000 $D=103
M3328 620 WL_0 4475 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=64710 $D=103
M3329 4476 WL_1 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=65200 $D=103
M3330 620 WL_2 4477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=68110 $D=103
M3331 4478 WL_3 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=68600 $D=103
M3332 620 WL_4 4479 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=71510 $D=103
M3333 4480 WL_5 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=72000 $D=103
M3334 620 WL_6 4481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=74910 $D=103
M3335 4482 WL_7 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=75400 $D=103
M3336 620 WL_8 4483 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=78310 $D=103
M3337 4484 WL_9 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=78800 $D=103
M3338 620 WL_10 4485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=81710 $D=103
M3339 4486 WL_11 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=82200 $D=103
M3340 620 WL_12 4487 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=85110 $D=103
M3341 4488 WL_13 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=85600 $D=103
M3342 620 WL_14 4489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=88510 $D=103
M3343 4490 WL_15 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=89000 $D=103
M3344 620 WL_16 4491 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=91910 $D=103
M3345 4492 WL_17 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=92400 $D=103
M3346 620 WL_18 4493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=95310 $D=103
M3347 4494 WL_19 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=95800 $D=103
M3348 620 WL_20 4495 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=98710 $D=103
M3349 4496 WL_21 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=99200 $D=103
M3350 620 WL_22 4497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=102110 $D=103
M3351 4498 WL_23 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=102600 $D=103
M3352 620 WL_24 4499 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=105510 $D=103
M3353 4500 WL_25 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=106000 $D=103
M3354 620 WL_26 4501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=108910 $D=103
M3355 4502 WL_27 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=109400 $D=103
M3356 620 WL_28 4503 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=112310 $D=103
M3357 4504 WL_29 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=112800 $D=103
M3358 620 WL_30 4505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=115710 $D=103
M3359 4506 WL_31 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=116200 $D=103
M3360 620 WL_32 4507 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=119110 $D=103
M3361 4508 WL_33 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=119600 $D=103
M3362 620 WL_34 4509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=122510 $D=103
M3363 4510 WL_35 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=123000 $D=103
M3364 620 WL_36 4511 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=125910 $D=103
M3365 4512 WL_37 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=126400 $D=103
M3366 620 WL_38 4513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=129310 $D=103
M3367 4514 WL_39 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=129800 $D=103
M3368 620 WL_40 4515 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=132710 $D=103
M3369 4516 WL_41 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=133200 $D=103
M3370 620 WL_42 4517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=136110 $D=103
M3371 4518 WL_43 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=136600 $D=103
M3372 620 WL_44 4519 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=139510 $D=103
M3373 4520 WL_45 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=140000 $D=103
M3374 620 WL_46 4521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=142910 $D=103
M3375 4522 WL_47 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=143400 $D=103
M3376 620 WL_48 4523 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=146310 $D=103
M3377 4524 WL_49 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=146800 $D=103
M3378 620 WL_50 4525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=149710 $D=103
M3379 4526 WL_51 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=150200 $D=103
M3380 620 WL_52 4527 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=153110 $D=103
M3381 4528 WL_53 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=153600 $D=103
M3382 620 WL_54 4529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=156510 $D=103
M3383 4530 WL_55 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=157000 $D=103
M3384 620 WL_56 4531 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=159910 $D=103
M3385 4532 WL_57 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=160400 $D=103
M3386 620 WL_58 4533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=163310 $D=103
M3387 4534 WL_59 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=163800 $D=103
M3388 620 WL_60 4535 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=166710 $D=103
M3389 4536 WL_61 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=167200 $D=103
M3390 620 WL_62 4537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=170110 $D=103
M3391 4538 WL_63 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=170600 $D=103
M3392 620 WL_64 4539 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=173510 $D=103
M3393 4540 WL_65 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=174000 $D=103
M3394 620 WL_66 4541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=176910 $D=103
M3395 4542 WL_67 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=177400 $D=103
M3396 620 WL_68 4543 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=180310 $D=103
M3397 4544 WL_69 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=180800 $D=103
M3398 620 WL_70 4545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=183710 $D=103
M3399 4546 WL_71 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=184200 $D=103
M3400 620 WL_72 4547 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=187110 $D=103
M3401 4548 WL_73 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=187600 $D=103
M3402 620 WL_74 4549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=190510 $D=103
M3403 4550 WL_75 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=191000 $D=103
M3404 620 WL_76 4551 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=193910 $D=103
M3405 4552 WL_77 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=194400 $D=103
M3406 620 WL_78 4553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=197310 $D=103
M3407 4554 WL_79 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=197800 $D=103
M3408 620 WL_80 4555 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=200710 $D=103
M3409 4556 WL_81 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=201200 $D=103
M3410 620 WL_82 4557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=204110 $D=103
M3411 4558 WL_83 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=204600 $D=103
M3412 620 WL_84 4559 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=207510 $D=103
M3413 4560 WL_85 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=208000 $D=103
M3414 620 WL_86 4561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=210910 $D=103
M3415 4562 WL_87 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=211400 $D=103
M3416 620 WL_88 4563 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=214310 $D=103
M3417 4564 WL_89 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=214800 $D=103
M3418 620 WL_90 4565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=217710 $D=103
M3419 4566 WL_91 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=218200 $D=103
M3420 620 WL_92 4567 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=221110 $D=103
M3421 4568 WL_93 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=221600 $D=103
M3422 620 WL_94 4569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=224510 $D=103
M3423 4570 WL_95 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=225000 $D=103
M3424 620 WL_96 4571 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=227910 $D=103
M3425 4572 WL_97 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=228400 $D=103
M3426 620 WL_98 4573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=231310 $D=103
M3427 4574 WL_99 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=231800 $D=103
M3428 620 WL_100 4575 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=234710 $D=103
M3429 4576 WL_101 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=235200 $D=103
M3430 620 WL_102 4577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=238110 $D=103
M3431 4578 WL_103 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=238600 $D=103
M3432 620 WL_104 4579 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=241510 $D=103
M3433 4580 WL_105 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=242000 $D=103
M3434 620 WL_106 4581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=244910 $D=103
M3435 4582 WL_107 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=245400 $D=103
M3436 620 WL_108 4583 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=248310 $D=103
M3437 4584 WL_109 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=248800 $D=103
M3438 620 WL_110 4585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=251710 $D=103
M3439 4586 WL_111 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=252200 $D=103
M3440 620 WL_112 4587 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=255110 $D=103
M3441 4588 WL_113 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=255600 $D=103
M3442 620 WL_114 4589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=258510 $D=103
M3443 4590 WL_115 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=259000 $D=103
M3444 620 WL_116 4591 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=261910 $D=103
M3445 4592 WL_117 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=262400 $D=103
M3446 620 WL_118 4593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=265310 $D=103
M3447 4594 WL_119 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=265800 $D=103
M3448 620 WL_120 4595 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=268710 $D=103
M3449 4596 WL_121 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=269200 $D=103
M3450 620 WL_122 4597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=272110 $D=103
M3451 4598 WL_123 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=272600 $D=103
M3452 620 WL_124 4599 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=275510 $D=103
M3453 4600 WL_125 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=276000 $D=103
M3454 620 WL_126 4601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=278910 $D=103
M3455 4602 WL_127 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=279400 $D=103
M3456 620 WL_128 4603 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=282310 $D=103
M3457 4604 WL_129 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=282800 $D=103
M3458 620 WL_130 4605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=285710 $D=103
M3459 4606 WL_131 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=286200 $D=103
M3460 620 WL_132 4607 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=289110 $D=103
M3461 4608 WL_133 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=289600 $D=103
M3462 620 WL_134 4609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=292510 $D=103
M3463 4610 WL_135 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=293000 $D=103
M3464 620 WL_136 4611 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=295910 $D=103
M3465 4612 WL_137 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=296400 $D=103
M3466 620 WL_138 4613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=299310 $D=103
M3467 4614 WL_139 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=299800 $D=103
M3468 620 WL_140 4615 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=302710 $D=103
M3469 4616 WL_141 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=303200 $D=103
M3470 620 WL_142 4617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=306110 $D=103
M3471 4618 WL_143 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=306600 $D=103
M3472 620 WL_144 4619 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=309510 $D=103
M3473 4620 WL_145 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=310000 $D=103
M3474 620 WL_146 4621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=312910 $D=103
M3475 4622 WL_147 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=313400 $D=103
M3476 620 WL_148 4623 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=316310 $D=103
M3477 4624 WL_149 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=316800 $D=103
M3478 620 WL_150 4625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=319710 $D=103
M3479 4626 WL_151 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=320200 $D=103
M3480 620 WL_152 4627 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=323110 $D=103
M3481 4628 WL_153 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=323600 $D=103
M3482 620 WL_154 4629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=326510 $D=103
M3483 4630 WL_155 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=327000 $D=103
M3484 620 WL_156 4631 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=329910 $D=103
M3485 4632 WL_157 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=330400 $D=103
M3486 620 WL_158 4633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=333310 $D=103
M3487 4634 WL_159 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=333800 $D=103
M3488 620 WL_160 4635 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=336710 $D=103
M3489 4636 WL_161 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=337200 $D=103
M3490 620 WL_162 4637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=340110 $D=103
M3491 4638 WL_163 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=340600 $D=103
M3492 620 WL_164 4639 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=343510 $D=103
M3493 4640 WL_165 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=344000 $D=103
M3494 620 WL_166 4641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=346910 $D=103
M3495 4642 WL_167 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=347400 $D=103
M3496 620 WL_168 4643 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=350310 $D=103
M3497 4644 WL_169 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=350800 $D=103
M3498 620 WL_170 4645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=353710 $D=103
M3499 4646 WL_171 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=354200 $D=103
M3500 620 WL_172 4647 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=357110 $D=103
M3501 4648 WL_173 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=357600 $D=103
M3502 620 WL_174 4649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=360510 $D=103
M3503 4650 WL_175 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=361000 $D=103
M3504 620 WL_176 4651 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=363910 $D=103
M3505 4652 WL_177 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=364400 $D=103
M3506 620 WL_178 4653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=367310 $D=103
M3507 4654 WL_179 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=367800 $D=103
M3508 620 WL_180 4655 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=370710 $D=103
M3509 4656 WL_181 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=371200 $D=103
M3510 620 WL_182 4657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=374110 $D=103
M3511 4658 WL_183 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=374600 $D=103
M3512 620 WL_184 4659 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=377510 $D=103
M3513 4660 WL_185 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=378000 $D=103
M3514 620 WL_186 4661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=380910 $D=103
M3515 4662 WL_187 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=381400 $D=103
M3516 620 WL_188 4663 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=384310 $D=103
M3517 4664 WL_189 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=384800 $D=103
M3518 620 WL_190 4665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=387710 $D=103
M3519 4666 WL_191 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=388200 $D=103
M3520 620 WL_192 4667 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=391110 $D=103
M3521 4668 WL_193 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=391600 $D=103
M3522 620 WL_194 4669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=394510 $D=103
M3523 4670 WL_195 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=395000 $D=103
M3524 620 WL_196 4671 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=397910 $D=103
M3525 4672 WL_197 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=398400 $D=103
M3526 620 WL_198 4673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=401310 $D=103
M3527 4674 WL_199 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=401800 $D=103
M3528 620 WL_200 4675 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=404710 $D=103
M3529 4676 WL_201 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=405200 $D=103
M3530 620 WL_202 4677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=408110 $D=103
M3531 4678 WL_203 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=408600 $D=103
M3532 620 WL_204 4679 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=411510 $D=103
M3533 4680 WL_205 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=412000 $D=103
M3534 620 WL_206 4681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=414910 $D=103
M3535 4682 WL_207 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=415400 $D=103
M3536 620 WL_208 4683 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=418310 $D=103
M3537 4684 WL_209 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=418800 $D=103
M3538 620 WL_210 4685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=421710 $D=103
M3539 4686 WL_211 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=422200 $D=103
M3540 620 WL_212 4687 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=425110 $D=103
M3541 4688 WL_213 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=425600 $D=103
M3542 620 WL_214 4689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=428510 $D=103
M3543 4690 WL_215 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=429000 $D=103
M3544 620 WL_216 4691 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=431910 $D=103
M3545 4692 WL_217 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=432400 $D=103
M3546 620 WL_218 4693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=435310 $D=103
M3547 4694 WL_219 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=435800 $D=103
M3548 620 WL_220 4695 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=438710 $D=103
M3549 4696 WL_221 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=439200 $D=103
M3550 620 WL_222 4697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=442110 $D=103
M3551 4698 WL_223 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=442600 $D=103
M3552 620 WL_224 4699 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=445510 $D=103
M3553 4700 WL_225 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=446000 $D=103
M3554 620 WL_226 4701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=448910 $D=103
M3555 4702 WL_227 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=449400 $D=103
M3556 620 WL_228 4703 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=452310 $D=103
M3557 4704 WL_229 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=452800 $D=103
M3558 620 WL_230 4705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=455710 $D=103
M3559 4706 WL_231 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=456200 $D=103
M3560 620 WL_232 4707 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=459110 $D=103
M3561 4708 WL_233 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=459600 $D=103
M3562 620 WL_234 4709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=462510 $D=103
M3563 4710 WL_235 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=463000 $D=103
M3564 620 WL_236 4711 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=465910 $D=103
M3565 4712 WL_237 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=466400 $D=103
M3566 620 WL_238 4713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=469310 $D=103
M3567 4714 WL_239 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=469800 $D=103
M3568 620 WL_240 4715 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=472710 $D=103
M3569 4716 WL_241 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=473200 $D=103
M3570 620 WL_242 4717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=476110 $D=103
M3571 4718 WL_243 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=476600 $D=103
M3572 620 WL_244 4719 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=479510 $D=103
M3573 4720 WL_245 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=480000 $D=103
M3574 620 WL_246 4721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=482910 $D=103
M3575 4722 WL_247 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=483400 $D=103
M3576 620 WL_248 4723 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=486310 $D=103
M3577 4724 WL_249 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=486800 $D=103
M3578 620 WL_250 4725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=489710 $D=103
M3579 4726 WL_251 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=490200 $D=103
M3580 620 WL_252 4727 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=493110 $D=103
M3581 4728 WL_253 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=493600 $D=103
M3582 620 WL_254 4729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=496510 $D=103
M3583 4730 WL_255 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138090 $Y=497000 $D=103
X3584 Q_0 VDD D_0 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 STUBDW_1 STUBDR__1 STUBDR_1 STUBDW__1 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 1134
+ 621 622 1135 623 1136 624 1137 625 1138 626 1139 627 1140 628 1141 629 1142 630 1143 631
+ 1144 632 1145 633 1146 634 1147 635 1148 636 1149 637 1150 638 1151 639 1152 640 1153 641
+ 1154 642 1155 643 1156 644 1157 645 1158 646 1159 647 1160 648 1161 649 1162 650 1163 651
+ 1164 652 1165 653 1166 654 1167 655 1168 656 1169 657 1170 658 1171 659 1172 660 1173 661
+ 1174 662 1175 663 1176 664 1177 665 1178 666 1179 667 1180 668 1181 669 1182 670 1183 671
+ 1184 672 1185 673 1186 674 1187 675 1188 676 1189 677 1190 678 1191 679 1192 680 1193 681
+ 1194 682 1195 683 1196 684 1197 685 1198 686 1199 687 1200 688 1201 689 1202 690 1203 691
+ 1204 692 1205 693 1206 694 1207 695 1208 696 1209 697 1210 698 1211 699 1212 700 1213 701
+ 1214 702 1215 703 1216 704 1217 705 1218 706 1219 707 1220 708 1221 709 1222 710 1223 711
+ 1224 712 1225 713 1226 714 1227 715 1228 716 1229 717 1230 718 1231 719 1232 720 1233 721
+ 1234 722 1235 723 1236 724 1237 725 1238 726 1239 727 1240 728 1241 729 1242 730 1243 731
+ 1244 732 1245 733 1246 734 1247 735 1248 736 1249 737 1250 738 1251 739 1252 740 1253 741
+ 1254 742 1255 743 1256 744 1257 745 1258 746 1259 747 1260 748 1261 749 1262 750 1263 751
+ 1264 752 1265 753 1266 754 1267 755 1268 756 1269 757 1270 758 1271 759 1272 760 1273 761
+ 1274 762 1275 763 1276 764 1277 765 1278 766 1279 767 1280 768 1281 769 1282 770 1283 771
+ 1284 772 1285 773 1286 774 1287 775 1288 776 1289 777 1290 778 1291 779 1292 780 1293 781
+ 1294 782 1295 783 1296 784 1297 785 1298 786 1299 787 1300 788 1301 789 1302 790 1303 791
+ 1304 792 1305 793 1306 794 1307 795 1308 796 1309 797 1310 798 1311 799 1312 800 1313 801
+ 1314 802 1315 803 1316 804 1317 805 1318 806 1319 807 1320 808 1321 809 1322 810 1323 811
+ 1324 812 1325 813 1326 814 1327 815 1328 816 1329 817 1330 818 1331 819 1332 820 1333 821
+ 1334 822 1335 823 1336 824 1337 825 1338 826 1339 827 1340 828 1341 829 1342 830 1343 831
+ 1344 832 1345 833 1346 834 1347 835 1348 836 1349 837 1350 838 1351 839 1352 840 1353 841
+ 1354 842 1355 843 1356 844 1357 845 1358 846 1359 847 1360 848 1361 849 1362 850 1363 851
+ 1364 852 1365 853 1366 854 1367 855 1368 856 1369 857 1370 858 1371 859 1372 860 1373 861
+ 1374 862 1375 863 1376 864 1377 865 1378 866 1379 867 1380 868 1381 869 1382 870 1383 871
+ 1384 872 1385 873 1386 874 1387 875 1388 876 1389 877 1390
+ ICV_89 $T=0 0 0 0 $X=-1000 $Y=-1000
X3585 Q_1 VDD D_1 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 561 562 563 564 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 1391
+ 1392 1393 1394 1395 1396 1397 1398 1399 1400 1401 1402 1403 1404 1405 1406 1407 1408 1409 1410 1411
+ 1412 1413 1414 1415 1416 1417 1418 1419 1420 1421 1422 1423 1424 1425 1426 1427 1428 1429 1430 1431
+ 1432 1433 1434 1435 1436 1437 1438 1439 1440 1441 1442 1443 1444 1445 1446 1447 1448 1449 1450 1451
+ 1452 1453 1454 1455 1456 1457 1458 1459 1460 1461 1462 1463 1464 1465 1466 1467 1468 1469 1470 1471
+ 1472 1473 1474 1475 1476 1477 1478 1479 1480 1481 1482 1483 1484 1485 1486 1487 1488 1489 1490 1491
+ 1492 1493 1494 1495 1496 1497 1498 1499 1500 1501 1502 1503 1504 1505 1506 1507 1508 1509 1510 1511
+ 1512 1513 1514 1515 1516 1517 1518 1519 1520 1521 1522 1523 1524 1525 1526 1527 1528 1529 1530 1531
+ 1532 1533 1534 1535 1536 1537 1538 1539 1540 1541 1542 1543 1544 1545 1546 1547 1548 1549 1550 1551
+ 1552 1553 1554 1555 1556 1557 1558 1559 1560 1561 1562 1563 1564 1565 1566 1567 1568 1569 1570 1571
+ 1572 1573 1574 1575 1576 1577 1578 1579 1580 1581 1582 1583 1584 1585 1586 1587 1588 1589 1590 1591
+ 1592 1593 1594 1595 1596 1597 1598 1599 1600 1601 1602 1603 1604 1605 1606 1607 1608 1609 1610 1611
+ 1612 1613 1614 1615 1616 1617 1618 1619 1620 1621 1622 1623 1624 1625 1626 1627 1628 1629 1630 1631
+ 1632 1633 1634 1635 1636 1637 1638 1639 1640 1641 1642 1643 1644 1645 1646 1647 1648 1649 1650 1651
+ 1652 1653 1654 1655 1656 1657 1658 1659 1660 1661 1662 1663 1664 1665 1666 1667 1668 1669 1670 1671
+ 1672 1673 1674 1675 1676 1677 1678 1679 1680 1681 1682 1683 1684 1685 1686 1687 1688 1689 1690 1691
+ 1692 1693 1694 1695 1696 1697 1698 1699 1700 1701 1702 1703 1704 1705 1706 1707 1708 1709 1710 1711
+ 1712 1713 1714 1715 1716 1717 1718 1719 1720 1721 1722 1723 1724 1725 1726 1727 1728 1729 1730 1731
+ 1732 1733 1734 1735 1736 1737 1738 1739 1740 1741 1742 1743 1744 1745 1746 1747 1748 1749 1750 1751
+ 1752 1753 1754 1755 1756 1757 1758 1759 1760 1761 1762 1763 1764 1765 1766 1767 1768 1769 1770 1771
+ 1772 1773 1774 1775 1776 1777 1778 1779 1780 1781 1782 1783 1784 1785 1786 1787 1788 1789 1790 1791
+ 1792 1793 1794 1795 1796 1797 1798 1799 1800 1801 1802 1803 1804 1805 1806 1807 1808 1809 1810 1811
+ 1812 1813 1814 1815 1816 1817 1818 1819 1820 1821 1822 1823 1824 1825 1826 1827 1828 1829 1830 1831
+ 1832 1833 1834 1835 1836 1837 1838 1839 1840 1841 1842 1843 1844 1845 1846 1847 1848 1849 1850 1851
+ 1852 1853 1854 1855 1856 1857 1858 1859 1860 1861 1862 1863 1864 1865 1866 1867 1868 1869 1870 1871
+ 1872 1873 1874 1875 1876 1877 1878 1879 1880 1881 1882 1883 1884 1885 1886 1887 1888 1889 1890 1891
+ 1892 1893 1894 1895 1896 1897 1898 1899 1900 1901 1902 1903 1904
+ ICV_84 $T=38400 0 1 180 $X=18200 $Y=-1000
X3586 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_98 $T=0 0 0 90 $X=37400 $Y=62320
X3587 Q_2 VDD D_2 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 565 566 567 568 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 1905
+ 1906 1907 1908 1909 1910 1911 1912 1913 1914 1915 1916 1917 1918 1919 1920 1921 1922 1923 1924 1925
+ 1926 1927 1928 1929 1930 1931 1932 1933 1934 1935 1936 1937 1938 1939 1940 1941 1942 1943 1944 1945
+ 1946 1947 1948 1949 1950 1951 1952 1953 1954 1955 1956 1957 1958 1959 1960 1961 1962 1963 1964 1965
+ 1966 1967 1968 1969 1970 1971 1972 1973 1974 1975 1976 1977 1978 1979 1980 1981 1982 1983 1984 1985
+ 1986 1987 1988 1989 1990 1991 1992 1993 1994 1995 1996 1997 1998 1999 2000 2001 2002 2003 2004 2005
+ 2006 2007 2008 2009 2010 2011 2012 2013 2014 2015 2016 2017 2018 2019 2020 2021 2022 2023 2024 2025
+ 2026 2027 2028 2029 2030 2031 2032 2033 2034 2035 2036 2037 2038 2039 2040 2041 2042 2043 2044 2045
+ 2046 2047 2048 2049 2050 2051 2052 2053 2054 2055 2056 2057 2058 2059 2060 2061 2062 2063 2064 2065
+ 2066 2067 2068 2069 2070 2071 2072 2073 2074 2075 2076 2077 2078 2079 2080 2081 2082 2083 2084 2085
+ 2086 2087 2088 2089 2090 2091 2092 2093 2094 2095 2096 2097 2098 2099 2100 2101 2102 2103 2104 2105
+ 2106 2107 2108 2109 2110 2111 2112 2113 2114 2115 2116 2117 2118 2119 2120 2121 2122 2123 2124 2125
+ 2126 2127 2128 2129 2130 2131 2132 2133 2134 2135 2136 2137 2138 2139 2140 2141 2142 2143 2144 2145
+ 2146 2147 2148 2149 2150 2151 2152 2153 2154 2155 2156 2157 2158 2159 2160 2161 2162 2163 2164 2165
+ 2166 2167 2168 2169 2170 2171 2172 2173 2174 2175 2176 2177 2178 2179 2180 2181 2182 2183 2184 2185
+ 2186 2187 2188 2189 2190 2191 2192 2193 2194 2195 2196 2197 2198 2199 2200 2201 2202 2203 2204 2205
+ 2206 2207 2208 2209 2210 2211 2212 2213 2214 2215 2216 2217 2218 2219 2220 2221 2222 2223 2224 2225
+ 2226 2227 2228 2229 2230 2231 2232 2233 2234 2235 2236 2237 2238 2239 2240 2241 2242 2243 2244 2245
+ 2246 2247 2248 2249 2250 2251 2252 2253 2254 2255 2256 2257 2258 2259 2260 2261 2262 2263 2264 2265
+ 2266 2267 2268 2269 2270 2271 2272 2273 2274 2275 2276 2277 2278 2279 2280 2281 2282 2283 2284 2285
+ 2286 2287 2288 2289 2290 2291 2292 2293 2294 2295 2296 2297 2298 2299 2300 2301 2302 2303 2304 2305
+ 2306 2307 2308 2309 2310 2311 2312 2313 2314 2315 2316 2317 2318 2319 2320 2321 2322 2323 2324 2325
+ 2326 2327 2328 2329 2330 2331 2332 2333 2334 2335 2336 2337 2338 2339 2340 2341 2342 2343 2344 2345
+ 2346 2347 2348 2349 2350 2351 2352 2353 2354 2355 2356 2357 2358 2359 2360 2361 2362 2363 2364 2365
+ 2366 2367 2368 2369 2370 2371 2372 2373 2374 2375 2376 2377 2378 2379 2380 2381 2382 2383 2384 2385
+ 2386 2387 2388 2389 2390 2391 2392 2393 2394 2395 2396 2397 2398 2399 2400 2401 2402 2403 2404 2405
+ 2406 2407 2408 2409 2410 2411 2412 2413 2414 2415 2416 2417 2418
+ ICV_79 $T=39600 0 0 0 $X=38600 $Y=-1000
X3588 Q_3 VDD D_3 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 569 570 571 572 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 2419
+ 2420 2421 2422 2423 2424 2425 2426 2427 2428 2429 2430 2431 2432 2433 2434 2435 2436 2437 2438 2439
+ 2440 2441 2442 2443 2444 2445 2446 2447 2448 2449 2450 2451 2452 2453 2454 2455 2456 2457 2458 2459
+ 2460 2461 2462 2463 2464 2465 2466 2467 2468 2469 2470 2471 2472 2473 2474 2475 2476 2477 2478 2479
+ 2480 2481 2482 2483 2484 2485 2486 2487 2488 2489 2490 2491 2492 2493 2494 2495 2496 2497 2498 2499
+ 2500 2501 2502 2503 2504 2505 2506 2507 2508 2509 2510 2511 2512 2513 2514 2515 2516 2517 2518 2519
+ 2520 2521 2522 2523 2524 2525 2526 2527 2528 2529 2530 2531 2532 2533 2534 2535 2536 2537 2538 2539
+ 2540 2541 2542 2543 2544 2545 2546 2547 2548 2549 2550 2551 2552 2553 2554 2555 2556 2557 2558 2559
+ 2560 2561 2562 2563 2564 2565 2566 2567 2568 2569 2570 2571 2572 2573 2574 2575 2576 2577 2578 2579
+ 2580 2581 2582 2583 2584 2585 2586 2587 2588 2589 2590 2591 2592 2593 2594 2595 2596 2597 2598 2599
+ 2600 2601 2602 2603 2604 2605 2606 2607 2608 2609 2610 2611 2612 2613 2614 2615 2616 2617 2618 2619
+ 2620 2621 2622 2623 2624 2625 2626 2627 2628 2629 2630 2631 2632 2633 2634 2635 2636 2637 2638 2639
+ 2640 2641 2642 2643 2644 2645 2646 2647 2648 2649 2650 2651 2652 2653 2654 2655 2656 2657 2658 2659
+ 2660 2661 2662 2663 2664 2665 2666 2667 2668 2669 2670 2671 2672 2673 2674 2675 2676 2677 2678 2679
+ 2680 2681 2682 2683 2684 2685 2686 2687 2688 2689 2690 2691 2692 2693 2694 2695 2696 2697 2698 2699
+ 2700 2701 2702 2703 2704 2705 2706 2707 2708 2709 2710 2711 2712 2713 2714 2715 2716 2717 2718 2719
+ 2720 2721 2722 2723 2724 2725 2726 2727 2728 2729 2730 2731 2732 2733 2734 2735 2736 2737 2738 2739
+ 2740 2741 2742 2743 2744 2745 2746 2747 2748 2749 2750 2751 2752 2753 2754 2755 2756 2757 2758 2759
+ 2760 2761 2762 2763 2764 2765 2766 2767 2768 2769 2770 2771 2772 2773 2774 2775 2776 2777 2778 2779
+ 2780 2781 2782 2783 2784 2785 2786 2787 2788 2789 2790 2791 2792 2793 2794 2795 2796 2797 2798 2799
+ 2800 2801 2802 2803 2804 2805 2806 2807 2808 2809 2810 2811 2812 2813 2814 2815 2816 2817 2818 2819
+ 2820 2821 2822 2823 2824 2825 2826 2827 2828 2829 2830 2831 2832 2833 2834 2835 2836 2837 2838 2839
+ 2840 2841 2842 2843 2844 2845 2846 2847 2848 2849 2850 2851 2852 2853 2854 2855 2856 2857 2858 2859
+ 2860 2861 2862 2863 2864 2865 2866 2867 2868 2869 2870 2871 2872 2873 2874 2875 2876 2877 2878 2879
+ 2880 2881 2882 2883 2884 2885 2886 2887 2888 2889 2890 2891 2892 2893 2894 2895 2896 2897 2898 2899
+ 2900 2901 2902 2903 2904 2905 2906 2907 2908 2909 2910 2911 2912 2913 2914 2915 2916 2917 2918 2919
+ 2920 2921 2922 2923 2924 2925 2926 2927 2928 2929 2930 2931 2932
+ ICV_74 $T=78000 0 1 180 $X=57800 $Y=-1000
X3589 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_97 $T=0 0 0 90 $X=77000 $Y=62320
X3590 Q_4 VDD D_4 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 573 574 575 576 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 2933
+ 2934 2935 2936 2937 2938 2939 2940 2941 2942 2943 2944 2945 2946 2947 2948 2949 2950 2951 2952 2953
+ 2954 2955 2956 2957 2958 2959 2960 2961 2962 2963 2964 2965 2966 2967 2968 2969 2970 2971 2972 2973
+ 2974 2975 2976 2977 2978 2979 2980 2981 2982 2983 2984 2985 2986 2987 2988 2989 2990 2991 2992 2993
+ 2994 2995 2996 2997 2998 2999 3000 3001 3002 3003 3004 3005 3006 3007 3008 3009 3010 3011 3012 3013
+ 3014 3015 3016 3017 3018 3019 3020 3021 3022 3023 3024 3025 3026 3027 3028 3029 3030 3031 3032 3033
+ 3034 3035 3036 3037 3038 3039 3040 3041 3042 3043 3044 3045 3046 3047 3048 3049 3050 3051 3052 3053
+ 3054 3055 3056 3057 3058 3059 3060 3061 3062 3063 3064 3065 3066 3067 3068 3069 3070 3071 3072 3073
+ 3074 3075 3076 3077 3078 3079 3080 3081 3082 3083 3084 3085 3086 3087 3088 3089 3090 3091 3092 3093
+ 3094 3095 3096 3097 3098 3099 3100 3101 3102 3103 3104 3105 3106 3107 3108 3109 3110 3111 3112 3113
+ 3114 3115 3116 3117 3118 3119 3120 3121 3122 3123 3124 3125 3126 3127 3128 3129 3130 3131 3132 3133
+ 3134 3135 3136 3137 3138 3139 3140 3141 3142 3143 3144 3145 3146 3147 3148 3149 3150 3151 3152 3153
+ 3154 3155 3156 3157 3158 3159 3160 3161 3162 3163 3164 3165 3166 3167 3168 3169 3170 3171 3172 3173
+ 3174 3175 3176 3177 3178 3179 3180 3181 3182 3183 3184 3185 3186 3187 3188 3189 3190 3191 3192 3193
+ 3194 3195 3196 3197 3198 3199 3200 3201 3202 3203 3204 3205 3206 3207 3208 3209 3210 3211 3212 3213
+ 3214 3215 3216 3217 3218 3219 3220 3221 3222 3223 3224 3225 3226 3227 3228 3229 3230 3231 3232 3233
+ 3234 3235 3236 3237 3238 3239 3240 3241 3242 3243 3244 3245 3246 3247 3248 3249 3250 3251 3252 3253
+ 3254 3255 3256 3257 3258 3259 3260 3261 3262 3263 3264 3265 3266 3267 3268 3269 3270 3271 3272 3273
+ 3274 3275 3276 3277 3278 3279 3280 3281 3282 3283 3284 3285 3286 3287 3288 3289 3290 3291 3292 3293
+ 3294 3295 3296 3297 3298 3299 3300 3301 3302 3303 3304 3305 3306 3307 3308 3309 3310 3311 3312 3313
+ 3314 3315 3316 3317 3318 3319 3320 3321 3322 3323 3324 3325 3326 3327 3328 3329 3330 3331 3332 3333
+ 3334 3335 3336 3337 3338 3339 3340 3341 3342 3343 3344 3345 3346 3347 3348 3349 3350 3351 3352 3353
+ 3354 3355 3356 3357 3358 3359 3360 3361 3362 3363 3364 3365 3366 3367 3368 3369 3370 3371 3372 3373
+ 3374 3375 3376 3377 3378 3379 3380 3381 3382 3383 3384 3385 3386 3387 3388 3389 3390 3391 3392 3393
+ 3394 3395 3396 3397 3398 3399 3400 3401 3402 3403 3404 3405 3406 3407 3408 3409 3410 3411 3412 3413
+ 3414 3415 3416 3417 3418 3419 3420 3421 3422 3423 3424 3425 3426 3427 3428 3429 3430 3431 3432 3433
+ 3434 3435 3436 3437 3438 3439 3440 3441 3442 3443 3444 3445 3446
+ ICV_69 $T=79200 0 0 0 $X=78200 $Y=-1000
X3591 Q_5 VDD D_5 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 577 578 579 580 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 3447
+ 3448 3449 3450 3451 3452 3453 3454 3455 3456 3457 3458 3459 3460 3461 3462 3463 3464 3465 3466 3467
+ 3468 3469 3470 3471 3472 3473 3474 3475 3476 3477 3478 3479 3480 3481 3482 3483 3484 3485 3486 3487
+ 3488 3489 3490 3491 3492 3493 3494 3495 3496 3497 3498 3499 3500 3501 3502 3503 3504 3505 3506 3507
+ 3508 3509 3510 3511 3512 3513 3514 3515 3516 3517 3518 3519 3520 3521 3522 3523 3524 3525 3526 3527
+ 3528 3529 3530 3531 3532 3533 3534 3535 3536 3537 3538 3539 3540 3541 3542 3543 3544 3545 3546 3547
+ 3548 3549 3550 3551 3552 3553 3554 3555 3556 3557 3558 3559 3560 3561 3562 3563 3564 3565 3566 3567
+ 3568 3569 3570 3571 3572 3573 3574 3575 3576 3577 3578 3579 3580 3581 3582 3583 3584 3585 3586 3587
+ 3588 3589 3590 3591 3592 3593 3594 3595 3596 3597 3598 3599 3600 3601 3602 3603 3604 3605 3606 3607
+ 3608 3609 3610 3611 3612 3613 3614 3615 3616 3617 3618 3619 3620 3621 3622 3623 3624 3625 3626 3627
+ 3628 3629 3630 3631 3632 3633 3634 3635 3636 3637 3638 3639 3640 3641 3642 3643 3644 3645 3646 3647
+ 3648 3649 3650 3651 3652 3653 3654 3655 3656 3657 3658 3659 3660 3661 3662 3663 3664 3665 3666 3667
+ 3668 3669 3670 3671 3672 3673 3674 3675 3676 3677 3678 3679 3680 3681 3682 3683 3684 3685 3686 3687
+ 3688 3689 3690 3691 3692 3693 3694 3695 3696 3697 3698 3699 3700 3701 3702 3703 3704 3705 3706 3707
+ 3708 3709 3710 3711 3712 3713 3714 3715 3716 3717 3718 3719 3720 3721 3722 3723 3724 3725 3726 3727
+ 3728 3729 3730 3731 3732 3733 3734 3735 3736 3737 3738 3739 3740 3741 3742 3743 3744 3745 3746 3747
+ 3748 3749 3750 3751 3752 3753 3754 3755 3756 3757 3758 3759 3760 3761 3762 3763 3764 3765 3766 3767
+ 3768 3769 3770 3771 3772 3773 3774 3775 3776 3777 3778 3779 3780 3781 3782 3783 3784 3785 3786 3787
+ 3788 3789 3790 3791 3792 3793 3794 3795 3796 3797 3798 3799 3800 3801 3802 3803 3804 3805 3806 3807
+ 3808 3809 3810 3811 3812 3813 3814 3815 3816 3817 3818 3819 3820 3821 3822 3823 3824 3825 3826 3827
+ 3828 3829 3830 3831 3832 3833 3834 3835 3836 3837 3838 3839 3840 3841 3842 3843 3844 3845 3846 3847
+ 3848 3849 3850 3851 3852 3853 3854 3855 3856 3857 3858 3859 3860 3861 3862 3863 3864 3865 3866 3867
+ 3868 3869 3870 3871 3872 3873 3874 3875 3876 3877 3878 3879 3880 3881 3882 3883 3884 3885 3886 3887
+ 3888 3889 3890 3891 3892 3893 3894 3895 3896 3897 3898 3899 3900 3901 3902 3903 3904 3905 3906 3907
+ 3908 3909 3910 3911 3912 3913 3914 3915 3916 3917 3918 3919 3920 3921 3922 3923 3924 3925 3926 3927
+ 3928 3929 3930 3931 3932 3933 3934 3935 3936 3937 3938 3939 3940 3941 3942 3943 3944 3945 3946 3947
+ 3948 3949 3950 3951 3952 3953 3954 3955 3956 3957 3958 3959 3960
+ ICV_64 $T=117600 0 1 180 $X=97400 $Y=-1000
X3592 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18
+ WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38
+ WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58
+ WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78
+ WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97 WL_98
+ WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118
+ WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137 WL_138
+ WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157 WL_158
+ WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177 WL_178
+ WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197 WL_198
+ WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217 WL_218
+ WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237 WL_238
+ WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ ICV_96 $T=0 0 0 90 $X=116600 $Y=62320
X3593 Q_6 VDD D_6 VSS WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15
+ WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35
+ WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55
+ WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75
+ WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95
+ WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115
+ WL_116 WL_117 WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135
+ WL_136 WL_137 WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155
+ WL_156 WL_157 WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175
+ WL_176 WL_177 WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195
+ WL_196 WL_197 WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215
+ WL_216 WL_217 WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235
+ WL_236 WL_237 WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255
+ WE GTP_0 OE_ GTP_1 581 582 583 584 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 3961
+ 3962 3963 3964 3965 3966 3967 3968 3969 3970 3971 3972 3973 3974 3975 3976 3977 3978 3979 3980 3981
+ 3982 3983 3984 3985 3986 3987 3988 3989 3990 3991 3992 3993 3994 3995 3996 3997 3998 3999 4000 4001
+ 4002 4003 4004 4005 4006 4007 4008 4009 4010 4011 4012 4013 4014 4015 4016 4017 4018 4019 4020 4021
+ 4022 4023 4024 4025 4026 4027 4028 4029 4030 4031 4032 4033 4034 4035 4036 4037 4038 4039 4040 4041
+ 4042 4043 4044 4045 4046 4047 4048 4049 4050 4051 4052 4053 4054 4055 4056 4057 4058 4059 4060 4061
+ 4062 4063 4064 4065 4066 4067 4068 4069 4070 4071 4072 4073 4074 4075 4076 4077 4078 4079 4080 4081
+ 4082 4083 4084 4085 4086 4087 4088 4089 4090 4091 4092 4093 4094 4095 4096 4097 4098 4099 4100 4101
+ 4102 4103 4104 4105 4106 4107 4108 4109 4110 4111 4112 4113 4114 4115 4116 4117 4118 4119 4120 4121
+ 4122 4123 4124 4125 4126 4127 4128 4129 4130 4131 4132 4133 4134 4135 4136 4137 4138 4139 4140 4141
+ 4142 4143 4144 4145 4146 4147 4148 4149 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161
+ 4162 4163 4164 4165 4166 4167 4168 4169 4170 4171 4172 4173 4174 4175 4176 4177 4178 4179 4180 4181
+ 4182 4183 4184 4185 4186 4187 4188 4189 4190 4191 4192 4193 4194 4195 4196 4197 4198 4199 4200 4201
+ 4202 4203 4204 4205 4206 4207 4208 4209 4210 4211 4212 4213 4214 4215 4216 4217 4218 4219 4220 4221
+ 4222 4223 4224 4225 4226 4227 4228 4229 4230 4231 4232 4233 4234 4235 4236 4237 4238 4239 4240 4241
+ 4242 4243 4244 4245 4246 4247 4248 4249 4250 4251 4252 4253 4254 4255 4256 4257 4258 4259 4260 4261
+ 4262 4263 4264 4265 4266 4267 4268 4269 4270 4271 4272 4273 4274 4275 4276 4277 4278 4279 4280 4281
+ 4282 4283 4284 4285 4286 4287 4288 4289 4290 4291 4292 4293 4294 4295 4296 4297 4298 4299 4300 4301
+ 4302 4303 4304 4305 4306 4307 4308 4309 4310 4311 4312 4313 4314 4315 4316 4317 4318 4319 4320 4321
+ 4322 4323 4324 4325 4326 4327 4328 4329 4330 4331 4332 4333 4334 4335 4336 4337 4338 4339 4340 4341
+ 4342 4343 4344 4345 4346 4347 4348 4349 4350 4351 4352 4353 4354 4355 4356 4357 4358 4359 4360 4361
+ 4362 4363 4364 4365 4366 4367 4368 4369 4370 4371 4372 4373 4374 4375 4376 4377 4378 4379 4380 4381
+ 4382 4383 4384 4385 4386 4387 4388 4389 4390 4391 4392 4393 4394 4395 4396 4397 4398 4399 4400 4401
+ 4402 4403 4404 4405 4406 4407 4408 4409 4410 4411 4412 4413 4414 4415 4416 4417 4418 4419 4420 4421
+ 4422 4423 4424 4425 4426 4427 4428 4429 4430 4431 4432 4433 4434 4435 4436 4437 4438 4439 4440 4441
+ 4442 4443 4444 4445 4446 4447 4448 4449 4450 4451 4452 4453 4454 4455 4456 4457 4458 4459 4460 4461
+ 4462 4463 4464 4465 4466 4467 4468 4469 4470 4471 4472 4473 4474
+ ICV_55 $T=118800 0 0 0 $X=117800 $Y=-1000
X3594 VSS VDD D_7 Q_7 585 588 587 586 A0 A0_ YP1_3 YP1_2 YP1_1 YP1_0 YP0_3 YP0_2 YP0_1 YP0_0 GTP_2 WE
+ GTP_0 OE_ GTP_1 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605
+ 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ ICV_91 $T=0 0 0 90 $X=137000 $Y=-1000
X3595 VSS VDD WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17
+ WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37
+ WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57
+ WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77
+ WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 WL_97
+ WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117
+ WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 WL_128 WL_129 WL_130 WL_131 WL_132 WL_133 WL_134 WL_135 WL_136 WL_137
+ WL_138 WL_139 WL_140 WL_141 WL_142 WL_143 WL_144 WL_145 WL_146 WL_147 WL_148 WL_149 WL_150 WL_151 WL_152 WL_153 WL_154 WL_155 WL_156 WL_157
+ WL_158 WL_159 WL_160 WL_161 WL_162 WL_163 WL_164 WL_165 WL_166 WL_167 WL_168 WL_169 WL_170 WL_171 WL_172 WL_173 WL_174 WL_175 WL_176 WL_177
+ WL_178 WL_179 WL_180 WL_181 WL_182 WL_183 WL_184 WL_185 WL_186 WL_187 WL_188 WL_189 WL_190 WL_191 WL_192 WL_193 WL_194 WL_195 WL_196 WL_197
+ WL_198 WL_199 WL_200 WL_201 WL_202 WL_203 WL_204 WL_205 WL_206 WL_207 WL_208 WL_209 WL_210 WL_211 WL_212 WL_213 WL_214 WL_215 WL_216 WL_217
+ WL_218 WL_219 WL_220 WL_221 WL_222 WL_223 WL_224 WL_225 WL_226 WL_227 WL_228 WL_229 WL_230 WL_231 WL_232 WL_233 WL_234 WL_235 WL_236 WL_237
+ WL_238 WL_239 WL_240 WL_241 WL_242 WL_243 WL_244 WL_245 WL_246 WL_247 WL_248 WL_249 WL_250 WL_251 WL_252 WL_253 WL_254 WL_255 619 618
+ 617 616 615 614 613 612 611 610 609 608 607 606 605 604 603 602 601 600 599 598
+ 597 596 595 594 593 592 591 590 4475 878 4476 879 4477 880 4478 881 4479 882 4480 883
+ 4481 884 4482 885 4483 886 4484 887 4485 888 4486 889 4487 890 4488 891 4489 892 4490 893
+ 4491 894 4492 895 4493 896 4494 897 4495 898 4496 899 4497 900 4498 901 4499 902 4500 903
+ 4501 904 4502 905 4503 906 4504 907 4505 908 4506 909 4507 910 4508 911 4509 912 4510 913
+ 4511 914 4512 915 4513 916 4514 917 4515 918 4516 919 4517 920 4518 921 4519 922 4520 923
+ 4521 924 4522 925 4523 926 4524 927 4525 928 4526 929 4527 930 4528 931 4529 932 4530 933
+ 4531 934 4532 935 4533 936 4534 937 4535 938 4536 939 4537 940 4538 941 4539 942 4540 943
+ 4541 944 4542 945 4543 946 4544 947 4545 948 4546 949 4547 950 4548 951 4549 952 4550 953
+ 4551 954 4552 955 4553 956 4554 957 4555 958 4556 959 4557 960 4558 961 4559 962 4560 963
+ 4561 964 4562 965 4563 966 4564 967 4565 968 4566 969 4567 970 4568 971 4569 972 4570 973
+ 4571 974 4572 975 4573 976 4574 977 4575 978 4576 979 4577 980 4578 981 4579 982 4580 983
+ 4581 984 4582 985 4583 986 4584 987 4585 988 4586 989 4587 990 4588 991 4589 992 4590 993
+ 4591 994 4592 995 4593 996 4594 997 4595 998 4596 999 4597 1000 4598 1001 4599 1002 4600 1003
+ 4601 1004 4602 1005 4603 1006 4604 1007 4605 1008 4606 1009 4607 1010 4608 1011 4609 1012 4610 1013
+ 4611 1014 4612 1015 4613 1016 4614 1017 4615 1018 4616 1019 4617 1020 4618 1021 4619 1022 4620 1023
+ 4621 1024 4622 1025 4623 1026 4624 1027 4625 1028 4626 1029 4627 1030 4628 1031 4629 1032 4630 1033
+ 4631 1034 4632 1035 4633 1036 4634 1037 4635 1038 4636 1039 4637 1040 4638 1041 4639 1042 4640 1043
+ 4641 1044 4642 1045 4643 1046 4644 1047 4645 1048 4646 1049 4647 1050 4648 1051 4649 1052 4650 1053
+ 4651 1054 4652 1055 4653 1056 4654 1057 4655 1058 4656 1059 4657 1060 4658 1061 4659 1062 4660 1063
+ 4661 1064 4662 1065 4663 1066 4664 1067 4665 1068 4666 1069 4667 1070 4668 1071 4669 1072 4670 1073
+ 4671 1074 4672 1075 4673 1076 4674 1077 4675 1078 4676 1079 4677 1080 4678 1081 4679 1082 4680 1083
+ 4681 1084 4682 1085 4683 1086 4684 1087 4685 1088 4686 1089 4687 1090 4688 1091 4689 1092 4690 1093
+ 4691 1094 4692 1095 4693 1096 4694 1097 4695 1098 4696 1099 4697 1100 4698 1101 4699 1102 4700 1103
+ 4701 1104 4702 1105 4703 1106 4704 1107 4705 1108 4706 1109 4707 1110 4708 1111 4709 1112 4710 1113
+ 4711 1114 4712 1115 4713 1116 4714 1117 4715 1118 4716 1119 4717 1120 4718 1121 4719 1122 4720 1123
+ 4721 1124 4722 1125 4723 1126 4724 1127 4725 1128 4726 1129 4727 1130 4728 1131 4729 1132 4730 1133
+ ICV_90 $T=0 0 0 90 $X=137000 $Y=61500
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT base_flme_nvpv 2 4 7 8
** N=18 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 4 8 7 4 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=380 $Y=850 $D=103
M1 8 7 4 4 lpnfet w=2e-07 l=1e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=850 $D=103
M2 2 8 7 2 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=370 $Y=260 $D=192
M3 8 7 2 2 lppfet w=1.5e-07 l=1.2e-07 m=1 par=1 nf=1 ngcon=1 $X=710 $Y=260 $D=192
.ENDS
***************************************
.SUBCKT SIGN_MEM VDD VSS D<7> Q<7> Q<6> D<6> D<5> Q<5> Q<4> D<4> D<3> Q<3> Q<2> D<2> D<1> Q<1> Q<0> D<0> A<11> A<10>
+ A<9> A<8> A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> CEN WEN CLK D<8> Q<8> Q<9> D<9> D<10> Q<10> Q<11>
+ D<11> D<12> Q<12> Q<13> D<13> D<14> Q<14> Q<15> D<15>
** N=5892 EP=49 IP=17697 FDC=420541
M0 4857 63 5115 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=74950 $D=103
M1 5116 64 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=75440 $D=103
M2 4857 65 5117 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=78350 $D=103
M3 5118 66 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=78840 $D=103
M4 4857 67 5119 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=81750 $D=103
M5 5120 68 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=82240 $D=103
M6 4857 69 5121 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=85150 $D=103
M7 5122 70 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=85640 $D=103
M8 4857 71 5123 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=88550 $D=103
M9 5124 72 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=89040 $D=103
M10 4857 73 5125 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=91950 $D=103
M11 5126 74 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=92440 $D=103
M12 4857 75 5127 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=95350 $D=103
M13 5128 76 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=95840 $D=103
M14 4857 77 5129 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=98750 $D=103
M15 5130 78 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=99240 $D=103
M16 4857 79 5131 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=102150 $D=103
M17 5132 80 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=102640 $D=103
M18 4857 81 5133 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=105550 $D=103
M19 5134 82 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=106040 $D=103
M20 4857 83 5135 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=108950 $D=103
M21 5136 84 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=109440 $D=103
M22 4857 85 5137 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=112350 $D=103
M23 5138 86 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=112840 $D=103
M24 4857 87 5139 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=115750 $D=103
M25 5140 88 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=116240 $D=103
M26 4857 89 5141 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=119150 $D=103
M27 5142 90 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=119640 $D=103
M28 4857 91 5143 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=122550 $D=103
M29 5144 92 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=123040 $D=103
M30 4857 93 5145 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=125950 $D=103
M31 5146 94 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=126440 $D=103
M32 4857 95 5147 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=129350 $D=103
M33 5148 96 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=129840 $D=103
M34 4857 97 5149 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=132750 $D=103
M35 5150 98 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=133240 $D=103
M36 4857 99 5151 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=136150 $D=103
M37 5152 100 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=136640 $D=103
M38 4857 101 5153 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=139550 $D=103
M39 5154 102 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=140040 $D=103
M40 4857 103 5155 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=142950 $D=103
M41 5156 104 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=143440 $D=103
M42 4857 105 5157 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=146350 $D=103
M43 5158 106 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=146840 $D=103
M44 4857 107 5159 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=149750 $D=103
M45 5160 108 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=150240 $D=103
M46 4857 109 5161 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=153150 $D=103
M47 5162 110 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=153640 $D=103
M48 4857 111 5163 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=156550 $D=103
M49 5164 112 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=157040 $D=103
M50 4857 113 5165 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=159950 $D=103
M51 5166 114 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=160440 $D=103
M52 4857 115 5167 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=163350 $D=103
M53 5168 116 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=163840 $D=103
M54 4857 117 5169 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=166750 $D=103
M55 5170 118 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=167240 $D=103
M56 4857 119 5171 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=170150 $D=103
M57 5172 120 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=170640 $D=103
M58 4857 121 5173 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=173550 $D=103
M59 5174 122 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=174040 $D=103
M60 4857 123 5175 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=176950 $D=103
M61 5176 124 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=177440 $D=103
M62 4857 125 5177 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=180350 $D=103
M63 5178 126 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=180840 $D=103
M64 4857 127 5179 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=183750 $D=103
M65 5180 128 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=184240 $D=103
M66 4857 129 5181 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=187150 $D=103
M67 5182 130 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=187640 $D=103
M68 4857 131 5183 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=190550 $D=103
M69 5184 132 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=191040 $D=103
M70 4857 133 5185 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=193950 $D=103
M71 5186 134 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=194440 $D=103
M72 4857 135 5187 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=197350 $D=103
M73 5188 136 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=197840 $D=103
M74 4857 137 5189 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=200750 $D=103
M75 5190 138 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=201240 $D=103
M76 4857 139 5191 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=204150 $D=103
M77 5192 140 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=204640 $D=103
M78 4857 141 5193 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=207550 $D=103
M79 5194 142 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=208040 $D=103
M80 4857 143 5195 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=210950 $D=103
M81 5196 144 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=211440 $D=103
M82 4857 145 5197 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=214350 $D=103
M83 5198 146 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=214840 $D=103
M84 4857 147 5199 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=217750 $D=103
M85 5200 148 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=218240 $D=103
M86 4857 149 5201 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=221150 $D=103
M87 5202 150 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=221640 $D=103
M88 4857 151 5203 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=224550 $D=103
M89 5204 152 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=225040 $D=103
M90 4857 153 5205 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=227950 $D=103
M91 5206 154 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=228440 $D=103
M92 4857 155 5207 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=231350 $D=103
M93 5208 156 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=231840 $D=103
M94 4857 157 5209 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=234750 $D=103
M95 5210 158 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=235240 $D=103
M96 4857 159 5211 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=238150 $D=103
M97 5212 160 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=238640 $D=103
M98 4857 161 5213 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=241550 $D=103
M99 5214 162 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=242040 $D=103
M100 4857 163 5215 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=244950 $D=103
M101 5216 164 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=245440 $D=103
M102 4857 165 5217 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=248350 $D=103
M103 5218 166 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=248840 $D=103
M104 4857 167 5219 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=251750 $D=103
M105 5220 168 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=252240 $D=103
M106 4857 169 5221 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=255150 $D=103
M107 5222 170 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=255640 $D=103
M108 4857 171 5223 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=258550 $D=103
M109 5224 172 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=259040 $D=103
M110 4857 173 5225 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=261950 $D=103
M111 5226 174 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=262440 $D=103
M112 4857 175 5227 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=265350 $D=103
M113 5228 176 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=265840 $D=103
M114 4857 177 5229 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=268750 $D=103
M115 5230 178 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=269240 $D=103
M116 4857 179 5231 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=272150 $D=103
M117 5232 180 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=272640 $D=103
M118 4857 181 5233 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=275550 $D=103
M119 5234 182 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=276040 $D=103
M120 4857 183 5235 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=278950 $D=103
M121 5236 184 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=279440 $D=103
M122 4857 185 5237 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=282350 $D=103
M123 5238 186 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=282840 $D=103
M124 4857 187 5239 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=285750 $D=103
M125 5240 188 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=286240 $D=103
M126 4857 189 5241 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=289150 $D=103
M127 5242 190 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=289640 $D=103
M128 4857 191 5243 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=292550 $D=103
M129 5244 192 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=293040 $D=103
M130 4857 193 5245 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=295950 $D=103
M131 5246 194 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=296440 $D=103
M132 4857 195 5247 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=299350 $D=103
M133 5248 196 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=299840 $D=103
M134 4857 197 5249 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=302750 $D=103
M135 5250 198 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=303240 $D=103
M136 4857 199 5251 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=306150 $D=103
M137 5252 200 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=306640 $D=103
M138 4857 201 5253 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=309550 $D=103
M139 5254 202 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=310040 $D=103
M140 4857 203 5255 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=312950 $D=103
M141 5256 204 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=313440 $D=103
M142 4857 205 5257 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=316350 $D=103
M143 5258 206 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=316840 $D=103
M144 4857 207 5259 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=319750 $D=103
M145 5260 208 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=320240 $D=103
M146 4857 209 5261 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=323150 $D=103
M147 5262 210 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=323640 $D=103
M148 4857 211 5263 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=326550 $D=103
M149 5264 212 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=327040 $D=103
M150 4857 213 5265 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=329950 $D=103
M151 5266 214 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=330440 $D=103
M152 4857 215 5267 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=333350 $D=103
M153 5268 216 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=333840 $D=103
M154 4857 217 5269 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=336750 $D=103
M155 5270 218 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=337240 $D=103
M156 4857 219 5271 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=340150 $D=103
M157 5272 220 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=340640 $D=103
M158 4857 221 5273 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=343550 $D=103
M159 5274 222 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=344040 $D=103
M160 4857 223 5275 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=346950 $D=103
M161 5276 224 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=347440 $D=103
M162 4857 225 5277 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=350350 $D=103
M163 5278 226 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=350840 $D=103
M164 4857 227 5279 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=353750 $D=103
M165 5280 228 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=354240 $D=103
M166 4857 229 5281 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=357150 $D=103
M167 5282 230 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=357640 $D=103
M168 4857 231 5283 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=360550 $D=103
M169 5284 232 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=361040 $D=103
M170 4857 233 5285 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=363950 $D=103
M171 5286 234 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=364440 $D=103
M172 4857 235 5287 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=367350 $D=103
M173 5288 236 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=367840 $D=103
M174 4857 237 5289 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=370750 $D=103
M175 5290 238 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=371240 $D=103
M176 4857 239 5291 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=374150 $D=103
M177 5292 240 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=374640 $D=103
M178 4857 241 5293 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=377550 $D=103
M179 5294 242 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=378040 $D=103
M180 4857 243 5295 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=380950 $D=103
M181 5296 244 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=381440 $D=103
M182 4857 245 5297 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=384350 $D=103
M183 5298 246 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=384840 $D=103
M184 4857 247 5299 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=387750 $D=103
M185 5300 248 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=388240 $D=103
M186 4857 249 5301 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=391150 $D=103
M187 5302 250 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=391640 $D=103
M188 4857 251 5303 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=394550 $D=103
M189 5304 252 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=395040 $D=103
M190 4857 253 5305 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=397950 $D=103
M191 5306 254 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=398440 $D=103
M192 4857 255 5307 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=401350 $D=103
M193 5308 256 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=401840 $D=103
M194 4857 257 5309 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=404750 $D=103
M195 5310 258 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=405240 $D=103
M196 4857 259 5311 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=408150 $D=103
M197 5312 260 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=408640 $D=103
M198 4857 261 5313 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=411550 $D=103
M199 5314 262 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=412040 $D=103
M200 4857 263 5315 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=414950 $D=103
M201 5316 264 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=415440 $D=103
M202 4857 265 5317 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=418350 $D=103
M203 5318 266 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=418840 $D=103
M204 4857 267 5319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=421750 $D=103
M205 5320 268 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=422240 $D=103
M206 4857 269 5321 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=425150 $D=103
M207 5322 270 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=425640 $D=103
M208 4857 271 5323 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=428550 $D=103
M209 5324 272 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=429040 $D=103
M210 4857 273 5325 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=431950 $D=103
M211 5326 274 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=432440 $D=103
M212 4857 275 5327 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=435350 $D=103
M213 5328 276 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=435840 $D=103
M214 4857 277 5329 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=438750 $D=103
M215 5330 278 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=439240 $D=103
M216 4857 279 5331 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=442150 $D=103
M217 5332 280 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=442640 $D=103
M218 4857 281 5333 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=445550 $D=103
M219 5334 282 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=446040 $D=103
M220 4857 283 5335 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=448950 $D=103
M221 5336 284 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=449440 $D=103
M222 4857 285 5337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=452350 $D=103
M223 5338 286 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=452840 $D=103
M224 4857 287 5339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=455750 $D=103
M225 5340 288 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=456240 $D=103
M226 4857 289 5341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=459150 $D=103
M227 5342 290 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=459640 $D=103
M228 4857 291 5343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=462550 $D=103
M229 5344 292 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=463040 $D=103
M230 4857 293 5345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=465950 $D=103
M231 5346 294 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=466440 $D=103
M232 4857 295 5347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=469350 $D=103
M233 5348 296 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=469840 $D=103
M234 4857 297 5349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=472750 $D=103
M235 5350 298 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=473240 $D=103
M236 4857 299 5351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=476150 $D=103
M237 5352 300 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=476640 $D=103
M238 4857 301 5353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=479550 $D=103
M239 5354 302 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=480040 $D=103
M240 4857 303 5355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=482950 $D=103
M241 5356 304 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=483440 $D=103
M242 4857 305 5357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=486350 $D=103
M243 5358 306 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=486840 $D=103
M244 4857 307 5359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=489750 $D=103
M245 5360 308 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=490240 $D=103
M246 4857 309 5361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=493150 $D=103
M247 5362 310 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=493640 $D=103
M248 4857 311 5363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=496550 $D=103
M249 5364 312 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=497040 $D=103
M250 4857 313 5365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=499950 $D=103
M251 5366 314 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=500440 $D=103
M252 4857 315 5367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=503350 $D=103
M253 5368 316 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=503840 $D=103
M254 4857 317 5369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=506750 $D=103
M255 5370 318 4857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=507240 $D=103
M256 341 VSS 3333 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=511190 $D=103
M257 3336 VSS 341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=12500 $Y=511680 $D=103
M258 342 VSS 3334 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13360 $Y=511190 $D=103
M259 3335 VSS 342 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13360 $Y=511680 $D=103
M260 467 VSS 3590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13700 $Y=511190 $D=103
M261 3591 VSS 467 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=13700 $Y=511680 $D=103
M262 468 VSS 3589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14560 $Y=511190 $D=103
M263 3592 VSS 468 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14560 $Y=511680 $D=103
M264 593 VSS 4353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14900 $Y=511190 $D=103
M265 4356 VSS 593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=14900 $Y=511680 $D=103
M266 594 VSS 4354 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15760 $Y=511190 $D=103
M267 4355 VSS 594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=15760 $Y=511680 $D=103
M268 719 VSS 4606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16100 $Y=511190 $D=103
M269 4607 VSS 719 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16100 $Y=511680 $D=103
M270 720 VSS 4605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16960 $Y=511190 $D=103
M271 4608 VSS 720 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=16960 $Y=511680 $D=103
M272 343 VSS 3337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17300 $Y=511190 $D=103
M273 3340 VSS 343 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=17300 $Y=511680 $D=103
M274 344 VSS 3338 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18160 $Y=511190 $D=103
M275 3339 VSS 344 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18160 $Y=511680 $D=103
M276 469 VSS 3594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18500 $Y=511190 $D=103
M277 3595 VSS 469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=18500 $Y=511680 $D=103
M278 470 VSS 3593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19360 $Y=511190 $D=103
M279 3596 VSS 470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19360 $Y=511680 $D=103
M280 595 VSS 4357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19700 $Y=511190 $D=103
M281 4360 VSS 595 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=19700 $Y=511680 $D=103
M282 596 VSS 4358 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=20560 $Y=511190 $D=103
M283 4359 VSS 596 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=20560 $Y=511680 $D=103
M284 721 VSS 4610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=20900 $Y=511190 $D=103
M285 4611 VSS 721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=20900 $Y=511680 $D=103
M286 722 VSS 4609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=21760 $Y=511190 $D=103
M287 4612 VSS 722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=21760 $Y=511680 $D=103
M288 345 VSS 3341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=22100 $Y=511190 $D=103
M289 3344 VSS 345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=22100 $Y=511680 $D=103
M290 346 VSS 3342 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=22960 $Y=511190 $D=103
M291 3343 VSS 346 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=22960 $Y=511680 $D=103
M292 471 VSS 3598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=23300 $Y=511190 $D=103
M293 3599 VSS 471 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=23300 $Y=511680 $D=103
M294 472 VSS 3597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=24160 $Y=511190 $D=103
M295 3600 VSS 472 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=24160 $Y=511680 $D=103
M296 597 VSS 4361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=24500 $Y=511190 $D=103
M297 4364 VSS 597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=24500 $Y=511680 $D=103
M298 598 VSS 4362 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=25360 $Y=511190 $D=103
M299 4363 VSS 598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=25360 $Y=511680 $D=103
M300 723 VSS 4614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=25700 $Y=511190 $D=103
M301 4615 VSS 723 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=25700 $Y=511680 $D=103
M302 724 VSS 4613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=26560 $Y=511190 $D=103
M303 4616 VSS 724 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=26560 $Y=511680 $D=103
M304 347 VSS 3345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=26900 $Y=511190 $D=103
M305 3348 VSS 347 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=26900 $Y=511680 $D=103
M306 348 VSS 3346 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=27760 $Y=511190 $D=103
M307 3347 VSS 348 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=27760 $Y=511680 $D=103
M308 473 VSS 3602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=28100 $Y=511190 $D=103
M309 3603 VSS 473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=28100 $Y=511680 $D=103
M310 474 VSS 3601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=28960 $Y=511190 $D=103
M311 3604 VSS 474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=28960 $Y=511680 $D=103
M312 599 VSS 4365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=29300 $Y=511190 $D=103
M313 4368 VSS 599 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=29300 $Y=511680 $D=103
M314 600 VSS 4366 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=30160 $Y=511190 $D=103
M315 4367 VSS 600 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=30160 $Y=511680 $D=103
M316 725 VSS 4618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=30500 $Y=511190 $D=103
M317 4619 VSS 725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=30500 $Y=511680 $D=103
M318 726 VSS 4617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=31360 $Y=511190 $D=103
M319 4620 VSS 726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=31360 $Y=511680 $D=103
M320 349 VSS 3349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=31700 $Y=511190 $D=103
M321 3352 VSS 349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=31700 $Y=511680 $D=103
M322 350 VSS 3350 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=32560 $Y=511190 $D=103
M323 3351 VSS 350 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=32560 $Y=511680 $D=103
M324 475 VSS 3606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=32900 $Y=511190 $D=103
M325 3607 VSS 475 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=32900 $Y=511680 $D=103
M326 476 VSS 3605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=33760 $Y=511190 $D=103
M327 3608 VSS 476 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=33760 $Y=511680 $D=103
M328 601 VSS 4369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=34100 $Y=511190 $D=103
M329 4372 VSS 601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=34100 $Y=511680 $D=103
M330 602 VSS 4370 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=34960 $Y=511190 $D=103
M331 4371 VSS 602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=34960 $Y=511680 $D=103
M332 727 VSS 4622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=35300 $Y=511190 $D=103
M333 4623 VSS 727 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=35300 $Y=511680 $D=103
M334 728 VSS 4621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=36160 $Y=511190 $D=103
M335 4624 VSS 728 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=36160 $Y=511680 $D=103
M336 351 VSS 3353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=36500 $Y=511190 $D=103
M337 3356 VSS 351 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=36500 $Y=511680 $D=103
M338 352 VSS 3354 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=37360 $Y=511190 $D=103
M339 3355 VSS 352 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=37360 $Y=511680 $D=103
M340 477 VSS 3610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=37700 $Y=511190 $D=103
M341 3611 VSS 477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=37700 $Y=511680 $D=103
M342 478 VSS 3609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38560 $Y=511190 $D=103
M343 3612 VSS 478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38560 $Y=511680 $D=103
M344 603 VSS 4373 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38900 $Y=511190 $D=103
M345 4376 VSS 603 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=38900 $Y=511680 $D=103
M346 604 VSS 4374 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39760 $Y=511190 $D=103
M347 4375 VSS 604 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=39760 $Y=511680 $D=103
M348 729 VSS 4626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=40100 $Y=511190 $D=103
M349 4627 VSS 729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=40100 $Y=511680 $D=103
M350 730 VSS 4625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=40960 $Y=511190 $D=103
M351 4628 VSS 730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=40960 $Y=511680 $D=103
M352 353 VSS 3357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=41300 $Y=511190 $D=103
M353 3360 VSS 353 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=41300 $Y=511680 $D=103
M354 354 VSS 3358 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=42160 $Y=511190 $D=103
M355 3359 VSS 354 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=42160 $Y=511680 $D=103
M356 479 VSS 3614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=42500 $Y=511190 $D=103
M357 3615 VSS 479 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=42500 $Y=511680 $D=103
M358 480 VSS 3613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=43360 $Y=511190 $D=103
M359 3616 VSS 480 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=43360 $Y=511680 $D=103
M360 605 VSS 4377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=43700 $Y=511190 $D=103
M361 4380 VSS 605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=43700 $Y=511680 $D=103
M362 606 VSS 4378 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=44560 $Y=511190 $D=103
M363 4379 VSS 606 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=44560 $Y=511680 $D=103
M364 731 VSS 4630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=44900 $Y=511190 $D=103
M365 4631 VSS 731 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=44900 $Y=511680 $D=103
M366 732 VSS 4629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=45760 $Y=511190 $D=103
M367 4632 VSS 732 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=45760 $Y=511680 $D=103
M368 355 VSS 3361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=46100 $Y=511190 $D=103
M369 3364 VSS 355 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=46100 $Y=511680 $D=103
M370 356 VSS 3362 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=46960 $Y=511190 $D=103
M371 3363 VSS 356 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=46960 $Y=511680 $D=103
M372 481 VSS 3618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=47300 $Y=511190 $D=103
M373 3619 VSS 481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=47300 $Y=511680 $D=103
M374 482 VSS 3617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=48160 $Y=511190 $D=103
M375 3620 VSS 482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=48160 $Y=511680 $D=103
M376 607 VSS 4381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=48500 $Y=511190 $D=103
M377 4384 VSS 607 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=48500 $Y=511680 $D=103
M378 608 VSS 4382 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=49360 $Y=511190 $D=103
M379 4383 VSS 608 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=49360 $Y=511680 $D=103
M380 733 VSS 4634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=49700 $Y=511190 $D=103
M381 4635 VSS 733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=49700 $Y=511680 $D=103
M382 734 VSS 4633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=50560 $Y=511190 $D=103
M383 4636 VSS 734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=50560 $Y=511680 $D=103
M384 357 VSS 3365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=52100 $Y=511190 $D=103
M385 3368 VSS 357 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=52100 $Y=511680 $D=103
M386 358 VSS 3366 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=52960 $Y=511190 $D=103
M387 3367 VSS 358 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=52960 $Y=511680 $D=103
M388 483 VSS 3622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=53300 $Y=511190 $D=103
M389 3623 VSS 483 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=53300 $Y=511680 $D=103
M390 484 VSS 3621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=54160 $Y=511190 $D=103
M391 3624 VSS 484 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=54160 $Y=511680 $D=103
M392 609 VSS 4385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=54500 $Y=511190 $D=103
M393 4388 VSS 609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=54500 $Y=511680 $D=103
M394 610 VSS 4386 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=55360 $Y=511190 $D=103
M395 4387 VSS 610 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=55360 $Y=511680 $D=103
M396 735 VSS 4638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=55700 $Y=511190 $D=103
M397 4639 VSS 735 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=55700 $Y=511680 $D=103
M398 736 VSS 4637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=56560 $Y=511190 $D=103
M399 4640 VSS 736 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=56560 $Y=511680 $D=103
M400 359 VSS 3369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=56900 $Y=511190 $D=103
M401 3372 VSS 359 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=56900 $Y=511680 $D=103
M402 360 VSS 3370 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=57760 $Y=511190 $D=103
M403 3371 VSS 360 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=57760 $Y=511680 $D=103
M404 485 VSS 3626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58100 $Y=511190 $D=103
M405 3627 VSS 485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58100 $Y=511680 $D=103
M406 486 VSS 3625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58960 $Y=511190 $D=103
M407 3628 VSS 486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=58960 $Y=511680 $D=103
M408 611 VSS 4389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=59300 $Y=511190 $D=103
M409 4392 VSS 611 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=59300 $Y=511680 $D=103
M410 612 VSS 4390 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=60160 $Y=511190 $D=103
M411 4391 VSS 612 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=60160 $Y=511680 $D=103
M412 737 VSS 4642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=60500 $Y=511190 $D=103
M413 4643 VSS 737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=60500 $Y=511680 $D=103
M414 738 VSS 4641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=61360 $Y=511190 $D=103
M415 4644 VSS 738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=61360 $Y=511680 $D=103
M416 361 VSS 3373 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=61700 $Y=511190 $D=103
M417 3376 VSS 361 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=61700 $Y=511680 $D=103
M418 362 VSS 3374 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=62560 $Y=511190 $D=103
M419 3375 VSS 362 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=62560 $Y=511680 $D=103
M420 487 VSS 3630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=62900 $Y=511190 $D=103
M421 3631 VSS 487 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=62900 $Y=511680 $D=103
M422 488 VSS 3629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=63760 $Y=511190 $D=103
M423 3632 VSS 488 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=63760 $Y=511680 $D=103
M424 613 VSS 4393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=64100 $Y=511190 $D=103
M425 4396 VSS 613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=64100 $Y=511680 $D=103
M426 614 VSS 4394 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=64960 $Y=511190 $D=103
M427 4395 VSS 614 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=64960 $Y=511680 $D=103
M428 739 VSS 4646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=65300 $Y=511190 $D=103
M429 4647 VSS 739 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=65300 $Y=511680 $D=103
M430 740 VSS 4645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=66160 $Y=511190 $D=103
M431 4648 VSS 740 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=66160 $Y=511680 $D=103
M432 363 VSS 3377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=66500 $Y=511190 $D=103
M433 3380 VSS 363 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=66500 $Y=511680 $D=103
M434 364 VSS 3378 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=67360 $Y=511190 $D=103
M435 3379 VSS 364 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=67360 $Y=511680 $D=103
M436 489 VSS 3634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=67700 $Y=511190 $D=103
M437 3635 VSS 489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=67700 $Y=511680 $D=103
M438 490 VSS 3633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=68560 $Y=511190 $D=103
M439 3636 VSS 490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=68560 $Y=511680 $D=103
M440 615 VSS 4397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=68900 $Y=511190 $D=103
M441 4400 VSS 615 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=68900 $Y=511680 $D=103
M442 616 VSS 4398 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=69760 $Y=511190 $D=103
M443 4399 VSS 616 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=69760 $Y=511680 $D=103
M444 741 VSS 4650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=70100 $Y=511190 $D=103
M445 4651 VSS 741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=70100 $Y=511680 $D=103
M446 742 VSS 4649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=70960 $Y=511190 $D=103
M447 4652 VSS 742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=70960 $Y=511680 $D=103
M448 365 VSS 3381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=71300 $Y=511190 $D=103
M449 3384 VSS 365 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=71300 $Y=511680 $D=103
M450 366 VSS 3382 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=72160 $Y=511190 $D=103
M451 3383 VSS 366 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=72160 $Y=511680 $D=103
M452 491 VSS 3638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=72500 $Y=511190 $D=103
M453 3639 VSS 491 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=72500 $Y=511680 $D=103
M454 492 VSS 3637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=73360 $Y=511190 $D=103
M455 3640 VSS 492 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=73360 $Y=511680 $D=103
M456 617 VSS 4401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=73700 $Y=511190 $D=103
M457 4404 VSS 617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=73700 $Y=511680 $D=103
M458 618 VSS 4402 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=74560 $Y=511190 $D=103
M459 4403 VSS 618 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=74560 $Y=511680 $D=103
M460 743 VSS 4654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=74900 $Y=511190 $D=103
M461 4655 VSS 743 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=74900 $Y=511680 $D=103
M462 744 VSS 4653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=75760 $Y=511190 $D=103
M463 4656 VSS 744 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=75760 $Y=511680 $D=103
M464 367 VSS 3385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=76100 $Y=511190 $D=103
M465 3388 VSS 367 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=76100 $Y=511680 $D=103
M466 368 VSS 3386 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=76960 $Y=511190 $D=103
M467 3387 VSS 368 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=76960 $Y=511680 $D=103
M468 493 VSS 3642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77300 $Y=511190 $D=103
M469 3643 VSS 493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=77300 $Y=511680 $D=103
M470 494 VSS 3641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=78160 $Y=511190 $D=103
M471 3644 VSS 494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=78160 $Y=511680 $D=103
M472 619 VSS 4405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=78500 $Y=511190 $D=103
M473 4408 VSS 619 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=78500 $Y=511680 $D=103
M474 620 VSS 4406 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79360 $Y=511190 $D=103
M475 4407 VSS 620 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79360 $Y=511680 $D=103
M476 745 VSS 4658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79700 $Y=511190 $D=103
M477 4659 VSS 745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=79700 $Y=511680 $D=103
M478 746 VSS 4657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=80560 $Y=511190 $D=103
M479 4660 VSS 746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=80560 $Y=511680 $D=103
M480 369 VSS 3389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=80900 $Y=511190 $D=103
M481 3392 VSS 369 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=80900 $Y=511680 $D=103
M482 370 VSS 3390 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=81760 $Y=511190 $D=103
M483 3391 VSS 370 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=81760 $Y=511680 $D=103
M484 495 VSS 3646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=82100 $Y=511190 $D=103
M485 3647 VSS 495 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=82100 $Y=511680 $D=103
M486 496 VSS 3645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=82960 $Y=511190 $D=103
M487 3648 VSS 496 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=82960 $Y=511680 $D=103
M488 621 VSS 4409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=83300 $Y=511190 $D=103
M489 4412 VSS 621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=83300 $Y=511680 $D=103
M490 622 VSS 4410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=84160 $Y=511190 $D=103
M491 4411 VSS 622 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=84160 $Y=511680 $D=103
M492 747 VSS 4662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=84500 $Y=511190 $D=103
M493 4663 VSS 747 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=84500 $Y=511680 $D=103
M494 748 VSS 4661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=85360 $Y=511190 $D=103
M495 4664 VSS 748 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=85360 $Y=511680 $D=103
M496 371 VSS 3393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=85700 $Y=511190 $D=103
M497 3396 VSS 371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=85700 $Y=511680 $D=103
M498 372 VSS 3394 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=86560 $Y=511190 $D=103
M499 3395 VSS 372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=86560 $Y=511680 $D=103
M500 497 VSS 3650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=86900 $Y=511190 $D=103
M501 3651 VSS 497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=86900 $Y=511680 $D=103
M502 498 VSS 3649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=87760 $Y=511190 $D=103
M503 3652 VSS 498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=87760 $Y=511680 $D=103
M504 319 VSS 3329 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=88100 $Y=511190 $D=103
M505 3332 VSS 319 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=88100 $Y=511680 $D=103
M506 320 VSS 3330 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=88960 $Y=511190 $D=103
M507 3331 VSS 320 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=88960 $Y=511680 $D=103
M508 321 VSS 5372 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=89300 $Y=511190 $D=103
M509 5373 VSS 321 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=89300 $Y=511680 $D=103
M510 322 50 5371 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=90160 $Y=511190 $D=103
M511 5374 50 322 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=90160 $Y=511680 $D=103
M512 373 50 3397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=91700 $Y=511190 $D=103
M513 3400 50 373 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=91700 $Y=511680 $D=103
M514 374 50 3398 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=92560 $Y=511190 $D=103
M515 3399 50 374 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=92560 $Y=511680 $D=103
M516 499 50 3654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=92900 $Y=511190 $D=103
M517 3655 50 499 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=92900 $Y=511680 $D=103
M518 500 50 3653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=93760 $Y=511190 $D=103
M519 3656 50 500 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=93760 $Y=511680 $D=103
M520 623 50 4413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=94100 $Y=511190 $D=103
M521 4416 50 623 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=94100 $Y=511680 $D=103
M522 624 50 4414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=94960 $Y=511190 $D=103
M523 4415 50 624 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=94960 $Y=511680 $D=103
M524 749 50 4666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=95300 $Y=511190 $D=103
M525 4667 50 749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=95300 $Y=511680 $D=103
M526 750 50 4665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=96160 $Y=511190 $D=103
M527 4668 50 750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=96160 $Y=511680 $D=103
M528 375 50 3401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=96500 $Y=511190 $D=103
M529 3404 50 375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=96500 $Y=511680 $D=103
M530 376 50 3402 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=97360 $Y=511190 $D=103
M531 3403 50 376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=97360 $Y=511680 $D=103
M532 501 50 3658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=97700 $Y=511190 $D=103
M533 3659 50 501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=97700 $Y=511680 $D=103
M534 502 50 3657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98560 $Y=511190 $D=103
M535 3660 50 502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98560 $Y=511680 $D=103
M536 625 50 4417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98900 $Y=511190 $D=103
M537 4420 50 625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=98900 $Y=511680 $D=103
M538 626 50 4418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=99760 $Y=511190 $D=103
M539 4419 50 626 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=99760 $Y=511680 $D=103
M540 751 50 4670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=100100 $Y=511190 $D=103
M541 4671 50 751 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=100100 $Y=511680 $D=103
M542 752 50 4669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=100960 $Y=511190 $D=103
M543 4672 50 752 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=100960 $Y=511680 $D=103
M544 377 50 3405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=101300 $Y=511190 $D=103
M545 3408 50 377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=101300 $Y=511680 $D=103
M546 378 50 3406 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=102160 $Y=511190 $D=103
M547 3407 50 378 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=102160 $Y=511680 $D=103
M548 503 50 3662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=102500 $Y=511190 $D=103
M549 3663 50 503 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=102500 $Y=511680 $D=103
M550 504 50 3661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=103360 $Y=511190 $D=103
M551 3664 50 504 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=103360 $Y=511680 $D=103
M552 627 50 4421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=103700 $Y=511190 $D=103
M553 4424 50 627 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=103700 $Y=511680 $D=103
M554 628 50 4422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=104560 $Y=511190 $D=103
M555 4423 50 628 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=104560 $Y=511680 $D=103
M556 753 50 4674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=104900 $Y=511190 $D=103
M557 4675 50 753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=104900 $Y=511680 $D=103
M558 754 50 4673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=105760 $Y=511190 $D=103
M559 4676 50 754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=105760 $Y=511680 $D=103
M560 379 50 3409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=106100 $Y=511190 $D=103
M561 3412 50 379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=106100 $Y=511680 $D=103
M562 380 50 3410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=106960 $Y=511190 $D=103
M563 3411 50 380 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=106960 $Y=511680 $D=103
M564 505 50 3666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=107300 $Y=511190 $D=103
M565 3667 50 505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=107300 $Y=511680 $D=103
M566 506 50 3665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=108160 $Y=511190 $D=103
M567 3668 50 506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=108160 $Y=511680 $D=103
M568 629 50 4425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=108500 $Y=511190 $D=103
M569 4428 50 629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=108500 $Y=511680 $D=103
M570 630 50 4426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=109360 $Y=511190 $D=103
M571 4427 50 630 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=109360 $Y=511680 $D=103
M572 755 50 4678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=109700 $Y=511190 $D=103
M573 4679 50 755 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=109700 $Y=511680 $D=103
M574 756 50 4677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=110560 $Y=511190 $D=103
M575 4680 50 756 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=110560 $Y=511680 $D=103
M576 381 50 3413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=110900 $Y=511190 $D=103
M577 3416 50 381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=110900 $Y=511680 $D=103
M578 382 50 3414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=111760 $Y=511190 $D=103
M579 3415 50 382 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=111760 $Y=511680 $D=103
M580 507 50 3670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=112100 $Y=511190 $D=103
M581 3671 50 507 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=112100 $Y=511680 $D=103
M582 508 50 3669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=112960 $Y=511190 $D=103
M583 3672 50 508 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=112960 $Y=511680 $D=103
M584 631 50 4429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=113300 $Y=511190 $D=103
M585 4432 50 631 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=113300 $Y=511680 $D=103
M586 632 50 4430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=114160 $Y=511190 $D=103
M587 4431 50 632 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=114160 $Y=511680 $D=103
M588 757 50 4682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=114500 $Y=511190 $D=103
M589 4683 50 757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=114500 $Y=511680 $D=103
M590 758 50 4681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=115360 $Y=511190 $D=103
M591 4684 50 758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=115360 $Y=511680 $D=103
M592 383 50 3417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=115700 $Y=511190 $D=103
M593 3420 50 383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=115700 $Y=511680 $D=103
M594 384 50 3418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=116560 $Y=511190 $D=103
M595 3419 50 384 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=116560 $Y=511680 $D=103
M596 509 50 3674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=116900 $Y=511190 $D=103
M597 3675 50 509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=116900 $Y=511680 $D=103
M598 510 50 3673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117760 $Y=511190 $D=103
M599 3676 50 510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=117760 $Y=511680 $D=103
M600 633 50 4433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118100 $Y=511190 $D=103
M601 4436 50 633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118100 $Y=511680 $D=103
M602 634 50 4434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118960 $Y=511190 $D=103
M603 4435 50 634 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=118960 $Y=511680 $D=103
M604 759 50 4686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=119300 $Y=511190 $D=103
M605 4687 50 759 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=119300 $Y=511680 $D=103
M606 760 50 4685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=120160 $Y=511190 $D=103
M607 4688 50 760 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=120160 $Y=511680 $D=103
M608 385 50 3421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=120500 $Y=511190 $D=103
M609 3424 50 385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=120500 $Y=511680 $D=103
M610 386 50 3422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=121360 $Y=511190 $D=103
M611 3423 50 386 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=121360 $Y=511680 $D=103
M612 511 50 3678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=121700 $Y=511190 $D=103
M613 3679 50 511 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=121700 $Y=511680 $D=103
M614 512 50 3677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=122560 $Y=511190 $D=103
M615 3680 50 512 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=122560 $Y=511680 $D=103
M616 635 50 4437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=122900 $Y=511190 $D=103
M617 4440 50 635 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=122900 $Y=511680 $D=103
M618 636 50 4438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=123760 $Y=511190 $D=103
M619 4439 50 636 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=123760 $Y=511680 $D=103
M620 761 50 4690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=124100 $Y=511190 $D=103
M621 4691 50 761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=124100 $Y=511680 $D=103
M622 762 50 4689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=124960 $Y=511190 $D=103
M623 4692 50 762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=124960 $Y=511680 $D=103
M624 387 50 3425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=125300 $Y=511190 $D=103
M625 3428 50 387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=125300 $Y=511680 $D=103
M626 388 50 3426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=126160 $Y=511190 $D=103
M627 3427 50 388 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=126160 $Y=511680 $D=103
M628 513 50 3682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=126500 $Y=511190 $D=103
M629 3683 50 513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=126500 $Y=511680 $D=103
M630 514 50 3681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=127360 $Y=511190 $D=103
M631 3684 50 514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=127360 $Y=511680 $D=103
M632 637 50 4441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=127700 $Y=511190 $D=103
M633 4444 50 637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=127700 $Y=511680 $D=103
M634 638 50 4442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=128560 $Y=511190 $D=103
M635 4443 50 638 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=128560 $Y=511680 $D=103
M636 763 50 4694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=128900 $Y=511190 $D=103
M637 4695 50 763 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=128900 $Y=511680 $D=103
M638 764 50 4693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=129760 $Y=511190 $D=103
M639 4696 50 764 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=129760 $Y=511680 $D=103
M640 389 50 3429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=131300 $Y=511190 $D=103
M641 3432 50 389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=131300 $Y=511680 $D=103
M642 390 50 3430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=132160 $Y=511190 $D=103
M643 3431 50 390 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=132160 $Y=511680 $D=103
M644 515 50 3686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=132500 $Y=511190 $D=103
M645 3687 50 515 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=132500 $Y=511680 $D=103
M646 516 50 3685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=133360 $Y=511190 $D=103
M647 3688 50 516 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=133360 $Y=511680 $D=103
M648 639 50 4445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=133700 $Y=511190 $D=103
M649 4448 50 639 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=133700 $Y=511680 $D=103
M650 640 50 4446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=134560 $Y=511190 $D=103
M651 4447 50 640 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=134560 $Y=511680 $D=103
M652 765 50 4698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=134900 $Y=511190 $D=103
M653 4699 50 765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=134900 $Y=511680 $D=103
M654 766 50 4697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=135760 $Y=511190 $D=103
M655 4700 50 766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=135760 $Y=511680 $D=103
M656 391 50 3433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=136100 $Y=511190 $D=103
M657 3436 50 391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=136100 $Y=511680 $D=103
M658 392 50 3434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=136960 $Y=511190 $D=103
M659 3435 50 392 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=136960 $Y=511680 $D=103
M660 517 50 3690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137300 $Y=511190 $D=103
M661 3691 50 517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=137300 $Y=511680 $D=103
M662 518 50 3689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138160 $Y=511190 $D=103
M663 3692 50 518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138160 $Y=511680 $D=103
M664 641 50 4449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138500 $Y=511190 $D=103
M665 4452 50 641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=138500 $Y=511680 $D=103
M666 642 50 4450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=139360 $Y=511190 $D=103
M667 4451 50 642 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=139360 $Y=511680 $D=103
M668 767 50 4702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=139700 $Y=511190 $D=103
M669 4703 50 767 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=139700 $Y=511680 $D=103
M670 768 50 4701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=140560 $Y=511190 $D=103
M671 4704 50 768 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=140560 $Y=511680 $D=103
M672 393 50 3437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=140900 $Y=511190 $D=103
M673 3440 50 393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=140900 $Y=511680 $D=103
M674 394 50 3438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=141760 $Y=511190 $D=103
M675 3439 50 394 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=141760 $Y=511680 $D=103
M676 519 50 3694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=142100 $Y=511190 $D=103
M677 3695 50 519 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=142100 $Y=511680 $D=103
M678 520 50 3693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=142960 $Y=511190 $D=103
M679 3696 50 520 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=142960 $Y=511680 $D=103
M680 643 50 4453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=143300 $Y=511190 $D=103
M681 4456 50 643 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=143300 $Y=511680 $D=103
M682 644 50 4454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=144160 $Y=511190 $D=103
M683 4455 50 644 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=144160 $Y=511680 $D=103
M684 769 50 4706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=144500 $Y=511190 $D=103
M685 4707 50 769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=144500 $Y=511680 $D=103
M686 770 50 4705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=145360 $Y=511190 $D=103
M687 4708 50 770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=145360 $Y=511680 $D=103
M688 395 50 3441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=145700 $Y=511190 $D=103
M689 3444 50 395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=145700 $Y=511680 $D=103
M690 396 50 3442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=146560 $Y=511190 $D=103
M691 3443 50 396 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=146560 $Y=511680 $D=103
M692 521 50 3698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=146900 $Y=511190 $D=103
M693 3699 50 521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=146900 $Y=511680 $D=103
M694 522 50 3697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=147760 $Y=511190 $D=103
M695 3700 50 522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=147760 $Y=511680 $D=103
M696 645 50 4457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=148100 $Y=511190 $D=103
M697 4460 50 645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=148100 $Y=511680 $D=103
M698 646 50 4458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=148960 $Y=511190 $D=103
M699 4459 50 646 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=148960 $Y=511680 $D=103
M700 771 50 4710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=149300 $Y=511190 $D=103
M701 4711 50 771 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=149300 $Y=511680 $D=103
M702 772 50 4709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=150160 $Y=511190 $D=103
M703 4712 50 772 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=150160 $Y=511680 $D=103
M704 397 50 3445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=150500 $Y=511190 $D=103
M705 3448 50 397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=150500 $Y=511680 $D=103
M706 398 50 3446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=151360 $Y=511190 $D=103
M707 3447 50 398 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=151360 $Y=511680 $D=103
M708 523 50 3702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=151700 $Y=511190 $D=103
M709 3703 50 523 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=151700 $Y=511680 $D=103
M710 524 50 3701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=152560 $Y=511190 $D=103
M711 3704 50 524 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=152560 $Y=511680 $D=103
M712 647 50 4461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=152900 $Y=511190 $D=103
M713 4464 50 647 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=152900 $Y=511680 $D=103
M714 648 50 4462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=153760 $Y=511190 $D=103
M715 4463 50 648 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=153760 $Y=511680 $D=103
M716 773 50 4714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=154100 $Y=511190 $D=103
M717 4715 50 773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=154100 $Y=511680 $D=103
M718 774 50 4713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=154960 $Y=511190 $D=103
M719 4716 50 774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=154960 $Y=511680 $D=103
M720 399 50 3449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=155300 $Y=511190 $D=103
M721 3452 50 399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=155300 $Y=511680 $D=103
M722 400 50 3450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=156160 $Y=511190 $D=103
M723 3451 50 400 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=156160 $Y=511680 $D=103
M724 525 50 3706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=156500 $Y=511190 $D=103
M725 3707 50 525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=156500 $Y=511680 $D=103
M726 526 50 3705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=157360 $Y=511190 $D=103
M727 3708 50 526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=157360 $Y=511680 $D=103
M728 649 50 4465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=157700 $Y=511190 $D=103
M729 4468 50 649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=157700 $Y=511680 $D=103
M730 650 50 4466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=158560 $Y=511190 $D=103
M731 4467 50 650 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=158560 $Y=511680 $D=103
M732 775 50 4718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=158900 $Y=511190 $D=103
M733 4719 50 775 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=158900 $Y=511680 $D=103
M734 776 50 4717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=159760 $Y=511190 $D=103
M735 4720 50 776 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=159760 $Y=511680 $D=103
M736 401 50 3453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=160100 $Y=511190 $D=103
M737 3456 50 401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=160100 $Y=511680 $D=103
M738 402 50 3454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=160960 $Y=511190 $D=103
M739 3455 50 402 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=160960 $Y=511680 $D=103
M740 527 50 3710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=161300 $Y=511190 $D=103
M741 3711 50 527 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=161300 $Y=511680 $D=103
M742 528 50 3709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=162160 $Y=511190 $D=103
M743 3712 50 528 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=162160 $Y=511680 $D=103
M744 651 50 4469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=162500 $Y=511190 $D=103
M745 4472 50 651 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=162500 $Y=511680 $D=103
M746 652 50 4470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=163360 $Y=511190 $D=103
M747 4471 50 652 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=163360 $Y=511680 $D=103
M748 777 50 4722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=163700 $Y=511190 $D=103
M749 4723 50 777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=163700 $Y=511680 $D=103
M750 778 50 4721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=164560 $Y=511190 $D=103
M751 4724 50 778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=164560 $Y=511680 $D=103
M752 403 50 3457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=164900 $Y=511190 $D=103
M753 3460 50 403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=164900 $Y=511680 $D=103
M754 404 50 3458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=165760 $Y=511190 $D=103
M755 3459 50 404 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=165760 $Y=511680 $D=103
M756 529 50 3714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=166100 $Y=511190 $D=103
M757 3715 50 529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=166100 $Y=511680 $D=103
M758 530 50 3713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=166960 $Y=511190 $D=103
M759 3716 50 530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=166960 $Y=511680 $D=103
M760 653 50 4473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=167300 $Y=511190 $D=103
M761 4476 50 653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=167300 $Y=511680 $D=103
M762 654 50 4474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=168160 $Y=511190 $D=103
M763 4475 50 654 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=168160 $Y=511680 $D=103
M764 779 50 4726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=168500 $Y=511190 $D=103
M765 4727 50 779 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=168500 $Y=511680 $D=103
M766 4858 63 4859 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=74950 $D=103
M767 4860 64 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=75440 $D=103
M768 4858 65 4861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=78350 $D=103
M769 4862 66 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=78840 $D=103
M770 4858 67 4863 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=81750 $D=103
M771 4864 68 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=82240 $D=103
M772 4858 69 4865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=85150 $D=103
M773 4866 70 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=85640 $D=103
M774 4858 71 4867 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=88550 $D=103
M775 4868 72 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=89040 $D=103
M776 4858 73 4869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=91950 $D=103
M777 4870 74 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=92440 $D=103
M778 4858 75 4871 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=95350 $D=103
M779 4872 76 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=95840 $D=103
M780 4858 77 4873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=98750 $D=103
M781 4874 78 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=99240 $D=103
M782 4858 79 4875 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=102150 $D=103
M783 4876 80 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=102640 $D=103
M784 4858 81 4877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=105550 $D=103
M785 4878 82 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=106040 $D=103
M786 4858 83 4879 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=108950 $D=103
M787 4880 84 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=109440 $D=103
M788 4858 85 4881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=112350 $D=103
M789 4882 86 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=112840 $D=103
M790 4858 87 4883 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=115750 $D=103
M791 4884 88 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=116240 $D=103
M792 4858 89 4885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=119150 $D=103
M793 4886 90 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=119640 $D=103
M794 4858 91 4887 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=122550 $D=103
M795 4888 92 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=123040 $D=103
M796 4858 93 4889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=125950 $D=103
M797 4890 94 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=126440 $D=103
M798 4858 95 4891 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=129350 $D=103
M799 4892 96 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=129840 $D=103
M800 4858 97 4893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=132750 $D=103
M801 4894 98 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=133240 $D=103
M802 4858 99 4895 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=136150 $D=103
M803 4896 100 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=136640 $D=103
M804 4858 101 4897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=139550 $D=103
M805 4898 102 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=140040 $D=103
M806 4858 103 4899 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=142950 $D=103
M807 4900 104 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=143440 $D=103
M808 4858 105 4901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=146350 $D=103
M809 4902 106 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=146840 $D=103
M810 4858 107 4903 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=149750 $D=103
M811 4904 108 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=150240 $D=103
M812 4858 109 4905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=153150 $D=103
M813 4906 110 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=153640 $D=103
M814 4858 111 4907 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=156550 $D=103
M815 4908 112 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=157040 $D=103
M816 4858 113 4909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=159950 $D=103
M817 4910 114 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=160440 $D=103
M818 4858 115 4911 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=163350 $D=103
M819 4912 116 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=163840 $D=103
M820 4858 117 4913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=166750 $D=103
M821 4914 118 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=167240 $D=103
M822 4858 119 4915 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=170150 $D=103
M823 4916 120 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=170640 $D=103
M824 4858 121 4917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=173550 $D=103
M825 4918 122 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=174040 $D=103
M826 4858 123 4919 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=176950 $D=103
M827 4920 124 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=177440 $D=103
M828 4858 125 4921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=180350 $D=103
M829 4922 126 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=180840 $D=103
M830 4858 127 4923 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=183750 $D=103
M831 4924 128 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=184240 $D=103
M832 4858 129 4925 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=187150 $D=103
M833 4926 130 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=187640 $D=103
M834 4858 131 4927 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=190550 $D=103
M835 4928 132 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=191040 $D=103
M836 4858 133 4929 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=193950 $D=103
M837 4930 134 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=194440 $D=103
M838 4858 135 4931 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=197350 $D=103
M839 4932 136 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=197840 $D=103
M840 4858 137 4933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=200750 $D=103
M841 4934 138 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=201240 $D=103
M842 4858 139 4935 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=204150 $D=103
M843 4936 140 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=204640 $D=103
M844 4858 141 4937 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=207550 $D=103
M845 4938 142 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=208040 $D=103
M846 4858 143 4939 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=210950 $D=103
M847 4940 144 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=211440 $D=103
M848 4858 145 4941 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=214350 $D=103
M849 4942 146 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=214840 $D=103
M850 4858 147 4943 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=217750 $D=103
M851 4944 148 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=218240 $D=103
M852 4858 149 4945 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=221150 $D=103
M853 4946 150 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=221640 $D=103
M854 4858 151 4947 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=224550 $D=103
M855 4948 152 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=225040 $D=103
M856 4858 153 4949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=227950 $D=103
M857 4950 154 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=228440 $D=103
M858 4858 155 4951 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=231350 $D=103
M859 4952 156 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=231840 $D=103
M860 4858 157 4953 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=234750 $D=103
M861 4954 158 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=235240 $D=103
M862 4858 159 4955 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=238150 $D=103
M863 4956 160 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=238640 $D=103
M864 4858 161 4957 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=241550 $D=103
M865 4958 162 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=242040 $D=103
M866 4858 163 4959 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=244950 $D=103
M867 4960 164 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=245440 $D=103
M868 4858 165 4961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=248350 $D=103
M869 4962 166 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=248840 $D=103
M870 4858 167 4963 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=251750 $D=103
M871 4964 168 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=252240 $D=103
M872 4858 169 4965 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=255150 $D=103
M873 4966 170 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=255640 $D=103
M874 4858 171 4967 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=258550 $D=103
M875 4968 172 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=259040 $D=103
M876 4858 173 4969 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=261950 $D=103
M877 4970 174 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=262440 $D=103
M878 4858 175 4971 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=265350 $D=103
M879 4972 176 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=265840 $D=103
M880 4858 177 4973 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=268750 $D=103
M881 4974 178 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=269240 $D=103
M882 4858 179 4975 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=272150 $D=103
M883 4976 180 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=272640 $D=103
M884 4858 181 4977 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=275550 $D=103
M885 4978 182 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=276040 $D=103
M886 4858 183 4979 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=278950 $D=103
M887 4980 184 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=279440 $D=103
M888 4858 185 4981 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=282350 $D=103
M889 4982 186 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=282840 $D=103
M890 4858 187 4983 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=285750 $D=103
M891 4984 188 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=286240 $D=103
M892 4858 189 4985 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=289150 $D=103
M893 4986 190 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=289640 $D=103
M894 4858 191 4987 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=292550 $D=103
M895 4988 192 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=293040 $D=103
M896 4858 193 4989 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=295950 $D=103
M897 4990 194 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=296440 $D=103
M898 4858 195 4991 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=299350 $D=103
M899 4992 196 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=299840 $D=103
M900 4858 197 4993 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=302750 $D=103
M901 4994 198 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=303240 $D=103
M902 4858 199 4995 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=306150 $D=103
M903 4996 200 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=306640 $D=103
M904 4858 201 4997 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=309550 $D=103
M905 4998 202 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=310040 $D=103
M906 4858 203 4999 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=312950 $D=103
M907 5000 204 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=313440 $D=103
M908 4858 205 5001 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=316350 $D=103
M909 5002 206 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=316840 $D=103
M910 4858 207 5003 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=319750 $D=103
M911 5004 208 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=320240 $D=103
M912 4858 209 5005 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=323150 $D=103
M913 5006 210 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=323640 $D=103
M914 4858 211 5007 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=326550 $D=103
M915 5008 212 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=327040 $D=103
M916 4858 213 5009 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=329950 $D=103
M917 5010 214 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=330440 $D=103
M918 4858 215 5011 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=333350 $D=103
M919 5012 216 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=333840 $D=103
M920 4858 217 5013 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=336750 $D=103
M921 5014 218 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=337240 $D=103
M922 4858 219 5015 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=340150 $D=103
M923 5016 220 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=340640 $D=103
M924 4858 221 5017 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=343550 $D=103
M925 5018 222 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=344040 $D=103
M926 4858 223 5019 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=346950 $D=103
M927 5020 224 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=347440 $D=103
M928 4858 225 5021 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=350350 $D=103
M929 5022 226 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=350840 $D=103
M930 4858 227 5023 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=353750 $D=103
M931 5024 228 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=354240 $D=103
M932 4858 229 5025 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=357150 $D=103
M933 5026 230 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=357640 $D=103
M934 4858 231 5027 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=360550 $D=103
M935 5028 232 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=361040 $D=103
M936 4858 233 5029 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=363950 $D=103
M937 5030 234 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=364440 $D=103
M938 4858 235 5031 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=367350 $D=103
M939 5032 236 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=367840 $D=103
M940 4858 237 5033 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=370750 $D=103
M941 5034 238 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=371240 $D=103
M942 4858 239 5035 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=374150 $D=103
M943 5036 240 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=374640 $D=103
M944 4858 241 5037 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=377550 $D=103
M945 5038 242 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=378040 $D=103
M946 4858 243 5039 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=380950 $D=103
M947 5040 244 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=381440 $D=103
M948 4858 245 5041 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=384350 $D=103
M949 5042 246 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=384840 $D=103
M950 4858 247 5043 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=387750 $D=103
M951 5044 248 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=388240 $D=103
M952 4858 249 5045 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=391150 $D=103
M953 5046 250 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=391640 $D=103
M954 4858 251 5047 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=394550 $D=103
M955 5048 252 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=395040 $D=103
M956 4858 253 5049 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=397950 $D=103
M957 5050 254 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=398440 $D=103
M958 4858 255 5051 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=401350 $D=103
M959 5052 256 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=401840 $D=103
M960 4858 257 5053 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=404750 $D=103
M961 5054 258 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=405240 $D=103
M962 4858 259 5055 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=408150 $D=103
M963 5056 260 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=408640 $D=103
M964 4858 261 5057 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=411550 $D=103
M965 5058 262 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=412040 $D=103
M966 4858 263 5059 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=414950 $D=103
M967 5060 264 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=415440 $D=103
M968 4858 265 5061 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=418350 $D=103
M969 5062 266 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=418840 $D=103
M970 4858 267 5063 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=421750 $D=103
M971 5064 268 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=422240 $D=103
M972 4858 269 5065 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=425150 $D=103
M973 5066 270 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=425640 $D=103
M974 4858 271 5067 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=428550 $D=103
M975 5068 272 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=429040 $D=103
M976 4858 273 5069 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=431950 $D=103
M977 5070 274 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=432440 $D=103
M978 4858 275 5071 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=435350 $D=103
M979 5072 276 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=435840 $D=103
M980 4858 277 5073 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=438750 $D=103
M981 5074 278 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=439240 $D=103
M982 4858 279 5075 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=442150 $D=103
M983 5076 280 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=442640 $D=103
M984 4858 281 5077 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=445550 $D=103
M985 5078 282 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=446040 $D=103
M986 4858 283 5079 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=448950 $D=103
M987 5080 284 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=449440 $D=103
M988 4858 285 5081 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=452350 $D=103
M989 5082 286 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=452840 $D=103
M990 4858 287 5083 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=455750 $D=103
M991 5084 288 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=456240 $D=103
M992 4858 289 5085 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=459150 $D=103
M993 5086 290 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=459640 $D=103
M994 4858 291 5087 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=462550 $D=103
M995 5088 292 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=463040 $D=103
M996 4858 293 5089 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=465950 $D=103
M997 5090 294 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=466440 $D=103
M998 4858 295 5091 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=469350 $D=103
M999 5092 296 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=469840 $D=103
M1000 4858 297 5093 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=472750 $D=103
M1001 5094 298 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=473240 $D=103
M1002 4858 299 5095 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=476150 $D=103
M1003 5096 300 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=476640 $D=103
M1004 4858 301 5097 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=479550 $D=103
M1005 5098 302 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=480040 $D=103
M1006 4858 303 5099 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=482950 $D=103
M1007 5100 304 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=483440 $D=103
M1008 4858 305 5101 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=486350 $D=103
M1009 5102 306 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=486840 $D=103
M1010 4858 307 5103 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=489750 $D=103
M1011 5104 308 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=490240 $D=103
M1012 4858 309 5105 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=493150 $D=103
M1013 5106 310 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=493640 $D=103
M1014 4858 311 5107 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=496550 $D=103
M1015 5108 312 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=497040 $D=103
M1016 4858 313 5109 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=499950 $D=103
M1017 5110 314 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=500440 $D=103
M1018 4858 315 5111 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=503350 $D=103
M1019 5112 316 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=503840 $D=103
M1020 4858 317 5113 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=506750 $D=103
M1021 5114 318 4858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=507240 $D=103
M1022 780 50 4725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=511190 $D=103
M1023 4728 50 780 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=169360 $Y=511680 $D=103
M1024 60 VSS 3718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=74950 $D=103
M1025 3719 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=75440 $D=103
M1026 60 VSS 3721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=78350 $D=103
M1027 3724 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=78840 $D=103
M1028 60 VSS 3726 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=81750 $D=103
M1029 3727 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=82240 $D=103
M1030 60 VSS 3729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=85150 $D=103
M1031 3732 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=85640 $D=103
M1032 60 VSS 3734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=88550 $D=103
M1033 3735 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=89040 $D=103
M1034 60 VSS 3737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=91950 $D=103
M1035 3740 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=92440 $D=103
M1036 60 VSS 3742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=95350 $D=103
M1037 3743 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=95840 $D=103
M1038 60 VSS 3745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=98750 $D=103
M1039 3748 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=99240 $D=103
M1040 60 VSS 3750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=102150 $D=103
M1041 3751 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=102640 $D=103
M1042 60 VSS 3753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=105550 $D=103
M1043 3756 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=106040 $D=103
M1044 60 VSS 3758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=108950 $D=103
M1045 3759 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=109440 $D=103
M1046 60 VSS 3761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=112350 $D=103
M1047 3764 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=112840 $D=103
M1048 60 VSS 3766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=115750 $D=103
M1049 3767 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=116240 $D=103
M1050 60 VSS 3769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=119150 $D=103
M1051 3772 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=119640 $D=103
M1052 60 VSS 3774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=122550 $D=103
M1053 3775 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=123040 $D=103
M1054 60 VSS 3777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=125950 $D=103
M1055 3780 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=126440 $D=103
M1056 60 VSS 3782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=129350 $D=103
M1057 3783 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=129840 $D=103
M1058 60 VSS 3785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=132750 $D=103
M1059 3788 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=133240 $D=103
M1060 60 VSS 3790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=136150 $D=103
M1061 3791 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=136640 $D=103
M1062 60 VSS 3793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=139550 $D=103
M1063 3796 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=140040 $D=103
M1064 60 VSS 3798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=142950 $D=103
M1065 3799 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=143440 $D=103
M1066 60 VSS 3801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=146350 $D=103
M1067 3804 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=146840 $D=103
M1068 60 VSS 3806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=149750 $D=103
M1069 3807 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=150240 $D=103
M1070 60 VSS 3809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=153150 $D=103
M1071 3812 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=153640 $D=103
M1072 60 VSS 3814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=156550 $D=103
M1073 3815 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=157040 $D=103
M1074 60 VSS 3817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=159950 $D=103
M1075 3820 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=160440 $D=103
M1076 60 VSS 3822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=163350 $D=103
M1077 3823 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=163840 $D=103
M1078 60 VSS 3825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=166750 $D=103
M1079 3828 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=167240 $D=103
M1080 60 VSS 3830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=170150 $D=103
M1081 3831 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=170640 $D=103
M1082 60 VSS 3833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=173550 $D=103
M1083 3836 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=174040 $D=103
M1084 60 VSS 3838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=176950 $D=103
M1085 3839 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=177440 $D=103
M1086 60 VSS 3841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=180350 $D=103
M1087 3844 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=180840 $D=103
M1088 60 VSS 3846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=183750 $D=103
M1089 3847 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=184240 $D=103
M1090 60 VSS 3849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=187150 $D=103
M1091 3852 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=187640 $D=103
M1092 60 VSS 3854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=190550 $D=103
M1093 3855 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=191040 $D=103
M1094 60 VSS 3857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=193950 $D=103
M1095 3860 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=194440 $D=103
M1096 60 VSS 3862 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=197350 $D=103
M1097 3863 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=197840 $D=103
M1098 60 VSS 3865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=200750 $D=103
M1099 3868 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=201240 $D=103
M1100 60 VSS 3870 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=204150 $D=103
M1101 3871 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=204640 $D=103
M1102 60 VSS 3873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=207550 $D=103
M1103 3876 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=208040 $D=103
M1104 60 VSS 3878 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=210950 $D=103
M1105 3879 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=211440 $D=103
M1106 60 VSS 3881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=214350 $D=103
M1107 3884 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=214840 $D=103
M1108 60 VSS 3886 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=217750 $D=103
M1109 3887 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=218240 $D=103
M1110 60 VSS 3889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=221150 $D=103
M1111 3892 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=221640 $D=103
M1112 60 VSS 3894 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=224550 $D=103
M1113 3895 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=225040 $D=103
M1114 60 VSS 3897 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=227950 $D=103
M1115 3900 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=228440 $D=103
M1116 60 VSS 3902 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=231350 $D=103
M1117 3903 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=231840 $D=103
M1118 60 VSS 3905 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=234750 $D=103
M1119 3908 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=235240 $D=103
M1120 60 VSS 3910 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=238150 $D=103
M1121 3911 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=238640 $D=103
M1122 60 VSS 3913 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=241550 $D=103
M1123 3916 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=242040 $D=103
M1124 60 VSS 3918 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=244950 $D=103
M1125 3919 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=245440 $D=103
M1126 60 VSS 3921 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=248350 $D=103
M1127 3924 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=248840 $D=103
M1128 60 VSS 3926 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=251750 $D=103
M1129 3927 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=252240 $D=103
M1130 60 VSS 3929 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=255150 $D=103
M1131 3932 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=255640 $D=103
M1132 60 VSS 3934 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=258550 $D=103
M1133 3935 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=259040 $D=103
M1134 60 VSS 3937 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=261950 $D=103
M1135 3940 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=262440 $D=103
M1136 60 VSS 3942 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=265350 $D=103
M1137 3943 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=265840 $D=103
M1138 60 VSS 3945 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=268750 $D=103
M1139 3948 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=269240 $D=103
M1140 60 VSS 3950 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=272150 $D=103
M1141 3951 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=272640 $D=103
M1142 60 VSS 3953 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=275550 $D=103
M1143 3956 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=276040 $D=103
M1144 60 VSS 3958 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=278950 $D=103
M1145 3959 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=279440 $D=103
M1146 60 VSS 3961 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=282350 $D=103
M1147 3964 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=282840 $D=103
M1148 60 VSS 3966 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=285750 $D=103
M1149 3967 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=286240 $D=103
M1150 60 VSS 3969 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=289150 $D=103
M1151 3972 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=289640 $D=103
M1152 60 VSS 3974 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=292550 $D=103
M1153 3975 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=293040 $D=103
M1154 60 VSS 3977 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=295950 $D=103
M1155 3980 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=296440 $D=103
M1156 60 VSS 3982 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=299350 $D=103
M1157 3983 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=299840 $D=103
M1158 60 VSS 3985 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=302750 $D=103
M1159 3988 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=303240 $D=103
M1160 60 VSS 3990 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=306150 $D=103
M1161 3991 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=306640 $D=103
M1162 60 VSS 3993 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=309550 $D=103
M1163 3996 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=310040 $D=103
M1164 60 VSS 3998 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=312950 $D=103
M1165 3999 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=313440 $D=103
M1166 60 VSS 4001 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=316350 $D=103
M1167 4004 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=316840 $D=103
M1168 60 VSS 4006 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=319750 $D=103
M1169 4007 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=320240 $D=103
M1170 60 VSS 4009 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=323150 $D=103
M1171 4012 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=323640 $D=103
M1172 60 VSS 4014 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=326550 $D=103
M1173 4015 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=327040 $D=103
M1174 60 VSS 4017 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=329950 $D=103
M1175 4020 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=330440 $D=103
M1176 60 VSS 4022 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=333350 $D=103
M1177 4023 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=333840 $D=103
M1178 60 VSS 4025 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=336750 $D=103
M1179 4028 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=337240 $D=103
M1180 60 VSS 4030 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=340150 $D=103
M1181 4031 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=340640 $D=103
M1182 60 VSS 4033 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=343550 $D=103
M1183 4036 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=344040 $D=103
M1184 60 VSS 4038 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=346950 $D=103
M1185 4039 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=347440 $D=103
M1186 60 VSS 4041 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=350350 $D=103
M1187 4044 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=350840 $D=103
M1188 60 VSS 4046 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=353750 $D=103
M1189 4047 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=354240 $D=103
M1190 60 VSS 4049 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=357150 $D=103
M1191 4052 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=357640 $D=103
M1192 60 VSS 4054 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=360550 $D=103
M1193 4055 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=361040 $D=103
M1194 60 VSS 4057 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=363950 $D=103
M1195 4060 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=364440 $D=103
M1196 60 VSS 4062 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=367350 $D=103
M1197 4063 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=367840 $D=103
M1198 60 VSS 4065 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=370750 $D=103
M1199 4068 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=371240 $D=103
M1200 60 VSS 4070 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=374150 $D=103
M1201 4071 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=374640 $D=103
M1202 60 VSS 4073 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=377550 $D=103
M1203 4076 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=378040 $D=103
M1204 60 VSS 4078 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=380950 $D=103
M1205 4079 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=381440 $D=103
M1206 60 VSS 4081 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=384350 $D=103
M1207 4084 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=384840 $D=103
M1208 60 VSS 4086 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=387750 $D=103
M1209 4087 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=388240 $D=103
M1210 60 VSS 4089 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=391150 $D=103
M1211 4092 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=391640 $D=103
M1212 60 VSS 4094 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=394550 $D=103
M1213 4095 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=395040 $D=103
M1214 60 VSS 4097 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=397950 $D=103
M1215 4100 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=398440 $D=103
M1216 60 VSS 4102 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=401350 $D=103
M1217 4103 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=401840 $D=103
M1218 60 VSS 4105 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=404750 $D=103
M1219 4108 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=405240 $D=103
M1220 60 VSS 4110 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=408150 $D=103
M1221 4111 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=408640 $D=103
M1222 60 VSS 4113 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=411550 $D=103
M1223 4116 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=412040 $D=103
M1224 60 VSS 4118 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=414950 $D=103
M1225 4119 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=415440 $D=103
M1226 60 VSS 4121 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=418350 $D=103
M1227 4124 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=418840 $D=103
M1228 60 VSS 4126 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=421750 $D=103
M1229 4127 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=422240 $D=103
M1230 60 VSS 4129 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=425150 $D=103
M1231 4132 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=425640 $D=103
M1232 60 VSS 4134 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=428550 $D=103
M1233 4135 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=429040 $D=103
M1234 60 VSS 4137 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=431950 $D=103
M1235 4140 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=432440 $D=103
M1236 60 VSS 4142 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=435350 $D=103
M1237 4143 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=435840 $D=103
M1238 60 VSS 4145 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=438750 $D=103
M1239 4148 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=439240 $D=103
M1240 60 VSS 4150 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=442150 $D=103
M1241 4151 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=442640 $D=103
M1242 60 VSS 4153 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=445550 $D=103
M1243 4156 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=446040 $D=103
M1244 60 VSS 4158 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=448950 $D=103
M1245 4159 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=449440 $D=103
M1246 60 VSS 4161 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=452350 $D=103
M1247 4164 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=452840 $D=103
M1248 60 VSS 4166 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=455750 $D=103
M1249 4167 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=456240 $D=103
M1250 60 VSS 4169 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=459150 $D=103
M1251 4172 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=459640 $D=103
M1252 60 VSS 4174 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=462550 $D=103
M1253 4175 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=463040 $D=103
M1254 60 VSS 4177 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=465950 $D=103
M1255 4180 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=466440 $D=103
M1256 60 VSS 4182 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=469350 $D=103
M1257 4183 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=469840 $D=103
M1258 60 VSS 4185 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=472750 $D=103
M1259 4188 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=473240 $D=103
M1260 60 VSS 4190 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=476150 $D=103
M1261 4191 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=476640 $D=103
M1262 60 VSS 4193 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=479550 $D=103
M1263 4196 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=480040 $D=103
M1264 60 VSS 4198 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=482950 $D=103
M1265 4199 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=483440 $D=103
M1266 60 VSS 4201 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=486350 $D=103
M1267 4204 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=486840 $D=103
M1268 60 VSS 4206 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=489750 $D=103
M1269 4207 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=490240 $D=103
M1270 60 VSS 4209 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=493150 $D=103
M1271 4212 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=493640 $D=103
M1272 60 VSS 4214 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=496550 $D=103
M1273 4215 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=497040 $D=103
M1274 60 VSS 4217 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=499950 $D=103
M1275 4220 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=500440 $D=103
M1276 60 VSS 4222 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=503350 $D=103
M1277 4223 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=503840 $D=103
M1278 60 VSS 4225 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=506750 $D=103
M1279 4228 VSS 60 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235080 $Y=507240 $D=103
M1280 61 VSS 3717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=74950 $D=103
M1281 3720 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=75440 $D=103
M1282 61 VSS 3722 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=78350 $D=103
M1283 3723 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=78840 $D=103
M1284 61 VSS 3725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=81750 $D=103
M1285 3728 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=82240 $D=103
M1286 61 VSS 3730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=85150 $D=103
M1287 3731 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=85640 $D=103
M1288 61 VSS 3733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=88550 $D=103
M1289 3736 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=89040 $D=103
M1290 61 VSS 3738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=91950 $D=103
M1291 3739 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=92440 $D=103
M1292 61 VSS 3741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=95350 $D=103
M1293 3744 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=95840 $D=103
M1294 61 VSS 3746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=98750 $D=103
M1295 3747 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=99240 $D=103
M1296 61 VSS 3749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=102150 $D=103
M1297 3752 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=102640 $D=103
M1298 61 VSS 3754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=105550 $D=103
M1299 3755 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=106040 $D=103
M1300 61 VSS 3757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=108950 $D=103
M1301 3760 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=109440 $D=103
M1302 61 VSS 3762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=112350 $D=103
M1303 3763 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=112840 $D=103
M1304 61 VSS 3765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=115750 $D=103
M1305 3768 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=116240 $D=103
M1306 61 VSS 3770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=119150 $D=103
M1307 3771 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=119640 $D=103
M1308 61 VSS 3773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=122550 $D=103
M1309 3776 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=123040 $D=103
M1310 61 VSS 3778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=125950 $D=103
M1311 3779 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=126440 $D=103
M1312 61 VSS 3781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=129350 $D=103
M1313 3784 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=129840 $D=103
M1314 61 VSS 3786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=132750 $D=103
M1315 3787 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=133240 $D=103
M1316 61 VSS 3789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=136150 $D=103
M1317 3792 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=136640 $D=103
M1318 61 VSS 3794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=139550 $D=103
M1319 3795 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=140040 $D=103
M1320 61 VSS 3797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=142950 $D=103
M1321 3800 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=143440 $D=103
M1322 61 VSS 3802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=146350 $D=103
M1323 3803 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=146840 $D=103
M1324 61 VSS 3805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=149750 $D=103
M1325 3808 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=150240 $D=103
M1326 61 VSS 3810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=153150 $D=103
M1327 3811 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=153640 $D=103
M1328 61 VSS 3813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=156550 $D=103
M1329 3816 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=157040 $D=103
M1330 61 VSS 3818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=159950 $D=103
M1331 3819 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=160440 $D=103
M1332 61 VSS 3821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=163350 $D=103
M1333 3824 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=163840 $D=103
M1334 61 VSS 3826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=166750 $D=103
M1335 3827 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=167240 $D=103
M1336 61 VSS 3829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=170150 $D=103
M1337 3832 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=170640 $D=103
M1338 61 VSS 3834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=173550 $D=103
M1339 3835 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=174040 $D=103
M1340 61 VSS 3837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=176950 $D=103
M1341 3840 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=177440 $D=103
M1342 61 VSS 3842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=180350 $D=103
M1343 3843 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=180840 $D=103
M1344 61 VSS 3845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=183750 $D=103
M1345 3848 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=184240 $D=103
M1346 61 VSS 3850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=187150 $D=103
M1347 3851 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=187640 $D=103
M1348 61 VSS 3853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=190550 $D=103
M1349 3856 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=191040 $D=103
M1350 61 VSS 3858 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=193950 $D=103
M1351 3859 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=194440 $D=103
M1352 61 VSS 3861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=197350 $D=103
M1353 3864 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=197840 $D=103
M1354 61 VSS 3866 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=200750 $D=103
M1355 3867 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=201240 $D=103
M1356 61 VSS 3869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=204150 $D=103
M1357 3872 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=204640 $D=103
M1358 61 VSS 3874 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=207550 $D=103
M1359 3875 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=208040 $D=103
M1360 61 VSS 3877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=210950 $D=103
M1361 3880 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=211440 $D=103
M1362 61 VSS 3882 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=214350 $D=103
M1363 3883 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=214840 $D=103
M1364 61 VSS 3885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=217750 $D=103
M1365 3888 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=218240 $D=103
M1366 61 VSS 3890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=221150 $D=103
M1367 3891 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=221640 $D=103
M1368 61 VSS 3893 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=224550 $D=103
M1369 3896 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=225040 $D=103
M1370 61 VSS 3898 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=227950 $D=103
M1371 3899 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=228440 $D=103
M1372 61 VSS 3901 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=231350 $D=103
M1373 3904 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=231840 $D=103
M1374 61 VSS 3906 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=234750 $D=103
M1375 3907 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=235240 $D=103
M1376 61 VSS 3909 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=238150 $D=103
M1377 3912 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=238640 $D=103
M1378 61 VSS 3914 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=241550 $D=103
M1379 3915 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=242040 $D=103
M1380 61 VSS 3917 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=244950 $D=103
M1381 3920 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=245440 $D=103
M1382 61 VSS 3922 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=248350 $D=103
M1383 3923 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=248840 $D=103
M1384 61 VSS 3925 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=251750 $D=103
M1385 3928 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=252240 $D=103
M1386 61 VSS 3930 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=255150 $D=103
M1387 3931 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=255640 $D=103
M1388 61 VSS 3933 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=258550 $D=103
M1389 3936 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=259040 $D=103
M1390 61 VSS 3938 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=261950 $D=103
M1391 3939 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=262440 $D=103
M1392 61 VSS 3941 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=265350 $D=103
M1393 3944 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=265840 $D=103
M1394 61 VSS 3946 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=268750 $D=103
M1395 3947 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=269240 $D=103
M1396 61 VSS 3949 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=272150 $D=103
M1397 3952 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=272640 $D=103
M1398 61 VSS 3954 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=275550 $D=103
M1399 3955 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=276040 $D=103
M1400 61 VSS 3957 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=278950 $D=103
M1401 3960 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=279440 $D=103
M1402 61 VSS 3962 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=282350 $D=103
M1403 3963 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=282840 $D=103
M1404 61 VSS 3965 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=285750 $D=103
M1405 3968 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=286240 $D=103
M1406 61 VSS 3970 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=289150 $D=103
M1407 3971 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=289640 $D=103
M1408 61 VSS 3973 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=292550 $D=103
M1409 3976 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=293040 $D=103
M1410 61 VSS 3978 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=295950 $D=103
M1411 3979 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=296440 $D=103
M1412 61 VSS 3981 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=299350 $D=103
M1413 3984 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=299840 $D=103
M1414 61 VSS 3986 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=302750 $D=103
M1415 3987 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=303240 $D=103
M1416 61 VSS 3989 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=306150 $D=103
M1417 3992 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=306640 $D=103
M1418 61 VSS 3994 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=309550 $D=103
M1419 3995 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=310040 $D=103
M1420 61 VSS 3997 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=312950 $D=103
M1421 4000 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=313440 $D=103
M1422 61 VSS 4002 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=316350 $D=103
M1423 4003 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=316840 $D=103
M1424 61 VSS 4005 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=319750 $D=103
M1425 4008 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=320240 $D=103
M1426 61 VSS 4010 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=323150 $D=103
M1427 4011 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=323640 $D=103
M1428 61 VSS 4013 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=326550 $D=103
M1429 4016 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=327040 $D=103
M1430 61 VSS 4018 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=329950 $D=103
M1431 4019 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=330440 $D=103
M1432 61 VSS 4021 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=333350 $D=103
M1433 4024 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=333840 $D=103
M1434 61 VSS 4026 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=336750 $D=103
M1435 4027 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=337240 $D=103
M1436 61 VSS 4029 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=340150 $D=103
M1437 4032 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=340640 $D=103
M1438 61 VSS 4034 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=343550 $D=103
M1439 4035 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=344040 $D=103
M1440 61 VSS 4037 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=346950 $D=103
M1441 4040 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=347440 $D=103
M1442 61 VSS 4042 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=350350 $D=103
M1443 4043 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=350840 $D=103
M1444 61 VSS 4045 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=353750 $D=103
M1445 4048 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=354240 $D=103
M1446 61 VSS 4050 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=357150 $D=103
M1447 4051 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=357640 $D=103
M1448 61 VSS 4053 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=360550 $D=103
M1449 4056 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=361040 $D=103
M1450 61 VSS 4058 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=363950 $D=103
M1451 4059 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=364440 $D=103
M1452 61 VSS 4061 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=367350 $D=103
M1453 4064 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=367840 $D=103
M1454 61 VSS 4066 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=370750 $D=103
M1455 4067 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=371240 $D=103
M1456 61 VSS 4069 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=374150 $D=103
M1457 4072 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=374640 $D=103
M1458 61 VSS 4074 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=377550 $D=103
M1459 4075 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=378040 $D=103
M1460 61 VSS 4077 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=380950 $D=103
M1461 4080 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=381440 $D=103
M1462 61 VSS 4082 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=384350 $D=103
M1463 4083 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=384840 $D=103
M1464 61 VSS 4085 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=387750 $D=103
M1465 4088 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=388240 $D=103
M1466 61 VSS 4090 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=391150 $D=103
M1467 4091 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=391640 $D=103
M1468 61 VSS 4093 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=394550 $D=103
M1469 4096 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=395040 $D=103
M1470 61 VSS 4098 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=397950 $D=103
M1471 4099 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=398440 $D=103
M1472 61 VSS 4101 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=401350 $D=103
M1473 4104 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=401840 $D=103
M1474 61 VSS 4106 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=404750 $D=103
M1475 4107 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=405240 $D=103
M1476 61 VSS 4109 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=408150 $D=103
M1477 4112 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=408640 $D=103
M1478 61 VSS 4114 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=411550 $D=103
M1479 4115 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=412040 $D=103
M1480 61 VSS 4117 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=414950 $D=103
M1481 4120 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=415440 $D=103
M1482 61 VSS 4122 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=418350 $D=103
M1483 4123 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=418840 $D=103
M1484 61 VSS 4125 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=421750 $D=103
M1485 4128 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=422240 $D=103
M1486 61 VSS 4130 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=425150 $D=103
M1487 4131 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=425640 $D=103
M1488 61 VSS 4133 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=428550 $D=103
M1489 4136 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=429040 $D=103
M1490 61 VSS 4138 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=431950 $D=103
M1491 4139 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=432440 $D=103
M1492 61 VSS 4141 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=435350 $D=103
M1493 4144 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=435840 $D=103
M1494 61 VSS 4146 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=438750 $D=103
M1495 4147 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=439240 $D=103
M1496 61 VSS 4149 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=442150 $D=103
M1497 4152 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=442640 $D=103
M1498 61 VSS 4154 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=445550 $D=103
M1499 4155 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=446040 $D=103
M1500 61 VSS 4157 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=448950 $D=103
M1501 4160 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=449440 $D=103
M1502 61 VSS 4162 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=452350 $D=103
M1503 4163 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=452840 $D=103
M1504 61 VSS 4165 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=455750 $D=103
M1505 4168 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=456240 $D=103
M1506 61 VSS 4170 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=459150 $D=103
M1507 4171 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=459640 $D=103
M1508 61 VSS 4173 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=462550 $D=103
M1509 4176 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=463040 $D=103
M1510 61 VSS 4178 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=465950 $D=103
M1511 4179 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=466440 $D=103
M1512 61 VSS 4181 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=469350 $D=103
M1513 4184 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=469840 $D=103
M1514 61 VSS 4186 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=472750 $D=103
M1515 4187 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=473240 $D=103
M1516 61 VSS 4189 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=476150 $D=103
M1517 4192 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=476640 $D=103
M1518 61 VSS 4194 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=479550 $D=103
M1519 4195 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=480040 $D=103
M1520 61 VSS 4197 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=482950 $D=103
M1521 4200 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=483440 $D=103
M1522 61 VSS 4202 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=486350 $D=103
M1523 4203 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=486840 $D=103
M1524 61 VSS 4205 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=489750 $D=103
M1525 4208 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=490240 $D=103
M1526 61 VSS 4210 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=493150 $D=103
M1527 4211 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=493640 $D=103
M1528 61 VSS 4213 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=496550 $D=103
M1529 4216 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=497040 $D=103
M1530 61 VSS 4218 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=499950 $D=103
M1531 4219 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=500440 $D=103
M1532 61 VSS 4221 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=503350 $D=103
M1533 4224 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=503840 $D=103
M1534 61 VSS 4226 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=506750 $D=103
M1535 4227 VSS 61 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=235940 $Y=507240 $D=103
M1536 5376 63 5377 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=74950 $D=103
M1537 5378 64 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=75440 $D=103
M1538 5376 65 5379 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=78350 $D=103
M1539 5380 66 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=78840 $D=103
M1540 5376 67 5381 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=81750 $D=103
M1541 5382 68 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=82240 $D=103
M1542 5376 69 5383 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=85150 $D=103
M1543 5384 70 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=85640 $D=103
M1544 5376 71 5385 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=88550 $D=103
M1545 5386 72 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=89040 $D=103
M1546 5376 73 5387 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=91950 $D=103
M1547 5388 74 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=92440 $D=103
M1548 5376 75 5389 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=95350 $D=103
M1549 5390 76 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=95840 $D=103
M1550 5376 77 5391 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=98750 $D=103
M1551 5392 78 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=99240 $D=103
M1552 5376 79 5393 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=102150 $D=103
M1553 5394 80 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=102640 $D=103
M1554 5376 81 5395 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=105550 $D=103
M1555 5396 82 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=106040 $D=103
M1556 5376 83 5397 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=108950 $D=103
M1557 5398 84 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=109440 $D=103
M1558 5376 85 5399 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=112350 $D=103
M1559 5400 86 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=112840 $D=103
M1560 5376 87 5401 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=115750 $D=103
M1561 5402 88 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=116240 $D=103
M1562 5376 89 5403 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=119150 $D=103
M1563 5404 90 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=119640 $D=103
M1564 5376 91 5405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=122550 $D=103
M1565 5406 92 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=123040 $D=103
M1566 5376 93 5407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=125950 $D=103
M1567 5408 94 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=126440 $D=103
M1568 5376 95 5409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=129350 $D=103
M1569 5410 96 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=129840 $D=103
M1570 5376 97 5411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=132750 $D=103
M1571 5412 98 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=133240 $D=103
M1572 5376 99 5413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=136150 $D=103
M1573 5414 100 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=136640 $D=103
M1574 5376 101 5415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=139550 $D=103
M1575 5416 102 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=140040 $D=103
M1576 5376 103 5417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=142950 $D=103
M1577 5418 104 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=143440 $D=103
M1578 5376 105 5419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=146350 $D=103
M1579 5420 106 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=146840 $D=103
M1580 5376 107 5421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=149750 $D=103
M1581 5422 108 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=150240 $D=103
M1582 5376 109 5423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=153150 $D=103
M1583 5424 110 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=153640 $D=103
M1584 5376 111 5425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=156550 $D=103
M1585 5426 112 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=157040 $D=103
M1586 5376 113 5427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=159950 $D=103
M1587 5428 114 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=160440 $D=103
M1588 5376 115 5429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=163350 $D=103
M1589 5430 116 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=163840 $D=103
M1590 5376 117 5431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=166750 $D=103
M1591 5432 118 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=167240 $D=103
M1592 5376 119 5433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=170150 $D=103
M1593 5434 120 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=170640 $D=103
M1594 5376 121 5435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=173550 $D=103
M1595 5436 122 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=174040 $D=103
M1596 5376 123 5437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=176950 $D=103
M1597 5438 124 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=177440 $D=103
M1598 5376 125 5439 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=180350 $D=103
M1599 5440 126 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=180840 $D=103
M1600 5376 127 5441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=183750 $D=103
M1601 5442 128 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=184240 $D=103
M1602 5376 129 5443 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=187150 $D=103
M1603 5444 130 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=187640 $D=103
M1604 5376 131 5445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=190550 $D=103
M1605 5446 132 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=191040 $D=103
M1606 5376 133 5447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=193950 $D=103
M1607 5448 134 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=194440 $D=103
M1608 5376 135 5449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=197350 $D=103
M1609 5450 136 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=197840 $D=103
M1610 5376 137 5451 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=200750 $D=103
M1611 5452 138 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=201240 $D=103
M1612 5376 139 5453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=204150 $D=103
M1613 5454 140 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=204640 $D=103
M1614 5376 141 5455 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=207550 $D=103
M1615 5456 142 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=208040 $D=103
M1616 5376 143 5457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=210950 $D=103
M1617 5458 144 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=211440 $D=103
M1618 5376 145 5459 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=214350 $D=103
M1619 5460 146 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=214840 $D=103
M1620 5376 147 5461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=217750 $D=103
M1621 5462 148 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=218240 $D=103
M1622 5376 149 5463 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=221150 $D=103
M1623 5464 150 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=221640 $D=103
M1624 5376 151 5465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=224550 $D=103
M1625 5466 152 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=225040 $D=103
M1626 5376 153 5467 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=227950 $D=103
M1627 5468 154 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=228440 $D=103
M1628 5376 155 5469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=231350 $D=103
M1629 5470 156 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=231840 $D=103
M1630 5376 157 5471 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=234750 $D=103
M1631 5472 158 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=235240 $D=103
M1632 5376 159 5473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=238150 $D=103
M1633 5474 160 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=238640 $D=103
M1634 5376 161 5475 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=241550 $D=103
M1635 5476 162 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=242040 $D=103
M1636 5376 163 5477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=244950 $D=103
M1637 5478 164 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=245440 $D=103
M1638 5376 165 5479 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=248350 $D=103
M1639 5480 166 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=248840 $D=103
M1640 5376 167 5481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=251750 $D=103
M1641 5482 168 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=252240 $D=103
M1642 5376 169 5483 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=255150 $D=103
M1643 5484 170 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=255640 $D=103
M1644 5376 171 5485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=258550 $D=103
M1645 5486 172 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=259040 $D=103
M1646 5376 173 5487 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=261950 $D=103
M1647 5488 174 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=262440 $D=103
M1648 5376 175 5489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=265350 $D=103
M1649 5490 176 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=265840 $D=103
M1650 5376 177 5491 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=268750 $D=103
M1651 5492 178 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=269240 $D=103
M1652 5376 179 5493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=272150 $D=103
M1653 5494 180 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=272640 $D=103
M1654 5376 181 5495 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=275550 $D=103
M1655 5496 182 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=276040 $D=103
M1656 5376 183 5497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=278950 $D=103
M1657 5498 184 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=279440 $D=103
M1658 5376 185 5499 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=282350 $D=103
M1659 5500 186 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=282840 $D=103
M1660 5376 187 5501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=285750 $D=103
M1661 5502 188 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=286240 $D=103
M1662 5376 189 5503 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=289150 $D=103
M1663 5504 190 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=289640 $D=103
M1664 5376 191 5505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=292550 $D=103
M1665 5506 192 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=293040 $D=103
M1666 5376 193 5507 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=295950 $D=103
M1667 5508 194 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=296440 $D=103
M1668 5376 195 5509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=299350 $D=103
M1669 5510 196 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=299840 $D=103
M1670 5376 197 5511 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=302750 $D=103
M1671 5512 198 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=303240 $D=103
M1672 5376 199 5513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=306150 $D=103
M1673 5514 200 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=306640 $D=103
M1674 5376 201 5515 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=309550 $D=103
M1675 5516 202 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=310040 $D=103
M1676 5376 203 5517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=312950 $D=103
M1677 5518 204 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=313440 $D=103
M1678 5376 205 5519 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=316350 $D=103
M1679 5520 206 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=316840 $D=103
M1680 5376 207 5521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=319750 $D=103
M1681 5522 208 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=320240 $D=103
M1682 5376 209 5523 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=323150 $D=103
M1683 5524 210 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=323640 $D=103
M1684 5376 211 5525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=326550 $D=103
M1685 5526 212 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=327040 $D=103
M1686 5376 213 5527 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=329950 $D=103
M1687 5528 214 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=330440 $D=103
M1688 5376 215 5529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=333350 $D=103
M1689 5530 216 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=333840 $D=103
M1690 5376 217 5531 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=336750 $D=103
M1691 5532 218 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=337240 $D=103
M1692 5376 219 5533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=340150 $D=103
M1693 5534 220 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=340640 $D=103
M1694 5376 221 5535 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=343550 $D=103
M1695 5536 222 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=344040 $D=103
M1696 5376 223 5537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=346950 $D=103
M1697 5538 224 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=347440 $D=103
M1698 5376 225 5539 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=350350 $D=103
M1699 5540 226 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=350840 $D=103
M1700 5376 227 5541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=353750 $D=103
M1701 5542 228 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=354240 $D=103
M1702 5376 229 5543 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=357150 $D=103
M1703 5544 230 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=357640 $D=103
M1704 5376 231 5545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=360550 $D=103
M1705 5546 232 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=361040 $D=103
M1706 5376 233 5547 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=363950 $D=103
M1707 5548 234 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=364440 $D=103
M1708 5376 235 5549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=367350 $D=103
M1709 5550 236 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=367840 $D=103
M1710 5376 237 5551 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=370750 $D=103
M1711 5552 238 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=371240 $D=103
M1712 5376 239 5553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=374150 $D=103
M1713 5554 240 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=374640 $D=103
M1714 5376 241 5555 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=377550 $D=103
M1715 5556 242 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=378040 $D=103
M1716 5376 243 5557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=380950 $D=103
M1717 5558 244 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=381440 $D=103
M1718 5376 245 5559 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=384350 $D=103
M1719 5560 246 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=384840 $D=103
M1720 5376 247 5561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=387750 $D=103
M1721 5562 248 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=388240 $D=103
M1722 5376 249 5563 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=391150 $D=103
M1723 5564 250 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=391640 $D=103
M1724 5376 251 5565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=394550 $D=103
M1725 5566 252 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=395040 $D=103
M1726 5376 253 5567 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=397950 $D=103
M1727 5568 254 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=398440 $D=103
M1728 5376 255 5569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=401350 $D=103
M1729 5570 256 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=401840 $D=103
M1730 5376 257 5571 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=404750 $D=103
M1731 5572 258 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=405240 $D=103
M1732 5376 259 5573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=408150 $D=103
M1733 5574 260 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=408640 $D=103
M1734 5376 261 5575 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=411550 $D=103
M1735 5576 262 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=412040 $D=103
M1736 5376 263 5577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=414950 $D=103
M1737 5578 264 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=415440 $D=103
M1738 5376 265 5579 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=418350 $D=103
M1739 5580 266 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=418840 $D=103
M1740 5376 267 5581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=421750 $D=103
M1741 5582 268 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=422240 $D=103
M1742 5376 269 5583 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=425150 $D=103
M1743 5584 270 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=425640 $D=103
M1744 5376 271 5585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=428550 $D=103
M1745 5586 272 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=429040 $D=103
M1746 5376 273 5587 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=431950 $D=103
M1747 5588 274 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=432440 $D=103
M1748 5376 275 5589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=435350 $D=103
M1749 5590 276 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=435840 $D=103
M1750 5376 277 5591 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=438750 $D=103
M1751 5592 278 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=439240 $D=103
M1752 5376 279 5593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=442150 $D=103
M1753 5594 280 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=442640 $D=103
M1754 5376 281 5595 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=445550 $D=103
M1755 5596 282 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=446040 $D=103
M1756 5376 283 5597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=448950 $D=103
M1757 5598 284 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=449440 $D=103
M1758 5376 285 5599 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=452350 $D=103
M1759 5600 286 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=452840 $D=103
M1760 5376 287 5601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=455750 $D=103
M1761 5602 288 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=456240 $D=103
M1762 5376 289 5603 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=459150 $D=103
M1763 5604 290 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=459640 $D=103
M1764 5376 291 5605 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=462550 $D=103
M1765 5606 292 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=463040 $D=103
M1766 5376 293 5607 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=465950 $D=103
M1767 5608 294 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=466440 $D=103
M1768 5376 295 5609 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=469350 $D=103
M1769 5610 296 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=469840 $D=103
M1770 5376 297 5611 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=472750 $D=103
M1771 5612 298 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=473240 $D=103
M1772 5376 299 5613 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=476150 $D=103
M1773 5614 300 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=476640 $D=103
M1774 5376 301 5615 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=479550 $D=103
M1775 5616 302 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=480040 $D=103
M1776 5376 303 5617 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=482950 $D=103
M1777 5618 304 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=483440 $D=103
M1778 5376 305 5619 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=486350 $D=103
M1779 5620 306 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=486840 $D=103
M1780 5376 307 5621 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=489750 $D=103
M1781 5622 308 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=490240 $D=103
M1782 5376 309 5623 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=493150 $D=103
M1783 5624 310 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=493640 $D=103
M1784 5376 311 5625 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=496550 $D=103
M1785 5626 312 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=497040 $D=103
M1786 5376 313 5627 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=499950 $D=103
M1787 5628 314 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=500440 $D=103
M1788 5376 315 5629 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=503350 $D=103
M1789 5630 316 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=503840 $D=103
M1790 5376 317 5631 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=506750 $D=103
M1791 5632 318 5376 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=507240 $D=103
M1792 405 50 3461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=511190 $D=103
M1793 3464 50 405 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=237480 $Y=511680 $D=103
M1794 406 50 3462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=238340 $Y=511190 $D=103
M1795 3463 50 406 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=238340 $Y=511680 $D=103
M1796 531 50 4230 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=238680 $Y=511190 $D=103
M1797 4231 50 531 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=238680 $Y=511680 $D=103
M1798 532 50 4229 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=239540 $Y=511190 $D=103
M1799 4232 50 532 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=239540 $Y=511680 $D=103
M1800 655 50 4477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=239880 $Y=511190 $D=103
M1801 4480 50 655 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=239880 $Y=511680 $D=103
M1802 656 50 4478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=240740 $Y=511190 $D=103
M1803 4479 50 656 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=240740 $Y=511680 $D=103
M1804 781 50 4730 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=241080 $Y=511190 $D=103
M1805 4731 50 781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=241080 $Y=511680 $D=103
M1806 782 50 4729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=241940 $Y=511190 $D=103
M1807 4732 50 782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=241940 $Y=511680 $D=103
M1808 407 50 3465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=242280 $Y=511190 $D=103
M1809 3468 50 407 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=242280 $Y=511680 $D=103
M1810 408 50 3466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=243140 $Y=511190 $D=103
M1811 3467 50 408 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=243140 $Y=511680 $D=103
M1812 533 50 4234 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=243480 $Y=511190 $D=103
M1813 4235 50 533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=243480 $Y=511680 $D=103
M1814 534 50 4233 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=244340 $Y=511190 $D=103
M1815 4236 50 534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=244340 $Y=511680 $D=103
M1816 657 50 4481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=244680 $Y=511190 $D=103
M1817 4484 50 657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=244680 $Y=511680 $D=103
M1818 658 50 4482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=245540 $Y=511190 $D=103
M1819 4483 50 658 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=245540 $Y=511680 $D=103
M1820 783 50 4734 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=245880 $Y=511190 $D=103
M1821 4735 50 783 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=245880 $Y=511680 $D=103
M1822 784 50 4733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=246740 $Y=511190 $D=103
M1823 4736 50 784 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=246740 $Y=511680 $D=103
M1824 409 50 3469 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=247080 $Y=511190 $D=103
M1825 3472 50 409 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=247080 $Y=511680 $D=103
M1826 410 50 3470 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=247940 $Y=511190 $D=103
M1827 3471 50 410 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=247940 $Y=511680 $D=103
M1828 535 50 4238 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=248280 $Y=511190 $D=103
M1829 4239 50 535 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=248280 $Y=511680 $D=103
M1830 536 50 4237 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=249140 $Y=511190 $D=103
M1831 4240 50 536 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=249140 $Y=511680 $D=103
M1832 659 50 4485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=249480 $Y=511190 $D=103
M1833 4488 50 659 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=249480 $Y=511680 $D=103
M1834 660 50 4486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=250340 $Y=511190 $D=103
M1835 4487 50 660 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=250340 $Y=511680 $D=103
M1836 785 50 4738 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=250680 $Y=511190 $D=103
M1837 4739 50 785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=250680 $Y=511680 $D=103
M1838 786 50 4737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=251540 $Y=511190 $D=103
M1839 4740 50 786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=251540 $Y=511680 $D=103
M1840 411 50 3473 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=251880 $Y=511190 $D=103
M1841 3476 50 411 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=251880 $Y=511680 $D=103
M1842 412 50 3474 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=252740 $Y=511190 $D=103
M1843 3475 50 412 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=252740 $Y=511680 $D=103
M1844 537 50 4242 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=253080 $Y=511190 $D=103
M1845 4243 50 537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=253080 $Y=511680 $D=103
M1846 538 50 4241 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=253940 $Y=511190 $D=103
M1847 4244 50 538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=253940 $Y=511680 $D=103
M1848 661 50 4489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=254280 $Y=511190 $D=103
M1849 4492 50 661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=254280 $Y=511680 $D=103
M1850 662 50 4490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=255140 $Y=511190 $D=103
M1851 4491 50 662 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=255140 $Y=511680 $D=103
M1852 787 50 4742 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=255480 $Y=511190 $D=103
M1853 4743 50 787 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=255480 $Y=511680 $D=103
M1854 788 50 4741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=256340 $Y=511190 $D=103
M1855 4744 50 788 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=256340 $Y=511680 $D=103
M1856 413 50 3477 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=256680 $Y=511190 $D=103
M1857 3480 50 413 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=256680 $Y=511680 $D=103
M1858 414 50 3478 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=257540 $Y=511190 $D=103
M1859 3479 50 414 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=257540 $Y=511680 $D=103
M1860 539 50 4246 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=257880 $Y=511190 $D=103
M1861 4247 50 539 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=257880 $Y=511680 $D=103
M1862 540 50 4245 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=258740 $Y=511190 $D=103
M1863 4248 50 540 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=258740 $Y=511680 $D=103
M1864 663 50 4493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=259080 $Y=511190 $D=103
M1865 4496 50 663 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=259080 $Y=511680 $D=103
M1866 664 50 4494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=259940 $Y=511190 $D=103
M1867 4495 50 664 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=259940 $Y=511680 $D=103
M1868 789 50 4746 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=260280 $Y=511190 $D=103
M1869 4747 50 789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=260280 $Y=511680 $D=103
M1870 790 50 4745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=261140 $Y=511190 $D=103
M1871 4748 50 790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=261140 $Y=511680 $D=103
M1872 415 50 3481 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=261480 $Y=511190 $D=103
M1873 3484 50 415 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=261480 $Y=511680 $D=103
M1874 416 50 3482 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=262340 $Y=511190 $D=103
M1875 3483 50 416 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=262340 $Y=511680 $D=103
M1876 541 50 4250 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=262680 $Y=511190 $D=103
M1877 4251 50 541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=262680 $Y=511680 $D=103
M1878 542 50 4249 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=263540 $Y=511190 $D=103
M1879 4252 50 542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=263540 $Y=511680 $D=103
M1880 665 50 4497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=263880 $Y=511190 $D=103
M1881 4500 50 665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=263880 $Y=511680 $D=103
M1882 666 50 4498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=264740 $Y=511190 $D=103
M1883 4499 50 666 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=264740 $Y=511680 $D=103
M1884 791 50 4750 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=265080 $Y=511190 $D=103
M1885 4751 50 791 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=265080 $Y=511680 $D=103
M1886 792 50 4749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=265940 $Y=511190 $D=103
M1887 4752 50 792 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=265940 $Y=511680 $D=103
M1888 417 50 3485 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=266280 $Y=511190 $D=103
M1889 3488 50 417 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=266280 $Y=511680 $D=103
M1890 418 50 3486 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=267140 $Y=511190 $D=103
M1891 3487 50 418 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=267140 $Y=511680 $D=103
M1892 543 50 4254 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=267480 $Y=511190 $D=103
M1893 4255 50 543 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=267480 $Y=511680 $D=103
M1894 544 50 4253 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=268340 $Y=511190 $D=103
M1895 4256 50 544 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=268340 $Y=511680 $D=103
M1896 667 50 4501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=268680 $Y=511190 $D=103
M1897 4504 50 667 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=268680 $Y=511680 $D=103
M1898 668 50 4502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=269540 $Y=511190 $D=103
M1899 4503 50 668 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=269540 $Y=511680 $D=103
M1900 793 50 4754 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=269880 $Y=511190 $D=103
M1901 4755 50 793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=269880 $Y=511680 $D=103
M1902 794 50 4753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=270740 $Y=511190 $D=103
M1903 4756 50 794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=270740 $Y=511680 $D=103
M1904 419 50 3489 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=271080 $Y=511190 $D=103
M1905 3492 50 419 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=271080 $Y=511680 $D=103
M1906 420 50 3490 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=271940 $Y=511190 $D=103
M1907 3491 50 420 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=271940 $Y=511680 $D=103
M1908 545 50 4258 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=272280 $Y=511190 $D=103
M1909 4259 50 545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=272280 $Y=511680 $D=103
M1910 546 50 4257 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=273140 $Y=511190 $D=103
M1911 4260 50 546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=273140 $Y=511680 $D=103
M1912 669 50 4505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=273480 $Y=511190 $D=103
M1913 4508 50 669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=273480 $Y=511680 $D=103
M1914 670 50 4506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=274340 $Y=511190 $D=103
M1915 4507 50 670 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=274340 $Y=511680 $D=103
M1916 795 50 4758 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=274680 $Y=511190 $D=103
M1917 4759 50 795 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=274680 $Y=511680 $D=103
M1918 796 50 4757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=275540 $Y=511190 $D=103
M1919 4760 50 796 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=275540 $Y=511680 $D=103
M1920 421 50 3493 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=277080 $Y=511190 $D=103
M1921 3496 50 421 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=277080 $Y=511680 $D=103
M1922 422 50 3494 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=277940 $Y=511190 $D=103
M1923 3495 50 422 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=277940 $Y=511680 $D=103
M1924 547 50 4262 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=278280 $Y=511190 $D=103
M1925 4263 50 547 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=278280 $Y=511680 $D=103
M1926 548 50 4261 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=279140 $Y=511190 $D=103
M1927 4264 50 548 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=279140 $Y=511680 $D=103
M1928 671 50 4509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=279480 $Y=511190 $D=103
M1929 4512 50 671 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=279480 $Y=511680 $D=103
M1930 672 50 4510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=280340 $Y=511190 $D=103
M1931 4511 50 672 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=280340 $Y=511680 $D=103
M1932 797 50 4762 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=280680 $Y=511190 $D=103
M1933 4763 50 797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=280680 $Y=511680 $D=103
M1934 798 50 4761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=281540 $Y=511190 $D=103
M1935 4764 50 798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=281540 $Y=511680 $D=103
M1936 423 50 3497 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=281880 $Y=511190 $D=103
M1937 3500 50 423 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=281880 $Y=511680 $D=103
M1938 424 50 3498 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=282740 $Y=511190 $D=103
M1939 3499 50 424 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=282740 $Y=511680 $D=103
M1940 549 50 4266 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=283080 $Y=511190 $D=103
M1941 4267 50 549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=283080 $Y=511680 $D=103
M1942 550 50 4265 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=283940 $Y=511190 $D=103
M1943 4268 50 550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=283940 $Y=511680 $D=103
M1944 673 50 4513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=284280 $Y=511190 $D=103
M1945 4516 50 673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=284280 $Y=511680 $D=103
M1946 674 50 4514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=285140 $Y=511190 $D=103
M1947 4515 50 674 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=285140 $Y=511680 $D=103
M1948 799 50 4766 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=285480 $Y=511190 $D=103
M1949 4767 50 799 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=285480 $Y=511680 $D=103
M1950 800 50 4765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=286340 $Y=511190 $D=103
M1951 4768 50 800 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=286340 $Y=511680 $D=103
M1952 425 50 3501 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=286680 $Y=511190 $D=103
M1953 3504 50 425 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=286680 $Y=511680 $D=103
M1954 426 50 3502 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=287540 $Y=511190 $D=103
M1955 3503 50 426 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=287540 $Y=511680 $D=103
M1956 551 50 4270 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=287880 $Y=511190 $D=103
M1957 4271 50 551 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=287880 $Y=511680 $D=103
M1958 552 50 4269 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=288740 $Y=511190 $D=103
M1959 4272 50 552 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=288740 $Y=511680 $D=103
M1960 675 50 4517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=289080 $Y=511190 $D=103
M1961 4520 50 675 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=289080 $Y=511680 $D=103
M1962 676 50 4518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=289940 $Y=511190 $D=103
M1963 4519 50 676 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=289940 $Y=511680 $D=103
M1964 801 50 4770 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=290280 $Y=511190 $D=103
M1965 4771 50 801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=290280 $Y=511680 $D=103
M1966 802 50 4769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=291140 $Y=511190 $D=103
M1967 4772 50 802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=291140 $Y=511680 $D=103
M1968 427 50 3505 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=291480 $Y=511190 $D=103
M1969 3508 50 427 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=291480 $Y=511680 $D=103
M1970 428 50 3506 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=292340 $Y=511190 $D=103
M1971 3507 50 428 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=292340 $Y=511680 $D=103
M1972 553 50 4274 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=292680 $Y=511190 $D=103
M1973 4275 50 553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=292680 $Y=511680 $D=103
M1974 554 50 4273 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=293540 $Y=511190 $D=103
M1975 4276 50 554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=293540 $Y=511680 $D=103
M1976 677 50 4521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=293880 $Y=511190 $D=103
M1977 4524 50 677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=293880 $Y=511680 $D=103
M1978 678 50 4522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=294740 $Y=511190 $D=103
M1979 4523 50 678 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=294740 $Y=511680 $D=103
M1980 803 50 4774 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=295080 $Y=511190 $D=103
M1981 4775 50 803 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=295080 $Y=511680 $D=103
M1982 804 50 4773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=295940 $Y=511190 $D=103
M1983 4776 50 804 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=295940 $Y=511680 $D=103
M1984 429 50 3509 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=296280 $Y=511190 $D=103
M1985 3512 50 429 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=296280 $Y=511680 $D=103
M1986 430 50 3510 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=297140 $Y=511190 $D=103
M1987 3511 50 430 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=297140 $Y=511680 $D=103
M1988 555 50 4278 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=297480 $Y=511190 $D=103
M1989 4279 50 555 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=297480 $Y=511680 $D=103
M1990 556 50 4277 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=298340 $Y=511190 $D=103
M1991 4280 50 556 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=298340 $Y=511680 $D=103
M1992 679 50 4525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=298680 $Y=511190 $D=103
M1993 4528 50 679 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=298680 $Y=511680 $D=103
M1994 680 50 4526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=299540 $Y=511190 $D=103
M1995 4527 50 680 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=299540 $Y=511680 $D=103
M1996 805 50 4778 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=299880 $Y=511190 $D=103
M1997 4779 50 805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=299880 $Y=511680 $D=103
M1998 806 50 4777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=300740 $Y=511190 $D=103
M1999 4780 50 806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=300740 $Y=511680 $D=103
M2000 431 50 3513 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=301080 $Y=511190 $D=103
M2001 3516 50 431 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=301080 $Y=511680 $D=103
M2002 432 50 3514 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=301940 $Y=511190 $D=103
M2003 3515 50 432 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=301940 $Y=511680 $D=103
M2004 557 50 4282 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=302280 $Y=511190 $D=103
M2005 4283 50 557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=302280 $Y=511680 $D=103
M2006 558 50 4281 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=303140 $Y=511190 $D=103
M2007 4284 50 558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=303140 $Y=511680 $D=103
M2008 681 50 4529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=303480 $Y=511190 $D=103
M2009 4532 50 681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=303480 $Y=511680 $D=103
M2010 682 50 4530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=304340 $Y=511190 $D=103
M2011 4531 50 682 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=304340 $Y=511680 $D=103
M2012 807 50 4782 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=304680 $Y=511190 $D=103
M2013 4783 50 807 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=304680 $Y=511680 $D=103
M2014 808 50 4781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=305540 $Y=511190 $D=103
M2015 4784 50 808 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=305540 $Y=511680 $D=103
M2016 433 50 3517 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=305880 $Y=511190 $D=103
M2017 3520 50 433 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=305880 $Y=511680 $D=103
M2018 434 50 3518 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=306740 $Y=511190 $D=103
M2019 3519 50 434 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=306740 $Y=511680 $D=103
M2020 559 50 4286 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=307080 $Y=511190 $D=103
M2021 4287 50 559 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=307080 $Y=511680 $D=103
M2022 560 50 4285 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=307940 $Y=511190 $D=103
M2023 4288 50 560 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=307940 $Y=511680 $D=103
M2024 683 50 4533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=308280 $Y=511190 $D=103
M2025 4536 50 683 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=308280 $Y=511680 $D=103
M2026 684 50 4534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=309140 $Y=511190 $D=103
M2027 4535 50 684 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=309140 $Y=511680 $D=103
M2028 809 50 4786 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=309480 $Y=511190 $D=103
M2029 4787 50 809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=309480 $Y=511680 $D=103
M2030 810 50 4785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=310340 $Y=511190 $D=103
M2031 4788 50 810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=310340 $Y=511680 $D=103
M2032 435 50 3521 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=310680 $Y=511190 $D=103
M2033 3524 50 435 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=310680 $Y=511680 $D=103
M2034 436 50 3522 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=311540 $Y=511190 $D=103
M2035 3523 50 436 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=311540 $Y=511680 $D=103
M2036 561 50 4290 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=311880 $Y=511190 $D=103
M2037 4291 50 561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=311880 $Y=511680 $D=103
M2038 562 50 4289 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=312740 $Y=511190 $D=103
M2039 4292 50 562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=312740 $Y=511680 $D=103
M2040 685 50 4537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=313080 $Y=511190 $D=103
M2041 4540 50 685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=313080 $Y=511680 $D=103
M2042 686 50 4538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=313940 $Y=511190 $D=103
M2043 4539 50 686 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=313940 $Y=511680 $D=103
M2044 811 50 4790 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=314280 $Y=511190 $D=103
M2045 4791 50 811 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=314280 $Y=511680 $D=103
M2046 812 50 4789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=315140 $Y=511190 $D=103
M2047 4792 50 812 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=315140 $Y=511680 $D=103
M2048 337 50 5889 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=316680 $Y=511190 $D=103
M2049 5892 50 337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=316680 $Y=511680 $D=103
M2050 338 VSS 5890 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=317540 $Y=511190 $D=103
M2051 5891 VSS 338 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=317540 $Y=511680 $D=103
M2052 339 VSS 3586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=317880 $Y=511190 $D=103
M2053 3587 VSS 339 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=317880 $Y=511680 $D=103
M2054 340 VSS 3585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=318740 $Y=511190 $D=103
M2055 3588 VSS 340 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=318740 $Y=511680 $D=103
M2056 687 VSS 4541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=319080 $Y=511190 $D=103
M2057 4544 VSS 687 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=319080 $Y=511680 $D=103
M2058 688 VSS 4542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=319940 $Y=511190 $D=103
M2059 4543 VSS 688 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=319940 $Y=511680 $D=103
M2060 813 VSS 4794 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=320280 $Y=511190 $D=103
M2061 4795 VSS 813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=320280 $Y=511680 $D=103
M2062 814 VSS 4793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=321140 $Y=511190 $D=103
M2063 4796 VSS 814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=321140 $Y=511680 $D=103
M2064 437 VSS 3525 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=321480 $Y=511190 $D=103
M2065 3528 VSS 437 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=321480 $Y=511680 $D=103
M2066 438 VSS 3526 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=322340 $Y=511190 $D=103
M2067 3527 VSS 438 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=322340 $Y=511680 $D=103
M2068 563 VSS 4294 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=322680 $Y=511190 $D=103
M2069 4295 VSS 563 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=322680 $Y=511680 $D=103
M2070 564 VSS 4293 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=323540 $Y=511190 $D=103
M2071 4296 VSS 564 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=323540 $Y=511680 $D=103
M2072 689 VSS 4545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=323880 $Y=511190 $D=103
M2073 4548 VSS 689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=323880 $Y=511680 $D=103
M2074 690 VSS 4546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=324740 $Y=511190 $D=103
M2075 4547 VSS 690 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=324740 $Y=511680 $D=103
M2076 815 VSS 4798 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=325080 $Y=511190 $D=103
M2077 4799 VSS 815 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=325080 $Y=511680 $D=103
M2078 816 VSS 4797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=325940 $Y=511190 $D=103
M2079 4800 VSS 816 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=325940 $Y=511680 $D=103
M2080 439 VSS 3529 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=326280 $Y=511190 $D=103
M2081 3532 VSS 439 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=326280 $Y=511680 $D=103
M2082 440 VSS 3530 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=327140 $Y=511190 $D=103
M2083 3531 VSS 440 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=327140 $Y=511680 $D=103
M2084 565 VSS 4298 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=327480 $Y=511190 $D=103
M2085 4299 VSS 565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=327480 $Y=511680 $D=103
M2086 566 VSS 4297 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=328340 $Y=511190 $D=103
M2087 4300 VSS 566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=328340 $Y=511680 $D=103
M2088 691 VSS 4549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=328680 $Y=511190 $D=103
M2089 4552 VSS 691 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=328680 $Y=511680 $D=103
M2090 692 VSS 4550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=329540 $Y=511190 $D=103
M2091 4551 VSS 692 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=329540 $Y=511680 $D=103
M2092 817 VSS 4802 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=329880 $Y=511190 $D=103
M2093 4803 VSS 817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=329880 $Y=511680 $D=103
M2094 818 VSS 4801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=330740 $Y=511190 $D=103
M2095 4804 VSS 818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=330740 $Y=511680 $D=103
M2096 441 VSS 3533 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=331080 $Y=511190 $D=103
M2097 3536 VSS 441 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=331080 $Y=511680 $D=103
M2098 442 VSS 3534 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=331940 $Y=511190 $D=103
M2099 3535 VSS 442 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=331940 $Y=511680 $D=103
M2100 567 VSS 4302 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=332280 $Y=511190 $D=103
M2101 4303 VSS 567 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=332280 $Y=511680 $D=103
M2102 568 VSS 4301 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=333140 $Y=511190 $D=103
M2103 4304 VSS 568 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=333140 $Y=511680 $D=103
M2104 693 VSS 4553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=333480 $Y=511190 $D=103
M2105 4556 VSS 693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=333480 $Y=511680 $D=103
M2106 694 VSS 4554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=334340 $Y=511190 $D=103
M2107 4555 VSS 694 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=334340 $Y=511680 $D=103
M2108 819 VSS 4806 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=334680 $Y=511190 $D=103
M2109 4807 VSS 819 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=334680 $Y=511680 $D=103
M2110 820 VSS 4805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=335540 $Y=511190 $D=103
M2111 4808 VSS 820 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=335540 $Y=511680 $D=103
M2112 443 VSS 3537 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=335880 $Y=511190 $D=103
M2113 3540 VSS 443 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=335880 $Y=511680 $D=103
M2114 444 VSS 3538 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=336740 $Y=511190 $D=103
M2115 3539 VSS 444 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=336740 $Y=511680 $D=103
M2116 569 VSS 4306 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=337080 $Y=511190 $D=103
M2117 4307 VSS 569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=337080 $Y=511680 $D=103
M2118 570 VSS 4305 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=337940 $Y=511190 $D=103
M2119 4308 VSS 570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=337940 $Y=511680 $D=103
M2120 695 VSS 4557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=338280 $Y=511190 $D=103
M2121 4560 VSS 695 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=338280 $Y=511680 $D=103
M2122 696 VSS 4558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=339140 $Y=511190 $D=103
M2123 4559 VSS 696 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=339140 $Y=511680 $D=103
M2124 821 VSS 4810 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=339480 $Y=511190 $D=103
M2125 4811 VSS 821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=339480 $Y=511680 $D=103
M2126 822 VSS 4809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=340340 $Y=511190 $D=103
M2127 4812 VSS 822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=340340 $Y=511680 $D=103
M2128 445 VSS 3541 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=340680 $Y=511190 $D=103
M2129 3544 VSS 445 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=340680 $Y=511680 $D=103
M2130 446 VSS 3542 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=341540 $Y=511190 $D=103
M2131 3543 VSS 446 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=341540 $Y=511680 $D=103
M2132 571 VSS 4310 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=341880 $Y=511190 $D=103
M2133 4311 VSS 571 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=341880 $Y=511680 $D=103
M2134 572 VSS 4309 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=342740 $Y=511190 $D=103
M2135 4312 VSS 572 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=342740 $Y=511680 $D=103
M2136 697 VSS 4561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=343080 $Y=511190 $D=103
M2137 4564 VSS 697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=343080 $Y=511680 $D=103
M2138 698 VSS 4562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=343940 $Y=511190 $D=103
M2139 4563 VSS 698 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=343940 $Y=511680 $D=103
M2140 823 VSS 4814 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=344280 $Y=511190 $D=103
M2141 4815 VSS 823 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=344280 $Y=511680 $D=103
M2142 824 VSS 4813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=345140 $Y=511190 $D=103
M2143 4816 VSS 824 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=345140 $Y=511680 $D=103
M2144 447 VSS 3545 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=345480 $Y=511190 $D=103
M2145 3548 VSS 447 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=345480 $Y=511680 $D=103
M2146 448 VSS 3546 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=346340 $Y=511190 $D=103
M2147 3547 VSS 448 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=346340 $Y=511680 $D=103
M2148 573 VSS 4314 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=346680 $Y=511190 $D=103
M2149 4315 VSS 573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=346680 $Y=511680 $D=103
M2150 574 VSS 4313 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=347540 $Y=511190 $D=103
M2151 4316 VSS 574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=347540 $Y=511680 $D=103
M2152 699 VSS 4565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=347880 $Y=511190 $D=103
M2153 4568 VSS 699 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=347880 $Y=511680 $D=103
M2154 700 VSS 4566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=348740 $Y=511190 $D=103
M2155 4567 VSS 700 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=348740 $Y=511680 $D=103
M2156 825 VSS 4818 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=349080 $Y=511190 $D=103
M2157 4819 VSS 825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=349080 $Y=511680 $D=103
M2158 826 VSS 4817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=349940 $Y=511190 $D=103
M2159 4820 VSS 826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=349940 $Y=511680 $D=103
M2160 449 VSS 3549 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=350280 $Y=511190 $D=103
M2161 3552 VSS 449 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=350280 $Y=511680 $D=103
M2162 450 VSS 3550 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=351140 $Y=511190 $D=103
M2163 3551 VSS 450 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=351140 $Y=511680 $D=103
M2164 575 VSS 4318 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=351480 $Y=511190 $D=103
M2165 4319 VSS 575 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=351480 $Y=511680 $D=103
M2166 576 VSS 4317 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=352340 $Y=511190 $D=103
M2167 4320 VSS 576 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=352340 $Y=511680 $D=103
M2168 701 VSS 4569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=352680 $Y=511190 $D=103
M2169 4572 VSS 701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=352680 $Y=511680 $D=103
M2170 702 VSS 4570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=353540 $Y=511190 $D=103
M2171 4571 VSS 702 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=353540 $Y=511680 $D=103
M2172 827 VSS 4822 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=353880 $Y=511190 $D=103
M2173 4823 VSS 827 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=353880 $Y=511680 $D=103
M2174 828 VSS 4821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=354740 $Y=511190 $D=103
M2175 4824 VSS 828 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=354740 $Y=511680 $D=103
M2176 451 VSS 3553 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=356280 $Y=511190 $D=103
M2177 3556 VSS 451 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=356280 $Y=511680 $D=103
M2178 452 VSS 3554 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=357140 $Y=511190 $D=103
M2179 3555 VSS 452 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=357140 $Y=511680 $D=103
M2180 577 VSS 4322 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=357480 $Y=511190 $D=103
M2181 4323 VSS 577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=357480 $Y=511680 $D=103
M2182 578 VSS 4321 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=358340 $Y=511190 $D=103
M2183 4324 VSS 578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=358340 $Y=511680 $D=103
M2184 703 VSS 4573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=358680 $Y=511190 $D=103
M2185 4576 VSS 703 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=358680 $Y=511680 $D=103
M2186 704 VSS 4574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=359540 $Y=511190 $D=103
M2187 4575 VSS 704 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=359540 $Y=511680 $D=103
M2188 829 VSS 4826 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=359880 $Y=511190 $D=103
M2189 4827 VSS 829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=359880 $Y=511680 $D=103
M2190 830 VSS 4825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=360740 $Y=511190 $D=103
M2191 4828 VSS 830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=360740 $Y=511680 $D=103
M2192 453 VSS 3557 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=361080 $Y=511190 $D=103
M2193 3560 VSS 453 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=361080 $Y=511680 $D=103
M2194 454 VSS 3558 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=361940 $Y=511190 $D=103
M2195 3559 VSS 454 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=361940 $Y=511680 $D=103
M2196 579 VSS 4326 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=362280 $Y=511190 $D=103
M2197 4327 VSS 579 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=362280 $Y=511680 $D=103
M2198 580 VSS 4325 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=363140 $Y=511190 $D=103
M2199 4328 VSS 580 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=363140 $Y=511680 $D=103
M2200 705 VSS 4577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=363480 $Y=511190 $D=103
M2201 4580 VSS 705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=363480 $Y=511680 $D=103
M2202 706 VSS 4578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=364340 $Y=511190 $D=103
M2203 4579 VSS 706 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=364340 $Y=511680 $D=103
M2204 831 VSS 4830 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=364680 $Y=511190 $D=103
M2205 4831 VSS 831 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=364680 $Y=511680 $D=103
M2206 832 VSS 4829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=365540 $Y=511190 $D=103
M2207 4832 VSS 832 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=365540 $Y=511680 $D=103
M2208 455 VSS 3561 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=365880 $Y=511190 $D=103
M2209 3564 VSS 455 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=365880 $Y=511680 $D=103
M2210 456 VSS 3562 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=366740 $Y=511190 $D=103
M2211 3563 VSS 456 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=366740 $Y=511680 $D=103
M2212 581 VSS 4330 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=367080 $Y=511190 $D=103
M2213 4331 VSS 581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=367080 $Y=511680 $D=103
M2214 582 VSS 4329 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=367940 $Y=511190 $D=103
M2215 4332 VSS 582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=367940 $Y=511680 $D=103
M2216 707 VSS 4581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=368280 $Y=511190 $D=103
M2217 4584 VSS 707 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=368280 $Y=511680 $D=103
M2218 708 VSS 4582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=369140 $Y=511190 $D=103
M2219 4583 VSS 708 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=369140 $Y=511680 $D=103
M2220 833 VSS 4834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=369480 $Y=511190 $D=103
M2221 4835 VSS 833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=369480 $Y=511680 $D=103
M2222 834 VSS 4833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=370340 $Y=511190 $D=103
M2223 4836 VSS 834 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=370340 $Y=511680 $D=103
M2224 457 VSS 3565 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=370680 $Y=511190 $D=103
M2225 3568 VSS 457 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=370680 $Y=511680 $D=103
M2226 458 VSS 3566 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=371540 $Y=511190 $D=103
M2227 3567 VSS 458 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=371540 $Y=511680 $D=103
M2228 583 VSS 4334 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=371880 $Y=511190 $D=103
M2229 4335 VSS 583 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=371880 $Y=511680 $D=103
M2230 584 VSS 4333 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=372740 $Y=511190 $D=103
M2231 4336 VSS 584 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=372740 $Y=511680 $D=103
M2232 709 VSS 4585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=373080 $Y=511190 $D=103
M2233 4588 VSS 709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=373080 $Y=511680 $D=103
M2234 710 VSS 4586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=373940 $Y=511190 $D=103
M2235 4587 VSS 710 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=373940 $Y=511680 $D=103
M2236 835 VSS 4838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=374280 $Y=511190 $D=103
M2237 4839 VSS 835 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=374280 $Y=511680 $D=103
M2238 836 VSS 4837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=375140 $Y=511190 $D=103
M2239 4840 VSS 836 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=375140 $Y=511680 $D=103
M2240 459 VSS 3569 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=375480 $Y=511190 $D=103
M2241 3572 VSS 459 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=375480 $Y=511680 $D=103
M2242 460 VSS 3570 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=376340 $Y=511190 $D=103
M2243 3571 VSS 460 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=376340 $Y=511680 $D=103
M2244 585 VSS 4338 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=376680 $Y=511190 $D=103
M2245 4339 VSS 585 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=376680 $Y=511680 $D=103
M2246 586 VSS 4337 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=377540 $Y=511190 $D=103
M2247 4340 VSS 586 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=377540 $Y=511680 $D=103
M2248 711 VSS 4589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=377880 $Y=511190 $D=103
M2249 4592 VSS 711 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=377880 $Y=511680 $D=103
M2250 712 VSS 4590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=378740 $Y=511190 $D=103
M2251 4591 VSS 712 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=378740 $Y=511680 $D=103
M2252 837 VSS 4842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=379080 $Y=511190 $D=103
M2253 4843 VSS 837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=379080 $Y=511680 $D=103
M2254 838 VSS 4841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=379940 $Y=511190 $D=103
M2255 4844 VSS 838 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=379940 $Y=511680 $D=103
M2256 461 VSS 3573 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=380280 $Y=511190 $D=103
M2257 3576 VSS 461 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=380280 $Y=511680 $D=103
M2258 462 VSS 3574 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=381140 $Y=511190 $D=103
M2259 3575 VSS 462 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=381140 $Y=511680 $D=103
M2260 587 VSS 4342 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=381480 $Y=511190 $D=103
M2261 4343 VSS 587 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=381480 $Y=511680 $D=103
M2262 588 VSS 4341 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=382340 $Y=511190 $D=103
M2263 4344 VSS 588 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=382340 $Y=511680 $D=103
M2264 713 VSS 4593 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=382680 $Y=511190 $D=103
M2265 4596 VSS 713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=382680 $Y=511680 $D=103
M2266 714 VSS 4594 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=383540 $Y=511190 $D=103
M2267 4595 VSS 714 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=383540 $Y=511680 $D=103
M2268 839 VSS 4846 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=383880 $Y=511190 $D=103
M2269 4847 VSS 839 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=383880 $Y=511680 $D=103
M2270 840 VSS 4845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=384740 $Y=511190 $D=103
M2271 4848 VSS 840 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=384740 $Y=511680 $D=103
M2272 463 VSS 3577 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=385080 $Y=511190 $D=103
M2273 3580 VSS 463 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=385080 $Y=511680 $D=103
M2274 464 VSS 3578 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=385940 $Y=511190 $D=103
M2275 3579 VSS 464 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=385940 $Y=511680 $D=103
M2276 589 VSS 4346 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=386280 $Y=511190 $D=103
M2277 4347 VSS 589 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=386280 $Y=511680 $D=103
M2278 590 VSS 4345 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=387140 $Y=511190 $D=103
M2279 4348 VSS 590 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=387140 $Y=511680 $D=103
M2280 715 VSS 4597 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=387480 $Y=511190 $D=103
M2281 4600 VSS 715 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=387480 $Y=511680 $D=103
M2282 716 VSS 4598 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=388340 $Y=511190 $D=103
M2283 4599 VSS 716 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=388340 $Y=511680 $D=103
M2284 841 VSS 4850 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=388680 $Y=511190 $D=103
M2285 4851 VSS 841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=388680 $Y=511680 $D=103
M2286 842 VSS 4849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=389540 $Y=511190 $D=103
M2287 4852 VSS 842 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=389540 $Y=511680 $D=103
M2288 465 VSS 3581 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=389880 $Y=511190 $D=103
M2289 3584 VSS 465 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=389880 $Y=511680 $D=103
M2290 466 VSS 3582 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=390740 $Y=511190 $D=103
M2291 3583 VSS 466 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=390740 $Y=511680 $D=103
M2292 591 VSS 4350 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=391080 $Y=511190 $D=103
M2293 4351 VSS 591 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=391080 $Y=511680 $D=103
M2294 592 VSS 4349 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=391940 $Y=511190 $D=103
M2295 4352 VSS 592 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=391940 $Y=511680 $D=103
M2296 717 VSS 4601 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=392280 $Y=511190 $D=103
M2297 4604 VSS 717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=392280 $Y=511680 $D=103
M2298 718 VSS 4602 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=393140 $Y=511190 $D=103
M2299 4603 VSS 718 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=393140 $Y=511680 $D=103
M2300 843 VSS 4854 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=393480 $Y=511190 $D=103
M2301 4855 VSS 843 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=393480 $Y=511680 $D=103
M2302 5375 63 5633 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=74950 $D=103
M2303 5634 64 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=75440 $D=103
M2304 5375 65 5635 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=78350 $D=103
M2305 5636 66 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=78840 $D=103
M2306 5375 67 5637 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=81750 $D=103
M2307 5638 68 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=82240 $D=103
M2308 5375 69 5639 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=85150 $D=103
M2309 5640 70 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=85640 $D=103
M2310 5375 71 5641 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=88550 $D=103
M2311 5642 72 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=89040 $D=103
M2312 5375 73 5643 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=91950 $D=103
M2313 5644 74 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=92440 $D=103
M2314 5375 75 5645 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=95350 $D=103
M2315 5646 76 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=95840 $D=103
M2316 5375 77 5647 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=98750 $D=103
M2317 5648 78 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=99240 $D=103
M2318 5375 79 5649 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=102150 $D=103
M2319 5650 80 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=102640 $D=103
M2320 5375 81 5651 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=105550 $D=103
M2321 5652 82 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=106040 $D=103
M2322 5375 83 5653 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=108950 $D=103
M2323 5654 84 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=109440 $D=103
M2324 5375 85 5655 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=112350 $D=103
M2325 5656 86 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=112840 $D=103
M2326 5375 87 5657 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=115750 $D=103
M2327 5658 88 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=116240 $D=103
M2328 5375 89 5659 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=119150 $D=103
M2329 5660 90 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=119640 $D=103
M2330 5375 91 5661 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=122550 $D=103
M2331 5662 92 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=123040 $D=103
M2332 5375 93 5663 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=125950 $D=103
M2333 5664 94 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=126440 $D=103
M2334 5375 95 5665 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=129350 $D=103
M2335 5666 96 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=129840 $D=103
M2336 5375 97 5667 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=132750 $D=103
M2337 5668 98 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=133240 $D=103
M2338 5375 99 5669 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=136150 $D=103
M2339 5670 100 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=136640 $D=103
M2340 5375 101 5671 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=139550 $D=103
M2341 5672 102 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=140040 $D=103
M2342 5375 103 5673 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=142950 $D=103
M2343 5674 104 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=143440 $D=103
M2344 5375 105 5675 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=146350 $D=103
M2345 5676 106 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=146840 $D=103
M2346 5375 107 5677 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=149750 $D=103
M2347 5678 108 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=150240 $D=103
M2348 5375 109 5679 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=153150 $D=103
M2349 5680 110 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=153640 $D=103
M2350 5375 111 5681 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=156550 $D=103
M2351 5682 112 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=157040 $D=103
M2352 5375 113 5683 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=159950 $D=103
M2353 5684 114 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=160440 $D=103
M2354 5375 115 5685 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=163350 $D=103
M2355 5686 116 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=163840 $D=103
M2356 5375 117 5687 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=166750 $D=103
M2357 5688 118 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=167240 $D=103
M2358 5375 119 5689 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=170150 $D=103
M2359 5690 120 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=170640 $D=103
M2360 5375 121 5691 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=173550 $D=103
M2361 5692 122 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=174040 $D=103
M2362 5375 123 5693 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=176950 $D=103
M2363 5694 124 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=177440 $D=103
M2364 5375 125 5695 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=180350 $D=103
M2365 5696 126 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=180840 $D=103
M2366 5375 127 5697 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=183750 $D=103
M2367 5698 128 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=184240 $D=103
M2368 5375 129 5699 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=187150 $D=103
M2369 5700 130 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=187640 $D=103
M2370 5375 131 5701 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=190550 $D=103
M2371 5702 132 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=191040 $D=103
M2372 5375 133 5703 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=193950 $D=103
M2373 5704 134 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=194440 $D=103
M2374 5375 135 5705 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=197350 $D=103
M2375 5706 136 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=197840 $D=103
M2376 5375 137 5707 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=200750 $D=103
M2377 5708 138 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=201240 $D=103
M2378 5375 139 5709 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=204150 $D=103
M2379 5710 140 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=204640 $D=103
M2380 5375 141 5711 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=207550 $D=103
M2381 5712 142 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=208040 $D=103
M2382 5375 143 5713 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=210950 $D=103
M2383 5714 144 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=211440 $D=103
M2384 5375 145 5715 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=214350 $D=103
M2385 5716 146 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=214840 $D=103
M2386 5375 147 5717 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=217750 $D=103
M2387 5718 148 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=218240 $D=103
M2388 5375 149 5719 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=221150 $D=103
M2389 5720 150 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=221640 $D=103
M2390 5375 151 5721 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=224550 $D=103
M2391 5722 152 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=225040 $D=103
M2392 5375 153 5723 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=227950 $D=103
M2393 5724 154 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=228440 $D=103
M2394 5375 155 5725 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=231350 $D=103
M2395 5726 156 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=231840 $D=103
M2396 5375 157 5727 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=234750 $D=103
M2397 5728 158 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=235240 $D=103
M2398 5375 159 5729 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=238150 $D=103
M2399 5730 160 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=238640 $D=103
M2400 5375 161 5731 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=241550 $D=103
M2401 5732 162 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=242040 $D=103
M2402 5375 163 5733 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=244950 $D=103
M2403 5734 164 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=245440 $D=103
M2404 5375 165 5735 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=248350 $D=103
M2405 5736 166 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=248840 $D=103
M2406 5375 167 5737 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=251750 $D=103
M2407 5738 168 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=252240 $D=103
M2408 5375 169 5739 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=255150 $D=103
M2409 5740 170 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=255640 $D=103
M2410 5375 171 5741 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=258550 $D=103
M2411 5742 172 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=259040 $D=103
M2412 5375 173 5743 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=261950 $D=103
M2413 5744 174 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=262440 $D=103
M2414 5375 175 5745 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=265350 $D=103
M2415 5746 176 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=265840 $D=103
M2416 5375 177 5747 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=268750 $D=103
M2417 5748 178 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=269240 $D=103
M2418 5375 179 5749 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=272150 $D=103
M2419 5750 180 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=272640 $D=103
M2420 5375 181 5751 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=275550 $D=103
M2421 5752 182 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=276040 $D=103
M2422 5375 183 5753 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=278950 $D=103
M2423 5754 184 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=279440 $D=103
M2424 5375 185 5755 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=282350 $D=103
M2425 5756 186 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=282840 $D=103
M2426 5375 187 5757 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=285750 $D=103
M2427 5758 188 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=286240 $D=103
M2428 5375 189 5759 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=289150 $D=103
M2429 5760 190 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=289640 $D=103
M2430 5375 191 5761 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=292550 $D=103
M2431 5762 192 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=293040 $D=103
M2432 5375 193 5763 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=295950 $D=103
M2433 5764 194 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=296440 $D=103
M2434 5375 195 5765 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=299350 $D=103
M2435 5766 196 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=299840 $D=103
M2436 5375 197 5767 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=302750 $D=103
M2437 5768 198 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=303240 $D=103
M2438 5375 199 5769 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=306150 $D=103
M2439 5770 200 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=306640 $D=103
M2440 5375 201 5771 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=309550 $D=103
M2441 5772 202 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=310040 $D=103
M2442 5375 203 5773 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=312950 $D=103
M2443 5774 204 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=313440 $D=103
M2444 5375 205 5775 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=316350 $D=103
M2445 5776 206 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=316840 $D=103
M2446 5375 207 5777 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=319750 $D=103
M2447 5778 208 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=320240 $D=103
M2448 5375 209 5779 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=323150 $D=103
M2449 5780 210 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=323640 $D=103
M2450 5375 211 5781 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=326550 $D=103
M2451 5782 212 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=327040 $D=103
M2452 5375 213 5783 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=329950 $D=103
M2453 5784 214 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=330440 $D=103
M2454 5375 215 5785 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=333350 $D=103
M2455 5786 216 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=333840 $D=103
M2456 5375 217 5787 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=336750 $D=103
M2457 5788 218 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=337240 $D=103
M2458 5375 219 5789 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=340150 $D=103
M2459 5790 220 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=340640 $D=103
M2460 5375 221 5791 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=343550 $D=103
M2461 5792 222 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=344040 $D=103
M2462 5375 223 5793 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=346950 $D=103
M2463 5794 224 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=347440 $D=103
M2464 5375 225 5795 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=350350 $D=103
M2465 5796 226 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=350840 $D=103
M2466 5375 227 5797 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=353750 $D=103
M2467 5798 228 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=354240 $D=103
M2468 5375 229 5799 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=357150 $D=103
M2469 5800 230 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=357640 $D=103
M2470 5375 231 5801 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=360550 $D=103
M2471 5802 232 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=361040 $D=103
M2472 5375 233 5803 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=363950 $D=103
M2473 5804 234 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=364440 $D=103
M2474 5375 235 5805 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=367350 $D=103
M2475 5806 236 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=367840 $D=103
M2476 5375 237 5807 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=370750 $D=103
M2477 5808 238 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=371240 $D=103
M2478 5375 239 5809 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=374150 $D=103
M2479 5810 240 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=374640 $D=103
M2480 5375 241 5811 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=377550 $D=103
M2481 5812 242 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=378040 $D=103
M2482 5375 243 5813 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=380950 $D=103
M2483 5814 244 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=381440 $D=103
M2484 5375 245 5815 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=384350 $D=103
M2485 5816 246 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=384840 $D=103
M2486 5375 247 5817 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=387750 $D=103
M2487 5818 248 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=388240 $D=103
M2488 5375 249 5819 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=391150 $D=103
M2489 5820 250 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=391640 $D=103
M2490 5375 251 5821 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=394550 $D=103
M2491 5822 252 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=395040 $D=103
M2492 5375 253 5823 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=397950 $D=103
M2493 5824 254 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=398440 $D=103
M2494 5375 255 5825 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=401350 $D=103
M2495 5826 256 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=401840 $D=103
M2496 5375 257 5827 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=404750 $D=103
M2497 5828 258 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=405240 $D=103
M2498 5375 259 5829 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=408150 $D=103
M2499 5830 260 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=408640 $D=103
M2500 5375 261 5831 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=411550 $D=103
M2501 5832 262 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=412040 $D=103
M2502 5375 263 5833 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=414950 $D=103
M2503 5834 264 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=415440 $D=103
M2504 5375 265 5835 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=418350 $D=103
M2505 5836 266 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=418840 $D=103
M2506 5375 267 5837 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=421750 $D=103
M2507 5838 268 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=422240 $D=103
M2508 5375 269 5839 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=425150 $D=103
M2509 5840 270 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=425640 $D=103
M2510 5375 271 5841 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=428550 $D=103
M2511 5842 272 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=429040 $D=103
M2512 5375 273 5843 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=431950 $D=103
M2513 5844 274 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=432440 $D=103
M2514 5375 275 5845 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=435350 $D=103
M2515 5846 276 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=435840 $D=103
M2516 5375 277 5847 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=438750 $D=103
M2517 5848 278 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=439240 $D=103
M2518 5375 279 5849 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=442150 $D=103
M2519 5850 280 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=442640 $D=103
M2520 5375 281 5851 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=445550 $D=103
M2521 5852 282 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=446040 $D=103
M2522 5375 283 5853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=448950 $D=103
M2523 5854 284 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=449440 $D=103
M2524 5375 285 5855 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=452350 $D=103
M2525 5856 286 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=452840 $D=103
M2526 5375 287 5857 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=455750 $D=103
M2527 5858 288 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=456240 $D=103
M2528 5375 289 5859 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=459150 $D=103
M2529 5860 290 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=459640 $D=103
M2530 5375 291 5861 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=462550 $D=103
M2531 5862 292 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=463040 $D=103
M2532 5375 293 5863 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=465950 $D=103
M2533 5864 294 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=466440 $D=103
M2534 5375 295 5865 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=469350 $D=103
M2535 5866 296 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=469840 $D=103
M2536 5375 297 5867 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=472750 $D=103
M2537 5868 298 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=473240 $D=103
M2538 5375 299 5869 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=476150 $D=103
M2539 5870 300 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=476640 $D=103
M2540 5375 301 5871 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=479550 $D=103
M2541 5872 302 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=480040 $D=103
M2542 5375 303 5873 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=482950 $D=103
M2543 5874 304 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=483440 $D=103
M2544 5375 305 5875 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=486350 $D=103
M2545 5876 306 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=486840 $D=103
M2546 5375 307 5877 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=489750 $D=103
M2547 5878 308 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=490240 $D=103
M2548 5375 309 5879 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=493150 $D=103
M2549 5880 310 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=493640 $D=103
M2550 5375 311 5881 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=496550 $D=103
M2551 5882 312 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=497040 $D=103
M2552 5375 313 5883 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=499950 $D=103
M2553 5884 314 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=500440 $D=103
M2554 5375 315 5885 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=503350 $D=103
M2555 5886 316 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=503840 $D=103
M2556 5375 317 5887 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=506750 $D=103
M2557 5888 318 5375 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=507240 $D=103
M2558 844 VSS 4853 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=511190 $D=103
M2559 4856 VSS 844 VSS lpnfet w=1.6e-07 l=1.3e-07 m=1 par=1 nf=1 ngcon=1 $X=394340 $Y=511680 $D=103
D2560 VSS 324 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=48230 $D=558
D2561 VSS 325 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=48830 $D=558
D2562 VSS 326 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=49430 $D=558
D2563 VSS 327 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=50030 $D=558
D2564 VSS 328 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=50630 $D=558
D2565 VSS 329 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=51230 $D=558
D2566 VSS 330 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=51830 $D=558
D2567 VSS 331 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=52430 $D=558
D2568 VSS 332 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=53030 $D=558
D2569 VSS 333 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=234850 $Y=53630 $D=558
D2570 VSS 51 tdndsx AREA=1.024e-13 perim=1.28e-06 $X=235610 $Y=55940 $D=558
X2571 VSS 323 VSS 51 SIGN_MEMFCIO8 $T=12410 10240 1 180 $X=9240 $Y=9240
X2572 VSS 323 VSS 51 SIGN_MEMFCIO8 $T=394590 10240 0 0 $X=393590 $Y=9240
X2573 VSS 51 SIGN_MEMFCSA8 $T=12410 22710 1 180 $X=9240 $Y=21710
X2574 VSS 51 SIGN_MEMFCSA8 $T=394590 22710 0 0 $X=393590 $Y=21710
X2837 VSS VSS 861 SIGN_MEMFLCCSTRAPR $T=12410 509800 1 180 $X=10210 $Y=508800
X2838 VSS VSS 861 SIGN_MEMFLCCSTRAPR $T=12410 513200 0 180 $X=10210 $Y=510500
X2839 VSS 50 862 SIGN_MEMFLCCSTRAPR $T=169610 509800 0 0 $X=168610 $Y=508800
X2840 VSS 50 862 SIGN_MEMFLCCSTRAPR $T=169610 513200 1 0 $X=168610 $Y=510500
X2841 VSS VSS 863 SIGN_MEMFLCCSTRAPR $T=394590 509800 0 0 $X=393590 $Y=508800
X2842 VSS VSS 863 SIGN_MEMFLCCSTRAPR $T=394590 513200 1 0 $X=393590 $Y=510500
X2843 VSS 63 64 ICV_42 $T=12410 73560 1 180 $X=10210 $Y=72560
X2844 VSS 65 66 ICV_42 $T=12410 76960 1 180 $X=10210 $Y=75960
X2845 VSS 67 68 ICV_42 $T=12410 80360 1 180 $X=10210 $Y=79360
X2846 VSS 69 70 ICV_42 $T=12410 83760 1 180 $X=10210 $Y=82760
X2847 VSS 71 72 ICV_42 $T=12410 87160 1 180 $X=10210 $Y=86160
X2848 VSS 73 74 ICV_42 $T=12410 90560 1 180 $X=10210 $Y=89560
X2849 VSS 75 76 ICV_42 $T=12410 93960 1 180 $X=10210 $Y=92960
X2850 VSS 77 78 ICV_42 $T=12410 97360 1 180 $X=10210 $Y=96360
X2851 VSS 79 80 ICV_42 $T=12410 100760 1 180 $X=10210 $Y=99760
X2852 VSS 81 82 ICV_42 $T=12410 104160 1 180 $X=10210 $Y=103160
X2853 VSS 83 84 ICV_42 $T=12410 107560 1 180 $X=10210 $Y=106560
X2854 VSS 85 86 ICV_42 $T=12410 110960 1 180 $X=10210 $Y=109960
X2855 VSS 87 88 ICV_42 $T=12410 114360 1 180 $X=10210 $Y=113360
X2856 VSS 89 90 ICV_42 $T=12410 117760 1 180 $X=10210 $Y=116760
X2857 VSS 91 92 ICV_42 $T=12410 121160 1 180 $X=10210 $Y=120160
X2858 VSS 93 94 ICV_42 $T=12410 124560 1 180 $X=10210 $Y=123560
X2859 VSS 95 96 ICV_42 $T=12410 127960 1 180 $X=10210 $Y=126960
X2860 VSS 97 98 ICV_42 $T=12410 131360 1 180 $X=10210 $Y=130360
X2861 VSS 99 100 ICV_42 $T=12410 134760 1 180 $X=10210 $Y=133760
X2862 VSS 101 102 ICV_42 $T=12410 138160 1 180 $X=10210 $Y=137160
X2863 VSS 103 104 ICV_42 $T=12410 141560 1 180 $X=10210 $Y=140560
X2864 VSS 105 106 ICV_42 $T=12410 144960 1 180 $X=10210 $Y=143960
X2865 VSS 107 108 ICV_42 $T=12410 148360 1 180 $X=10210 $Y=147360
X2866 VSS 109 110 ICV_42 $T=12410 151760 1 180 $X=10210 $Y=150760
X2867 VSS 111 112 ICV_42 $T=12410 155160 1 180 $X=10210 $Y=154160
X2868 VSS 113 114 ICV_42 $T=12410 158560 1 180 $X=10210 $Y=157560
X2869 VSS 115 116 ICV_42 $T=12410 161960 1 180 $X=10210 $Y=160960
X2870 VSS 117 118 ICV_42 $T=12410 165360 1 180 $X=10210 $Y=164360
X2871 VSS 119 120 ICV_42 $T=12410 168760 1 180 $X=10210 $Y=167760
X2872 VSS 121 122 ICV_42 $T=12410 172160 1 180 $X=10210 $Y=171160
X2873 VSS 123 124 ICV_42 $T=12410 175560 1 180 $X=10210 $Y=174560
X2874 VSS 125 126 ICV_42 $T=12410 178960 1 180 $X=10210 $Y=177960
X2875 VSS 127 128 ICV_42 $T=12410 182360 1 180 $X=10210 $Y=181360
X2876 VSS 129 130 ICV_42 $T=12410 185760 1 180 $X=10210 $Y=184760
X2877 VSS 131 132 ICV_42 $T=12410 189160 1 180 $X=10210 $Y=188160
X2878 VSS 133 134 ICV_42 $T=12410 192560 1 180 $X=10210 $Y=191560
X2879 VSS 135 136 ICV_42 $T=12410 195960 1 180 $X=10210 $Y=194960
X2880 VSS 137 138 ICV_42 $T=12410 199360 1 180 $X=10210 $Y=198360
X2881 VSS 139 140 ICV_42 $T=12410 202760 1 180 $X=10210 $Y=201760
X2882 VSS 141 142 ICV_42 $T=12410 206160 1 180 $X=10210 $Y=205160
X2883 VSS 143 144 ICV_42 $T=12410 209560 1 180 $X=10210 $Y=208560
X2884 VSS 145 146 ICV_42 $T=12410 212960 1 180 $X=10210 $Y=211960
X2885 VSS 147 148 ICV_42 $T=12410 216360 1 180 $X=10210 $Y=215360
X2886 VSS 149 150 ICV_42 $T=12410 219760 1 180 $X=10210 $Y=218760
X2887 VSS 151 152 ICV_42 $T=12410 223160 1 180 $X=10210 $Y=222160
X2888 VSS 153 154 ICV_42 $T=12410 226560 1 180 $X=10210 $Y=225560
X2889 VSS 155 156 ICV_42 $T=12410 229960 1 180 $X=10210 $Y=228960
X2890 VSS 157 158 ICV_42 $T=12410 233360 1 180 $X=10210 $Y=232360
X2891 VSS 159 160 ICV_42 $T=12410 236760 1 180 $X=10210 $Y=235760
X2892 VSS 161 162 ICV_42 $T=12410 240160 1 180 $X=10210 $Y=239160
X2893 VSS 163 164 ICV_42 $T=12410 243560 1 180 $X=10210 $Y=242560
X2894 VSS 165 166 ICV_42 $T=12410 246960 1 180 $X=10210 $Y=245960
X2895 VSS 167 168 ICV_42 $T=12410 250360 1 180 $X=10210 $Y=249360
X2896 VSS 169 170 ICV_42 $T=12410 253760 1 180 $X=10210 $Y=252760
X2897 VSS 171 172 ICV_42 $T=12410 257160 1 180 $X=10210 $Y=256160
X2898 VSS 173 174 ICV_42 $T=12410 260560 1 180 $X=10210 $Y=259560
X2899 VSS 175 176 ICV_42 $T=12410 263960 1 180 $X=10210 $Y=262960
X2900 VSS 177 178 ICV_42 $T=12410 267360 1 180 $X=10210 $Y=266360
X2901 VSS 179 180 ICV_42 $T=12410 270760 1 180 $X=10210 $Y=269760
X2902 VSS 181 182 ICV_42 $T=12410 274160 1 180 $X=10210 $Y=273160
X2903 VSS 183 184 ICV_42 $T=12410 277560 1 180 $X=10210 $Y=276560
X2904 VSS 185 186 ICV_42 $T=12410 280960 1 180 $X=10210 $Y=279960
X2905 VSS 187 188 ICV_42 $T=12410 284360 1 180 $X=10210 $Y=283360
X2906 VSS 189 190 ICV_42 $T=12410 287760 1 180 $X=10210 $Y=286760
X2907 VSS 191 192 ICV_42 $T=12410 291160 1 180 $X=10210 $Y=290160
X2908 VSS 193 194 ICV_42 $T=12410 294560 1 180 $X=10210 $Y=293560
X2909 VSS 195 196 ICV_42 $T=12410 297960 1 180 $X=10210 $Y=296960
X2910 VSS 197 198 ICV_42 $T=12410 301360 1 180 $X=10210 $Y=300360
X2911 VSS 199 200 ICV_42 $T=12410 304760 1 180 $X=10210 $Y=303760
X2912 VSS 201 202 ICV_42 $T=12410 308160 1 180 $X=10210 $Y=307160
X2913 VSS 203 204 ICV_42 $T=12410 311560 1 180 $X=10210 $Y=310560
X2914 VSS 205 206 ICV_42 $T=12410 314960 1 180 $X=10210 $Y=313960
X2915 VSS 207 208 ICV_42 $T=12410 318360 1 180 $X=10210 $Y=317360
X2916 VSS 209 210 ICV_42 $T=12410 321760 1 180 $X=10210 $Y=320760
X2917 VSS 211 212 ICV_42 $T=12410 325160 1 180 $X=10210 $Y=324160
X2918 VSS 213 214 ICV_42 $T=12410 328560 1 180 $X=10210 $Y=327560
X2919 VSS 215 216 ICV_42 $T=12410 331960 1 180 $X=10210 $Y=330960
X2920 VSS 217 218 ICV_42 $T=12410 335360 1 180 $X=10210 $Y=334360
X2921 VSS 219 220 ICV_42 $T=12410 338760 1 180 $X=10210 $Y=337760
X2922 VSS 221 222 ICV_42 $T=12410 342160 1 180 $X=10210 $Y=341160
X2923 VSS 223 224 ICV_42 $T=12410 345560 1 180 $X=10210 $Y=344560
X2924 VSS 225 226 ICV_42 $T=12410 348960 1 180 $X=10210 $Y=347960
X2925 VSS 227 228 ICV_42 $T=12410 352360 1 180 $X=10210 $Y=351360
X2926 VSS 229 230 ICV_42 $T=12410 355760 1 180 $X=10210 $Y=354760
X2927 VSS 231 232 ICV_42 $T=12410 359160 1 180 $X=10210 $Y=358160
X2928 VSS 233 234 ICV_42 $T=12410 362560 1 180 $X=10210 $Y=361560
X2929 VSS 235 236 ICV_42 $T=12410 365960 1 180 $X=10210 $Y=364960
X2930 VSS 237 238 ICV_42 $T=12410 369360 1 180 $X=10210 $Y=368360
X2931 VSS 239 240 ICV_42 $T=12410 372760 1 180 $X=10210 $Y=371760
X2932 VSS 241 242 ICV_42 $T=12410 376160 1 180 $X=10210 $Y=375160
X2933 VSS 243 244 ICV_42 $T=12410 379560 1 180 $X=10210 $Y=378560
X2934 VSS 245 246 ICV_42 $T=12410 382960 1 180 $X=10210 $Y=381960
X2935 VSS 247 248 ICV_42 $T=12410 386360 1 180 $X=10210 $Y=385360
X2936 VSS 249 250 ICV_42 $T=12410 389760 1 180 $X=10210 $Y=388760
X2937 VSS 251 252 ICV_42 $T=12410 393160 1 180 $X=10210 $Y=392160
X2938 VSS 253 254 ICV_42 $T=12410 396560 1 180 $X=10210 $Y=395560
X2939 VSS 255 256 ICV_42 $T=12410 399960 1 180 $X=10210 $Y=398960
X2940 VSS 257 258 ICV_42 $T=12410 403360 1 180 $X=10210 $Y=402360
X2941 VSS 259 260 ICV_42 $T=12410 406760 1 180 $X=10210 $Y=405760
X2942 VSS 261 262 ICV_42 $T=12410 410160 1 180 $X=10210 $Y=409160
X2943 VSS 263 264 ICV_42 $T=12410 413560 1 180 $X=10210 $Y=412560
X2944 VSS 265 266 ICV_42 $T=12410 416960 1 180 $X=10210 $Y=415960
X2945 VSS 267 268 ICV_42 $T=12410 420360 1 180 $X=10210 $Y=419360
X2946 VSS 269 270 ICV_42 $T=12410 423760 1 180 $X=10210 $Y=422760
X2947 VSS 271 272 ICV_42 $T=12410 427160 1 180 $X=10210 $Y=426160
X2948 VSS 273 274 ICV_42 $T=12410 430560 1 180 $X=10210 $Y=429560
X2949 VSS 275 276 ICV_42 $T=12410 433960 1 180 $X=10210 $Y=432960
X2950 VSS 277 278 ICV_42 $T=12410 437360 1 180 $X=10210 $Y=436360
X2951 VSS 279 280 ICV_42 $T=12410 440760 1 180 $X=10210 $Y=439760
X2952 VSS 281 282 ICV_42 $T=12410 444160 1 180 $X=10210 $Y=443160
X2953 VSS 283 284 ICV_42 $T=12410 447560 1 180 $X=10210 $Y=446560
X2954 VSS 285 286 ICV_42 $T=12410 450960 1 180 $X=10210 $Y=449960
X2955 VSS 287 288 ICV_42 $T=12410 454360 1 180 $X=10210 $Y=453360
X2956 VSS 289 290 ICV_42 $T=12410 457760 1 180 $X=10210 $Y=456760
X2957 VSS 291 292 ICV_42 $T=12410 461160 1 180 $X=10210 $Y=460160
X2958 VSS 293 294 ICV_42 $T=12410 464560 1 180 $X=10210 $Y=463560
X2959 VSS 295 296 ICV_42 $T=12410 467960 1 180 $X=10210 $Y=466960
X2960 VSS 297 298 ICV_42 $T=12410 471360 1 180 $X=10210 $Y=470360
X2961 VSS 299 300 ICV_42 $T=12410 474760 1 180 $X=10210 $Y=473760
X2962 VSS 301 302 ICV_42 $T=12410 478160 1 180 $X=10210 $Y=477160
X2963 VSS 303 304 ICV_42 $T=12410 481560 1 180 $X=10210 $Y=480560
X2964 VSS 305 306 ICV_42 $T=12410 484960 1 180 $X=10210 $Y=483960
X2965 VSS 307 308 ICV_42 $T=12410 488360 1 180 $X=10210 $Y=487360
X2966 VSS 309 310 ICV_42 $T=12410 491760 1 180 $X=10210 $Y=490760
X2967 VSS 311 312 ICV_42 $T=12410 495160 1 180 $X=10210 $Y=494160
X2968 VSS 313 314 ICV_42 $T=12410 498560 1 180 $X=10210 $Y=497560
X2969 VSS 315 316 ICV_42 $T=12410 501960 1 180 $X=10210 $Y=500960
X2970 VSS 317 318 ICV_42 $T=12410 505360 1 180 $X=10210 $Y=504360
X2971 VSS 63 64 ICV_42 $T=169610 73560 0 0 $X=168610 $Y=72560
X2972 VSS 65 66 ICV_42 $T=169610 76960 0 0 $X=168610 $Y=75960
X2973 VSS 67 68 ICV_42 $T=169610 80360 0 0 $X=168610 $Y=79360
X2974 VSS 69 70 ICV_42 $T=169610 83760 0 0 $X=168610 $Y=82760
X2975 VSS 71 72 ICV_42 $T=169610 87160 0 0 $X=168610 $Y=86160
X2976 VSS 73 74 ICV_42 $T=169610 90560 0 0 $X=168610 $Y=89560
X2977 VSS 75 76 ICV_42 $T=169610 93960 0 0 $X=168610 $Y=92960
X2978 VSS 77 78 ICV_42 $T=169610 97360 0 0 $X=168610 $Y=96360
X2979 VSS 79 80 ICV_42 $T=169610 100760 0 0 $X=168610 $Y=99760
X2980 VSS 81 82 ICV_42 $T=169610 104160 0 0 $X=168610 $Y=103160
X2981 VSS 83 84 ICV_42 $T=169610 107560 0 0 $X=168610 $Y=106560
X2982 VSS 85 86 ICV_42 $T=169610 110960 0 0 $X=168610 $Y=109960
X2983 VSS 87 88 ICV_42 $T=169610 114360 0 0 $X=168610 $Y=113360
X2984 VSS 89 90 ICV_42 $T=169610 117760 0 0 $X=168610 $Y=116760
X2985 VSS 91 92 ICV_42 $T=169610 121160 0 0 $X=168610 $Y=120160
X2986 VSS 93 94 ICV_42 $T=169610 124560 0 0 $X=168610 $Y=123560
X2987 VSS 95 96 ICV_42 $T=169610 127960 0 0 $X=168610 $Y=126960
X2988 VSS 97 98 ICV_42 $T=169610 131360 0 0 $X=168610 $Y=130360
X2989 VSS 99 100 ICV_42 $T=169610 134760 0 0 $X=168610 $Y=133760
X2990 VSS 101 102 ICV_42 $T=169610 138160 0 0 $X=168610 $Y=137160
X2991 VSS 103 104 ICV_42 $T=169610 141560 0 0 $X=168610 $Y=140560
X2992 VSS 105 106 ICV_42 $T=169610 144960 0 0 $X=168610 $Y=143960
X2993 VSS 107 108 ICV_42 $T=169610 148360 0 0 $X=168610 $Y=147360
X2994 VSS 109 110 ICV_42 $T=169610 151760 0 0 $X=168610 $Y=150760
X2995 VSS 111 112 ICV_42 $T=169610 155160 0 0 $X=168610 $Y=154160
X2996 VSS 113 114 ICV_42 $T=169610 158560 0 0 $X=168610 $Y=157560
X2997 VSS 115 116 ICV_42 $T=169610 161960 0 0 $X=168610 $Y=160960
X2998 VSS 117 118 ICV_42 $T=169610 165360 0 0 $X=168610 $Y=164360
X2999 VSS 119 120 ICV_42 $T=169610 168760 0 0 $X=168610 $Y=167760
X3000 VSS 121 122 ICV_42 $T=169610 172160 0 0 $X=168610 $Y=171160
X3001 VSS 123 124 ICV_42 $T=169610 175560 0 0 $X=168610 $Y=174560
X3002 VSS 125 126 ICV_42 $T=169610 178960 0 0 $X=168610 $Y=177960
X3003 VSS 127 128 ICV_42 $T=169610 182360 0 0 $X=168610 $Y=181360
X3004 VSS 129 130 ICV_42 $T=169610 185760 0 0 $X=168610 $Y=184760
X3005 VSS 131 132 ICV_42 $T=169610 189160 0 0 $X=168610 $Y=188160
X3006 VSS 133 134 ICV_42 $T=169610 192560 0 0 $X=168610 $Y=191560
X3007 VSS 135 136 ICV_42 $T=169610 195960 0 0 $X=168610 $Y=194960
X3008 VSS 137 138 ICV_42 $T=169610 199360 0 0 $X=168610 $Y=198360
X3009 VSS 139 140 ICV_42 $T=169610 202760 0 0 $X=168610 $Y=201760
X3010 VSS 141 142 ICV_42 $T=169610 206160 0 0 $X=168610 $Y=205160
X3011 VSS 143 144 ICV_42 $T=169610 209560 0 0 $X=168610 $Y=208560
X3012 VSS 145 146 ICV_42 $T=169610 212960 0 0 $X=168610 $Y=211960
X3013 VSS 147 148 ICV_42 $T=169610 216360 0 0 $X=168610 $Y=215360
X3014 VSS 149 150 ICV_42 $T=169610 219760 0 0 $X=168610 $Y=218760
X3015 VSS 151 152 ICV_42 $T=169610 223160 0 0 $X=168610 $Y=222160
X3016 VSS 153 154 ICV_42 $T=169610 226560 0 0 $X=168610 $Y=225560
X3017 VSS 155 156 ICV_42 $T=169610 229960 0 0 $X=168610 $Y=228960
X3018 VSS 157 158 ICV_42 $T=169610 233360 0 0 $X=168610 $Y=232360
X3019 VSS 159 160 ICV_42 $T=169610 236760 0 0 $X=168610 $Y=235760
X3020 VSS 161 162 ICV_42 $T=169610 240160 0 0 $X=168610 $Y=239160
X3021 VSS 163 164 ICV_42 $T=169610 243560 0 0 $X=168610 $Y=242560
X3022 VSS 165 166 ICV_42 $T=169610 246960 0 0 $X=168610 $Y=245960
X3023 VSS 167 168 ICV_42 $T=169610 250360 0 0 $X=168610 $Y=249360
X3024 VSS 169 170 ICV_42 $T=169610 253760 0 0 $X=168610 $Y=252760
X3025 VSS 171 172 ICV_42 $T=169610 257160 0 0 $X=168610 $Y=256160
X3026 VSS 173 174 ICV_42 $T=169610 260560 0 0 $X=168610 $Y=259560
X3027 VSS 175 176 ICV_42 $T=169610 263960 0 0 $X=168610 $Y=262960
X3028 VSS 177 178 ICV_42 $T=169610 267360 0 0 $X=168610 $Y=266360
X3029 VSS 179 180 ICV_42 $T=169610 270760 0 0 $X=168610 $Y=269760
X3030 VSS 181 182 ICV_42 $T=169610 274160 0 0 $X=168610 $Y=273160
X3031 VSS 183 184 ICV_42 $T=169610 277560 0 0 $X=168610 $Y=276560
X3032 VSS 185 186 ICV_42 $T=169610 280960 0 0 $X=168610 $Y=279960
X3033 VSS 187 188 ICV_42 $T=169610 284360 0 0 $X=168610 $Y=283360
X3034 VSS 189 190 ICV_42 $T=169610 287760 0 0 $X=168610 $Y=286760
X3035 VSS 191 192 ICV_42 $T=169610 291160 0 0 $X=168610 $Y=290160
X3036 VSS 193 194 ICV_42 $T=169610 294560 0 0 $X=168610 $Y=293560
X3037 VSS 195 196 ICV_42 $T=169610 297960 0 0 $X=168610 $Y=296960
X3038 VSS 197 198 ICV_42 $T=169610 301360 0 0 $X=168610 $Y=300360
X3039 VSS 199 200 ICV_42 $T=169610 304760 0 0 $X=168610 $Y=303760
X3040 VSS 201 202 ICV_42 $T=169610 308160 0 0 $X=168610 $Y=307160
X3041 VSS 203 204 ICV_42 $T=169610 311560 0 0 $X=168610 $Y=310560
X3042 VSS 205 206 ICV_42 $T=169610 314960 0 0 $X=168610 $Y=313960
X3043 VSS 207 208 ICV_42 $T=169610 318360 0 0 $X=168610 $Y=317360
X3044 VSS 209 210 ICV_42 $T=169610 321760 0 0 $X=168610 $Y=320760
X3045 VSS 211 212 ICV_42 $T=169610 325160 0 0 $X=168610 $Y=324160
X3046 VSS 213 214 ICV_42 $T=169610 328560 0 0 $X=168610 $Y=327560
X3047 VSS 215 216 ICV_42 $T=169610 331960 0 0 $X=168610 $Y=330960
X3048 VSS 217 218 ICV_42 $T=169610 335360 0 0 $X=168610 $Y=334360
X3049 VSS 219 220 ICV_42 $T=169610 338760 0 0 $X=168610 $Y=337760
X3050 VSS 221 222 ICV_42 $T=169610 342160 0 0 $X=168610 $Y=341160
X3051 VSS 223 224 ICV_42 $T=169610 345560 0 0 $X=168610 $Y=344560
X3052 VSS 225 226 ICV_42 $T=169610 348960 0 0 $X=168610 $Y=347960
X3053 VSS 227 228 ICV_42 $T=169610 352360 0 0 $X=168610 $Y=351360
X3054 VSS 229 230 ICV_42 $T=169610 355760 0 0 $X=168610 $Y=354760
X3055 VSS 231 232 ICV_42 $T=169610 359160 0 0 $X=168610 $Y=358160
X3056 VSS 233 234 ICV_42 $T=169610 362560 0 0 $X=168610 $Y=361560
X3057 VSS 235 236 ICV_42 $T=169610 365960 0 0 $X=168610 $Y=364960
X3058 VSS 237 238 ICV_42 $T=169610 369360 0 0 $X=168610 $Y=368360
X3059 VSS 239 240 ICV_42 $T=169610 372760 0 0 $X=168610 $Y=371760
X3060 VSS 241 242 ICV_42 $T=169610 376160 0 0 $X=168610 $Y=375160
X3061 VSS 243 244 ICV_42 $T=169610 379560 0 0 $X=168610 $Y=378560
X3062 VSS 245 246 ICV_42 $T=169610 382960 0 0 $X=168610 $Y=381960
X3063 VSS 247 248 ICV_42 $T=169610 386360 0 0 $X=168610 $Y=385360
X3064 VSS 249 250 ICV_42 $T=169610 389760 0 0 $X=168610 $Y=388760
X3065 VSS 251 252 ICV_42 $T=169610 393160 0 0 $X=168610 $Y=392160
X3066 VSS 253 254 ICV_42 $T=169610 396560 0 0 $X=168610 $Y=395560
X3067 VSS 255 256 ICV_42 $T=169610 399960 0 0 $X=168610 $Y=398960
X3068 VSS 257 258 ICV_42 $T=169610 403360 0 0 $X=168610 $Y=402360
X3069 VSS 259 260 ICV_42 $T=169610 406760 0 0 $X=168610 $Y=405760
X3070 VSS 261 262 ICV_42 $T=169610 410160 0 0 $X=168610 $Y=409160
X3071 VSS 263 264 ICV_42 $T=169610 413560 0 0 $X=168610 $Y=412560
X3072 VSS 265 266 ICV_42 $T=169610 416960 0 0 $X=168610 $Y=415960
X3073 VSS 267 268 ICV_42 $T=169610 420360 0 0 $X=168610 $Y=419360
X3074 VSS 269 270 ICV_42 $T=169610 423760 0 0 $X=168610 $Y=422760
X3075 VSS 271 272 ICV_42 $T=169610 427160 0 0 $X=168610 $Y=426160
X3076 VSS 273 274 ICV_42 $T=169610 430560 0 0 $X=168610 $Y=429560
X3077 VSS 275 276 ICV_42 $T=169610 433960 0 0 $X=168610 $Y=432960
X3078 VSS 277 278 ICV_42 $T=169610 437360 0 0 $X=168610 $Y=436360
X3079 VSS 279 280 ICV_42 $T=169610 440760 0 0 $X=168610 $Y=439760
X3080 VSS 281 282 ICV_42 $T=169610 444160 0 0 $X=168610 $Y=443160
X3081 VSS 283 284 ICV_42 $T=169610 447560 0 0 $X=168610 $Y=446560
X3082 VSS 285 286 ICV_42 $T=169610 450960 0 0 $X=168610 $Y=449960
X3083 VSS 287 288 ICV_42 $T=169610 454360 0 0 $X=168610 $Y=453360
X3084 VSS 289 290 ICV_42 $T=169610 457760 0 0 $X=168610 $Y=456760
X3085 VSS 291 292 ICV_42 $T=169610 461160 0 0 $X=168610 $Y=460160
X3086 VSS 293 294 ICV_42 $T=169610 464560 0 0 $X=168610 $Y=463560
X3087 VSS 295 296 ICV_42 $T=169610 467960 0 0 $X=168610 $Y=466960
X3088 VSS 297 298 ICV_42 $T=169610 471360 0 0 $X=168610 $Y=470360
X3089 VSS 299 300 ICV_42 $T=169610 474760 0 0 $X=168610 $Y=473760
X3090 VSS 301 302 ICV_42 $T=169610 478160 0 0 $X=168610 $Y=477160
X3091 VSS 303 304 ICV_42 $T=169610 481560 0 0 $X=168610 $Y=480560
X3092 VSS 305 306 ICV_42 $T=169610 484960 0 0 $X=168610 $Y=483960
X3093 VSS 307 308 ICV_42 $T=169610 488360 0 0 $X=168610 $Y=487360
X3094 VSS 309 310 ICV_42 $T=169610 491760 0 0 $X=168610 $Y=490760
X3095 VSS 311 312 ICV_42 $T=169610 495160 0 0 $X=168610 $Y=494160
X3096 VSS 313 314 ICV_42 $T=169610 498560 0 0 $X=168610 $Y=497560
X3097 VSS 315 316 ICV_42 $T=169610 501960 0 0 $X=168610 $Y=500960
X3098 VSS 317 318 ICV_42 $T=169610 505360 0 0 $X=168610 $Y=504360
X3099 VSS 63 64 ICV_42 $T=394590 73560 0 0 $X=393590 $Y=72560
X3100 VSS 65 66 ICV_42 $T=394590 76960 0 0 $X=393590 $Y=75960
X3101 VSS 67 68 ICV_42 $T=394590 80360 0 0 $X=393590 $Y=79360
X3102 VSS 69 70 ICV_42 $T=394590 83760 0 0 $X=393590 $Y=82760
X3103 VSS 71 72 ICV_42 $T=394590 87160 0 0 $X=393590 $Y=86160
X3104 VSS 73 74 ICV_42 $T=394590 90560 0 0 $X=393590 $Y=89560
X3105 VSS 75 76 ICV_42 $T=394590 93960 0 0 $X=393590 $Y=92960
X3106 VSS 77 78 ICV_42 $T=394590 97360 0 0 $X=393590 $Y=96360
X3107 VSS 79 80 ICV_42 $T=394590 100760 0 0 $X=393590 $Y=99760
X3108 VSS 81 82 ICV_42 $T=394590 104160 0 0 $X=393590 $Y=103160
X3109 VSS 83 84 ICV_42 $T=394590 107560 0 0 $X=393590 $Y=106560
X3110 VSS 85 86 ICV_42 $T=394590 110960 0 0 $X=393590 $Y=109960
X3111 VSS 87 88 ICV_42 $T=394590 114360 0 0 $X=393590 $Y=113360
X3112 VSS 89 90 ICV_42 $T=394590 117760 0 0 $X=393590 $Y=116760
X3113 VSS 91 92 ICV_42 $T=394590 121160 0 0 $X=393590 $Y=120160
X3114 VSS 93 94 ICV_42 $T=394590 124560 0 0 $X=393590 $Y=123560
X3115 VSS 95 96 ICV_42 $T=394590 127960 0 0 $X=393590 $Y=126960
X3116 VSS 97 98 ICV_42 $T=394590 131360 0 0 $X=393590 $Y=130360
X3117 VSS 99 100 ICV_42 $T=394590 134760 0 0 $X=393590 $Y=133760
X3118 VSS 101 102 ICV_42 $T=394590 138160 0 0 $X=393590 $Y=137160
X3119 VSS 103 104 ICV_42 $T=394590 141560 0 0 $X=393590 $Y=140560
X3120 VSS 105 106 ICV_42 $T=394590 144960 0 0 $X=393590 $Y=143960
X3121 VSS 107 108 ICV_42 $T=394590 148360 0 0 $X=393590 $Y=147360
X3122 VSS 109 110 ICV_42 $T=394590 151760 0 0 $X=393590 $Y=150760
X3123 VSS 111 112 ICV_42 $T=394590 155160 0 0 $X=393590 $Y=154160
X3124 VSS 113 114 ICV_42 $T=394590 158560 0 0 $X=393590 $Y=157560
X3125 VSS 115 116 ICV_42 $T=394590 161960 0 0 $X=393590 $Y=160960
X3126 VSS 117 118 ICV_42 $T=394590 165360 0 0 $X=393590 $Y=164360
X3127 VSS 119 120 ICV_42 $T=394590 168760 0 0 $X=393590 $Y=167760
X3128 VSS 121 122 ICV_42 $T=394590 172160 0 0 $X=393590 $Y=171160
X3129 VSS 123 124 ICV_42 $T=394590 175560 0 0 $X=393590 $Y=174560
X3130 VSS 125 126 ICV_42 $T=394590 178960 0 0 $X=393590 $Y=177960
X3131 VSS 127 128 ICV_42 $T=394590 182360 0 0 $X=393590 $Y=181360
X3132 VSS 129 130 ICV_42 $T=394590 185760 0 0 $X=393590 $Y=184760
X3133 VSS 131 132 ICV_42 $T=394590 189160 0 0 $X=393590 $Y=188160
X3134 VSS 133 134 ICV_42 $T=394590 192560 0 0 $X=393590 $Y=191560
X3135 VSS 135 136 ICV_42 $T=394590 195960 0 0 $X=393590 $Y=194960
X3136 VSS 137 138 ICV_42 $T=394590 199360 0 0 $X=393590 $Y=198360
X3137 VSS 139 140 ICV_42 $T=394590 202760 0 0 $X=393590 $Y=201760
X3138 VSS 141 142 ICV_42 $T=394590 206160 0 0 $X=393590 $Y=205160
X3139 VSS 143 144 ICV_42 $T=394590 209560 0 0 $X=393590 $Y=208560
X3140 VSS 145 146 ICV_42 $T=394590 212960 0 0 $X=393590 $Y=211960
X3141 VSS 147 148 ICV_42 $T=394590 216360 0 0 $X=393590 $Y=215360
X3142 VSS 149 150 ICV_42 $T=394590 219760 0 0 $X=393590 $Y=218760
X3143 VSS 151 152 ICV_42 $T=394590 223160 0 0 $X=393590 $Y=222160
X3144 VSS 153 154 ICV_42 $T=394590 226560 0 0 $X=393590 $Y=225560
X3145 VSS 155 156 ICV_42 $T=394590 229960 0 0 $X=393590 $Y=228960
X3146 VSS 157 158 ICV_42 $T=394590 233360 0 0 $X=393590 $Y=232360
X3147 VSS 159 160 ICV_42 $T=394590 236760 0 0 $X=393590 $Y=235760
X3148 VSS 161 162 ICV_42 $T=394590 240160 0 0 $X=393590 $Y=239160
X3149 VSS 163 164 ICV_42 $T=394590 243560 0 0 $X=393590 $Y=242560
X3150 VSS 165 166 ICV_42 $T=394590 246960 0 0 $X=393590 $Y=245960
X3151 VSS 167 168 ICV_42 $T=394590 250360 0 0 $X=393590 $Y=249360
X3152 VSS 169 170 ICV_42 $T=394590 253760 0 0 $X=393590 $Y=252760
X3153 VSS 171 172 ICV_42 $T=394590 257160 0 0 $X=393590 $Y=256160
X3154 VSS 173 174 ICV_42 $T=394590 260560 0 0 $X=393590 $Y=259560
X3155 VSS 175 176 ICV_42 $T=394590 263960 0 0 $X=393590 $Y=262960
X3156 VSS 177 178 ICV_42 $T=394590 267360 0 0 $X=393590 $Y=266360
X3157 VSS 179 180 ICV_42 $T=394590 270760 0 0 $X=393590 $Y=269760
X3158 VSS 181 182 ICV_42 $T=394590 274160 0 0 $X=393590 $Y=273160
X3159 VSS 183 184 ICV_42 $T=394590 277560 0 0 $X=393590 $Y=276560
X3160 VSS 185 186 ICV_42 $T=394590 280960 0 0 $X=393590 $Y=279960
X3161 VSS 187 188 ICV_42 $T=394590 284360 0 0 $X=393590 $Y=283360
X3162 VSS 189 190 ICV_42 $T=394590 287760 0 0 $X=393590 $Y=286760
X3163 VSS 191 192 ICV_42 $T=394590 291160 0 0 $X=393590 $Y=290160
X3164 VSS 193 194 ICV_42 $T=394590 294560 0 0 $X=393590 $Y=293560
X3165 VSS 195 196 ICV_42 $T=394590 297960 0 0 $X=393590 $Y=296960
X3166 VSS 197 198 ICV_42 $T=394590 301360 0 0 $X=393590 $Y=300360
X3167 VSS 199 200 ICV_42 $T=394590 304760 0 0 $X=393590 $Y=303760
X3168 VSS 201 202 ICV_42 $T=394590 308160 0 0 $X=393590 $Y=307160
X3169 VSS 203 204 ICV_42 $T=394590 311560 0 0 $X=393590 $Y=310560
X3170 VSS 205 206 ICV_42 $T=394590 314960 0 0 $X=393590 $Y=313960
X3171 VSS 207 208 ICV_42 $T=394590 318360 0 0 $X=393590 $Y=317360
X3172 VSS 209 210 ICV_42 $T=394590 321760 0 0 $X=393590 $Y=320760
X3173 VSS 211 212 ICV_42 $T=394590 325160 0 0 $X=393590 $Y=324160
X3174 VSS 213 214 ICV_42 $T=394590 328560 0 0 $X=393590 $Y=327560
X3175 VSS 215 216 ICV_42 $T=394590 331960 0 0 $X=393590 $Y=330960
X3176 VSS 217 218 ICV_42 $T=394590 335360 0 0 $X=393590 $Y=334360
X3177 VSS 219 220 ICV_42 $T=394590 338760 0 0 $X=393590 $Y=337760
X3178 VSS 221 222 ICV_42 $T=394590 342160 0 0 $X=393590 $Y=341160
X3179 VSS 223 224 ICV_42 $T=394590 345560 0 0 $X=393590 $Y=344560
X3180 VSS 225 226 ICV_42 $T=394590 348960 0 0 $X=393590 $Y=347960
X3181 VSS 227 228 ICV_42 $T=394590 352360 0 0 $X=393590 $Y=351360
X3182 VSS 229 230 ICV_42 $T=394590 355760 0 0 $X=393590 $Y=354760
X3183 VSS 231 232 ICV_42 $T=394590 359160 0 0 $X=393590 $Y=358160
X3184 VSS 233 234 ICV_42 $T=394590 362560 0 0 $X=393590 $Y=361560
X3185 VSS 235 236 ICV_42 $T=394590 365960 0 0 $X=393590 $Y=364960
X3186 VSS 237 238 ICV_42 $T=394590 369360 0 0 $X=393590 $Y=368360
X3187 VSS 239 240 ICV_42 $T=394590 372760 0 0 $X=393590 $Y=371760
X3188 VSS 241 242 ICV_42 $T=394590 376160 0 0 $X=393590 $Y=375160
X3189 VSS 243 244 ICV_42 $T=394590 379560 0 0 $X=393590 $Y=378560
X3190 VSS 245 246 ICV_42 $T=394590 382960 0 0 $X=393590 $Y=381960
X3191 VSS 247 248 ICV_42 $T=394590 386360 0 0 $X=393590 $Y=385360
X3192 VSS 249 250 ICV_42 $T=394590 389760 0 0 $X=393590 $Y=388760
X3193 VSS 251 252 ICV_42 $T=394590 393160 0 0 $X=393590 $Y=392160
X3194 VSS 253 254 ICV_42 $T=394590 396560 0 0 $X=393590 $Y=395560
X3195 VSS 255 256 ICV_42 $T=394590 399960 0 0 $X=393590 $Y=398960
X3196 VSS 257 258 ICV_42 $T=394590 403360 0 0 $X=393590 $Y=402360
X3197 VSS 259 260 ICV_42 $T=394590 406760 0 0 $X=393590 $Y=405760
X3198 VSS 261 262 ICV_42 $T=394590 410160 0 0 $X=393590 $Y=409160
X3199 VSS 263 264 ICV_42 $T=394590 413560 0 0 $X=393590 $Y=412560
X3200 VSS 265 266 ICV_42 $T=394590 416960 0 0 $X=393590 $Y=415960
X3201 VSS 267 268 ICV_42 $T=394590 420360 0 0 $X=393590 $Y=419360
X3202 VSS 269 270 ICV_42 $T=394590 423760 0 0 $X=393590 $Y=422760
X3203 VSS 271 272 ICV_42 $T=394590 427160 0 0 $X=393590 $Y=426160
X3204 VSS 273 274 ICV_42 $T=394590 430560 0 0 $X=393590 $Y=429560
X3205 VSS 275 276 ICV_42 $T=394590 433960 0 0 $X=393590 $Y=432960
X3206 VSS 277 278 ICV_42 $T=394590 437360 0 0 $X=393590 $Y=436360
X3207 VSS 279 280 ICV_42 $T=394590 440760 0 0 $X=393590 $Y=439760
X3208 VSS 281 282 ICV_42 $T=394590 444160 0 0 $X=393590 $Y=443160
X3209 VSS 283 284 ICV_42 $T=394590 447560 0 0 $X=393590 $Y=446560
X3210 VSS 285 286 ICV_42 $T=394590 450960 0 0 $X=393590 $Y=449960
X3211 VSS 287 288 ICV_42 $T=394590 454360 0 0 $X=393590 $Y=453360
X3212 VSS 289 290 ICV_42 $T=394590 457760 0 0 $X=393590 $Y=456760
X3213 VSS 291 292 ICV_42 $T=394590 461160 0 0 $X=393590 $Y=460160
X3214 VSS 293 294 ICV_42 $T=394590 464560 0 0 $X=393590 $Y=463560
X3215 VSS 295 296 ICV_42 $T=394590 467960 0 0 $X=393590 $Y=466960
X3216 VSS 297 298 ICV_42 $T=394590 471360 0 0 $X=393590 $Y=470360
X3217 VSS 299 300 ICV_42 $T=394590 474760 0 0 $X=393590 $Y=473760
X3218 VSS 301 302 ICV_42 $T=394590 478160 0 0 $X=393590 $Y=477160
X3219 VSS 303 304 ICV_42 $T=394590 481560 0 0 $X=393590 $Y=480560
X3220 VSS 305 306 ICV_42 $T=394590 484960 0 0 $X=393590 $Y=483960
X3221 VSS 307 308 ICV_42 $T=394590 488360 0 0 $X=393590 $Y=487360
X3222 VSS 309 310 ICV_42 $T=394590 491760 0 0 $X=393590 $Y=490760
X3223 VSS 311 312 ICV_42 $T=394590 495160 0 0 $X=393590 $Y=494160
X3224 VSS 313 314 ICV_42 $T=394590 498560 0 0 $X=393590 $Y=497560
X3225 VSS 315 316 ICV_42 $T=394590 501960 0 0 $X=393590 $Y=500960
X3226 VSS 317 318 ICV_42 $T=394590 505360 0 0 $X=393590 $Y=504360
X3492 VDD VSS 3329 3330 A8FCELLE_D_LP $T=88010 509800 0 0 $X=87790 $Y=509330
X3493 VDD VSS 3331 3332 A8FCELLE_D_LP $T=89210 513200 0 180 $X=87790 $Y=511170
X3494 VSS VDD 3333 3334 SIGN_MEMCCEG $T=12410 509800 0 0 $X=11410 $Y=508800
X3495 VSS VDD 3335 3336 SIGN_MEMCCEG $T=13610 513200 0 180 $X=11410 $Y=510500
X3496 VSS VDD 3337 3338 SIGN_MEMCCEG $T=17210 509800 0 0 $X=16210 $Y=508800
X3497 VSS VDD 3339 3340 SIGN_MEMCCEG $T=18410 513200 0 180 $X=16210 $Y=510500
X3498 VSS VDD 3341 3342 SIGN_MEMCCEG $T=22010 509800 0 0 $X=21010 $Y=508800
X3499 VSS VDD 3343 3344 SIGN_MEMCCEG $T=23210 513200 0 180 $X=21010 $Y=510500
X3500 VSS VDD 3345 3346 SIGN_MEMCCEG $T=26810 509800 0 0 $X=25810 $Y=508800
X3501 VSS VDD 3347 3348 SIGN_MEMCCEG $T=28010 513200 0 180 $X=25810 $Y=510500
X3502 VSS VDD 3349 3350 SIGN_MEMCCEG $T=31610 509800 0 0 $X=30610 $Y=508800
X3503 VSS VDD 3351 3352 SIGN_MEMCCEG $T=32810 513200 0 180 $X=30610 $Y=510500
X3504 VSS VDD 3353 3354 SIGN_MEMCCEG $T=36410 509800 0 0 $X=35410 $Y=508800
X3505 VSS VDD 3355 3356 SIGN_MEMCCEG $T=37610 513200 0 180 $X=35410 $Y=510500
X3506 VSS VDD 3357 3358 SIGN_MEMCCEG $T=41210 509800 0 0 $X=40210 $Y=508800
X3507 VSS VDD 3359 3360 SIGN_MEMCCEG $T=42410 513200 0 180 $X=40210 $Y=510500
X3508 VSS VDD 3361 3362 SIGN_MEMCCEG $T=46010 509800 0 0 $X=45010 $Y=508800
X3509 VSS VDD 3363 3364 SIGN_MEMCCEG $T=47210 513200 0 180 $X=45010 $Y=510500
X3510 VSS VDD 3365 3366 SIGN_MEMCCEG $T=52010 509800 0 0 $X=51010 $Y=508800
X3511 VSS VDD 3367 3368 SIGN_MEMCCEG $T=53210 513200 0 180 $X=51010 $Y=510500
X3512 VSS VDD 3369 3370 SIGN_MEMCCEG $T=56810 509800 0 0 $X=55810 $Y=508800
X3513 VSS VDD 3371 3372 SIGN_MEMCCEG $T=58010 513200 0 180 $X=55810 $Y=510500
X3514 VSS VDD 3373 3374 SIGN_MEMCCEG $T=61610 509800 0 0 $X=60610 $Y=508800
X3515 VSS VDD 3375 3376 SIGN_MEMCCEG $T=62810 513200 0 180 $X=60610 $Y=510500
X3516 VSS VDD 3377 3378 SIGN_MEMCCEG $T=66410 509800 0 0 $X=65410 $Y=508800
X3517 VSS VDD 3379 3380 SIGN_MEMCCEG $T=67610 513200 0 180 $X=65410 $Y=510500
X3518 VSS VDD 3381 3382 SIGN_MEMCCEG $T=71210 509800 0 0 $X=70210 $Y=508800
X3519 VSS VDD 3383 3384 SIGN_MEMCCEG $T=72410 513200 0 180 $X=70210 $Y=510500
X3520 VSS VDD 3385 3386 SIGN_MEMCCEG $T=76010 509800 0 0 $X=75010 $Y=508800
X3521 VSS VDD 3387 3388 SIGN_MEMCCEG $T=77210 513200 0 180 $X=75010 $Y=510500
X3522 VSS VDD 3389 3390 SIGN_MEMCCEG $T=80810 509800 0 0 $X=79810 $Y=508800
X3523 VSS VDD 3391 3392 SIGN_MEMCCEG $T=82010 513200 0 180 $X=79810 $Y=510500
X3524 VSS VDD 3393 3394 SIGN_MEMCCEG $T=85610 509800 0 0 $X=84610 $Y=508800
X3525 VSS VDD 3395 3396 SIGN_MEMCCEG $T=86810 513200 0 180 $X=84610 $Y=510500
X3526 VSS VDD 3397 3398 SIGN_MEMCCEG $T=91610 509800 0 0 $X=90610 $Y=508800
X3527 VSS VDD 3399 3400 SIGN_MEMCCEG $T=92810 513200 0 180 $X=90610 $Y=510500
X3528 VSS VDD 3401 3402 SIGN_MEMCCEG $T=96410 509800 0 0 $X=95410 $Y=508800
X3529 VSS VDD 3403 3404 SIGN_MEMCCEG $T=97610 513200 0 180 $X=95410 $Y=510500
X3530 VSS VDD 3405 3406 SIGN_MEMCCEG $T=101210 509800 0 0 $X=100210 $Y=508800
X3531 VSS VDD 3407 3408 SIGN_MEMCCEG $T=102410 513200 0 180 $X=100210 $Y=510500
X3532 VSS VDD 3409 3410 SIGN_MEMCCEG $T=106010 509800 0 0 $X=105010 $Y=508800
X3533 VSS VDD 3411 3412 SIGN_MEMCCEG $T=107210 513200 0 180 $X=105010 $Y=510500
X3534 VSS VDD 3413 3414 SIGN_MEMCCEG $T=110810 509800 0 0 $X=109810 $Y=508800
X3535 VSS VDD 3415 3416 SIGN_MEMCCEG $T=112010 513200 0 180 $X=109810 $Y=510500
X3536 VSS VDD 3417 3418 SIGN_MEMCCEG $T=115610 509800 0 0 $X=114610 $Y=508800
X3537 VSS VDD 3419 3420 SIGN_MEMCCEG $T=116810 513200 0 180 $X=114610 $Y=510500
X3538 VSS VDD 3421 3422 SIGN_MEMCCEG $T=120410 509800 0 0 $X=119410 $Y=508800
X3539 VSS VDD 3423 3424 SIGN_MEMCCEG $T=121610 513200 0 180 $X=119410 $Y=510500
X3540 VSS VDD 3425 3426 SIGN_MEMCCEG $T=125210 509800 0 0 $X=124210 $Y=508800
X3541 VSS VDD 3427 3428 SIGN_MEMCCEG $T=126410 513200 0 180 $X=124210 $Y=510500
X3542 VSS VDD 3429 3430 SIGN_MEMCCEG $T=131210 509800 0 0 $X=130210 $Y=508800
X3543 VSS VDD 3431 3432 SIGN_MEMCCEG $T=132410 513200 0 180 $X=130210 $Y=510500
X3544 VSS VDD 3433 3434 SIGN_MEMCCEG $T=136010 509800 0 0 $X=135010 $Y=508800
X3545 VSS VDD 3435 3436 SIGN_MEMCCEG $T=137210 513200 0 180 $X=135010 $Y=510500
X3546 VSS VDD 3437 3438 SIGN_MEMCCEG $T=140810 509800 0 0 $X=139810 $Y=508800
X3547 VSS VDD 3439 3440 SIGN_MEMCCEG $T=142010 513200 0 180 $X=139810 $Y=510500
X3548 VSS VDD 3441 3442 SIGN_MEMCCEG $T=145610 509800 0 0 $X=144610 $Y=508800
X3549 VSS VDD 3443 3444 SIGN_MEMCCEG $T=146810 513200 0 180 $X=144610 $Y=510500
X3550 VSS VDD 3445 3446 SIGN_MEMCCEG $T=150410 509800 0 0 $X=149410 $Y=508800
X3551 VSS VDD 3447 3448 SIGN_MEMCCEG $T=151610 513200 0 180 $X=149410 $Y=510500
X3552 VSS VDD 3449 3450 SIGN_MEMCCEG $T=155210 509800 0 0 $X=154210 $Y=508800
X3553 VSS VDD 3451 3452 SIGN_MEMCCEG $T=156410 513200 0 180 $X=154210 $Y=510500
X3554 VSS VDD 3453 3454 SIGN_MEMCCEG $T=160010 509800 0 0 $X=159010 $Y=508800
X3555 VSS VDD 3455 3456 SIGN_MEMCCEG $T=161210 513200 0 180 $X=159010 $Y=510500
X3556 VSS VDD 3457 3458 SIGN_MEMCCEG $T=164810 509800 0 0 $X=163810 $Y=508800
X3557 VSS VDD 3459 3460 SIGN_MEMCCEG $T=166010 513200 0 180 $X=163810 $Y=510500
X3558 VSS VDD 3461 3462 SIGN_MEMCCEG $T=237390 509800 0 0 $X=236390 $Y=508800
X3559 VSS VDD 3463 3464 SIGN_MEMCCEG $T=238590 513200 0 180 $X=236390 $Y=510500
X3560 VSS VDD 3465 3466 SIGN_MEMCCEG $T=242190 509800 0 0 $X=241190 $Y=508800
X3561 VSS VDD 3467 3468 SIGN_MEMCCEG $T=243390 513200 0 180 $X=241190 $Y=510500
X3562 VSS VDD 3469 3470 SIGN_MEMCCEG $T=246990 509800 0 0 $X=245990 $Y=508800
X3563 VSS VDD 3471 3472 SIGN_MEMCCEG $T=248190 513200 0 180 $X=245990 $Y=510500
X3564 VSS VDD 3473 3474 SIGN_MEMCCEG $T=251790 509800 0 0 $X=250790 $Y=508800
X3565 VSS VDD 3475 3476 SIGN_MEMCCEG $T=252990 513200 0 180 $X=250790 $Y=510500
X3566 VSS VDD 3477 3478 SIGN_MEMCCEG $T=256590 509800 0 0 $X=255590 $Y=508800
X3567 VSS VDD 3479 3480 SIGN_MEMCCEG $T=257790 513200 0 180 $X=255590 $Y=510500
X3568 VSS VDD 3481 3482 SIGN_MEMCCEG $T=261390 509800 0 0 $X=260390 $Y=508800
X3569 VSS VDD 3483 3484 SIGN_MEMCCEG $T=262590 513200 0 180 $X=260390 $Y=510500
X3570 VSS VDD 3485 3486 SIGN_MEMCCEG $T=266190 509800 0 0 $X=265190 $Y=508800
X3571 VSS VDD 3487 3488 SIGN_MEMCCEG $T=267390 513200 0 180 $X=265190 $Y=510500
X3572 VSS VDD 3489 3490 SIGN_MEMCCEG $T=270990 509800 0 0 $X=269990 $Y=508800
X3573 VSS VDD 3491 3492 SIGN_MEMCCEG $T=272190 513200 0 180 $X=269990 $Y=510500
X3574 VSS VDD 3493 3494 SIGN_MEMCCEG $T=276990 509800 0 0 $X=275990 $Y=508800
X3575 VSS VDD 3495 3496 SIGN_MEMCCEG $T=278190 513200 0 180 $X=275990 $Y=510500
X3576 VSS VDD 3497 3498 SIGN_MEMCCEG $T=281790 509800 0 0 $X=280790 $Y=508800
X3577 VSS VDD 3499 3500 SIGN_MEMCCEG $T=282990 513200 0 180 $X=280790 $Y=510500
X3578 VSS VDD 3501 3502 SIGN_MEMCCEG $T=286590 509800 0 0 $X=285590 $Y=508800
X3579 VSS VDD 3503 3504 SIGN_MEMCCEG $T=287790 513200 0 180 $X=285590 $Y=510500
X3580 VSS VDD 3505 3506 SIGN_MEMCCEG $T=291390 509800 0 0 $X=290390 $Y=508800
X3581 VSS VDD 3507 3508 SIGN_MEMCCEG $T=292590 513200 0 180 $X=290390 $Y=510500
X3582 VSS VDD 3509 3510 SIGN_MEMCCEG $T=296190 509800 0 0 $X=295190 $Y=508800
X3583 VSS VDD 3511 3512 SIGN_MEMCCEG $T=297390 513200 0 180 $X=295190 $Y=510500
X3584 VSS VDD 3513 3514 SIGN_MEMCCEG $T=300990 509800 0 0 $X=299990 $Y=508800
X3585 VSS VDD 3515 3516 SIGN_MEMCCEG $T=302190 513200 0 180 $X=299990 $Y=510500
X3586 VSS VDD 3517 3518 SIGN_MEMCCEG $T=305790 509800 0 0 $X=304790 $Y=508800
X3587 VSS VDD 3519 3520 SIGN_MEMCCEG $T=306990 513200 0 180 $X=304790 $Y=510500
X3588 VSS VDD 3521 3522 SIGN_MEMCCEG $T=310590 509800 0 0 $X=309590 $Y=508800
X3589 VSS VDD 3523 3524 SIGN_MEMCCEG $T=311790 513200 0 180 $X=309590 $Y=510500
X3590 VSS VDD 3525 3526 SIGN_MEMCCEG $T=321390 509800 0 0 $X=320390 $Y=508800
X3591 VSS VDD 3527 3528 SIGN_MEMCCEG $T=322590 513200 0 180 $X=320390 $Y=510500
X3592 VSS VDD 3529 3530 SIGN_MEMCCEG $T=326190 509800 0 0 $X=325190 $Y=508800
X3593 VSS VDD 3531 3532 SIGN_MEMCCEG $T=327390 513200 0 180 $X=325190 $Y=510500
X3594 VSS VDD 3533 3534 SIGN_MEMCCEG $T=330990 509800 0 0 $X=329990 $Y=508800
X3595 VSS VDD 3535 3536 SIGN_MEMCCEG $T=332190 513200 0 180 $X=329990 $Y=510500
X3596 VSS VDD 3537 3538 SIGN_MEMCCEG $T=335790 509800 0 0 $X=334790 $Y=508800
X3597 VSS VDD 3539 3540 SIGN_MEMCCEG $T=336990 513200 0 180 $X=334790 $Y=510500
X3598 VSS VDD 3541 3542 SIGN_MEMCCEG $T=340590 509800 0 0 $X=339590 $Y=508800
X3599 VSS VDD 3543 3544 SIGN_MEMCCEG $T=341790 513200 0 180 $X=339590 $Y=510500
X3600 VSS VDD 3545 3546 SIGN_MEMCCEG $T=345390 509800 0 0 $X=344390 $Y=508800
X3601 VSS VDD 3547 3548 SIGN_MEMCCEG $T=346590 513200 0 180 $X=344390 $Y=510500
X3602 VSS VDD 3549 3550 SIGN_MEMCCEG $T=350190 509800 0 0 $X=349190 $Y=508800
X3603 VSS VDD 3551 3552 SIGN_MEMCCEG $T=351390 513200 0 180 $X=349190 $Y=510500
X3604 VSS VDD 3553 3554 SIGN_MEMCCEG $T=356190 509800 0 0 $X=355190 $Y=508800
X3605 VSS VDD 3555 3556 SIGN_MEMCCEG $T=357390 513200 0 180 $X=355190 $Y=510500
X3606 VSS VDD 3557 3558 SIGN_MEMCCEG $T=360990 509800 0 0 $X=359990 $Y=508800
X3607 VSS VDD 3559 3560 SIGN_MEMCCEG $T=362190 513200 0 180 $X=359990 $Y=510500
X3608 VSS VDD 3561 3562 SIGN_MEMCCEG $T=365790 509800 0 0 $X=364790 $Y=508800
X3609 VSS VDD 3563 3564 SIGN_MEMCCEG $T=366990 513200 0 180 $X=364790 $Y=510500
X3610 VSS VDD 3565 3566 SIGN_MEMCCEG $T=370590 509800 0 0 $X=369590 $Y=508800
X3611 VSS VDD 3567 3568 SIGN_MEMCCEG $T=371790 513200 0 180 $X=369590 $Y=510500
X3612 VSS VDD 3569 3570 SIGN_MEMCCEG $T=375390 509800 0 0 $X=374390 $Y=508800
X3613 VSS VDD 3571 3572 SIGN_MEMCCEG $T=376590 513200 0 180 $X=374390 $Y=510500
X3614 VSS VDD 3573 3574 SIGN_MEMCCEG $T=380190 509800 0 0 $X=379190 $Y=508800
X3615 VSS VDD 3575 3576 SIGN_MEMCCEG $T=381390 513200 0 180 $X=379190 $Y=510500
X3616 VSS VDD 3577 3578 SIGN_MEMCCEG $T=384990 509800 0 0 $X=383990 $Y=508800
X3617 VSS VDD 3579 3580 SIGN_MEMCCEG $T=386190 513200 0 180 $X=383990 $Y=510500
X3618 VSS VDD 3581 3582 SIGN_MEMCCEG $T=389790 509800 0 0 $X=388790 $Y=508800
X3619 VSS VDD 3583 3584 SIGN_MEMCCEG $T=390990 513200 0 180 $X=388790 $Y=510500
X3620 VSS VDD 3585 3586 A8FCELLO_D_LP $T=318990 509800 1 180 $X=317570 $Y=509330
X3621 VSS VDD 3587 3588 A8FCELLO_D_LP $T=317790 513200 1 0 $X=317570 $Y=511170
X3622 VDD VSS 3589 3590 SIGN_MEMCCOP $T=14810 509800 1 180 $X=12610 $Y=508800
X3623 VDD VSS 3591 3592 SIGN_MEMCCOP $T=13610 513200 1 0 $X=12610 $Y=510500
X3624 VDD VSS 3593 3594 SIGN_MEMCCOP $T=19610 509800 1 180 $X=17410 $Y=508800
X3625 VDD VSS 3595 3596 SIGN_MEMCCOP $T=18410 513200 1 0 $X=17410 $Y=510500
X3626 VDD VSS 3597 3598 SIGN_MEMCCOP $T=24410 509800 1 180 $X=22210 $Y=508800
X3627 VDD VSS 3599 3600 SIGN_MEMCCOP $T=23210 513200 1 0 $X=22210 $Y=510500
X3628 VDD VSS 3601 3602 SIGN_MEMCCOP $T=29210 509800 1 180 $X=27010 $Y=508800
X3629 VDD VSS 3603 3604 SIGN_MEMCCOP $T=28010 513200 1 0 $X=27010 $Y=510500
X3630 VDD VSS 3605 3606 SIGN_MEMCCOP $T=34010 509800 1 180 $X=31810 $Y=508800
X3631 VDD VSS 3607 3608 SIGN_MEMCCOP $T=32810 513200 1 0 $X=31810 $Y=510500
X3632 VDD VSS 3609 3610 SIGN_MEMCCOP $T=38810 509800 1 180 $X=36610 $Y=508800
X3633 VDD VSS 3611 3612 SIGN_MEMCCOP $T=37610 513200 1 0 $X=36610 $Y=510500
X3634 VDD VSS 3613 3614 SIGN_MEMCCOP $T=43610 509800 1 180 $X=41410 $Y=508800
X3635 VDD VSS 3615 3616 SIGN_MEMCCOP $T=42410 513200 1 0 $X=41410 $Y=510500
X3636 VDD VSS 3617 3618 SIGN_MEMCCOP $T=48410 509800 1 180 $X=46210 $Y=508800
X3637 VDD VSS 3619 3620 SIGN_MEMCCOP $T=47210 513200 1 0 $X=46210 $Y=510500
X3638 VDD VSS 3621 3622 SIGN_MEMCCOP $T=54410 509800 1 180 $X=52210 $Y=508800
X3639 VDD VSS 3623 3624 SIGN_MEMCCOP $T=53210 513200 1 0 $X=52210 $Y=510500
X3640 VDD VSS 3625 3626 SIGN_MEMCCOP $T=59210 509800 1 180 $X=57010 $Y=508800
X3641 VDD VSS 3627 3628 SIGN_MEMCCOP $T=58010 513200 1 0 $X=57010 $Y=510500
X3642 VDD VSS 3629 3630 SIGN_MEMCCOP $T=64010 509800 1 180 $X=61810 $Y=508800
X3643 VDD VSS 3631 3632 SIGN_MEMCCOP $T=62810 513200 1 0 $X=61810 $Y=510500
X3644 VDD VSS 3633 3634 SIGN_MEMCCOP $T=68810 509800 1 180 $X=66610 $Y=508800
X3645 VDD VSS 3635 3636 SIGN_MEMCCOP $T=67610 513200 1 0 $X=66610 $Y=510500
X3646 VDD VSS 3637 3638 SIGN_MEMCCOP $T=73610 509800 1 180 $X=71410 $Y=508800
X3647 VDD VSS 3639 3640 SIGN_MEMCCOP $T=72410 513200 1 0 $X=71410 $Y=510500
X3648 VDD VSS 3641 3642 SIGN_MEMCCOP $T=78410 509800 1 180 $X=76210 $Y=508800
X3649 VDD VSS 3643 3644 SIGN_MEMCCOP $T=77210 513200 1 0 $X=76210 $Y=510500
X3650 VDD VSS 3645 3646 SIGN_MEMCCOP $T=83210 509800 1 180 $X=81010 $Y=508800
X3651 VDD VSS 3647 3648 SIGN_MEMCCOP $T=82010 513200 1 0 $X=81010 $Y=510500
X3652 VDD VSS 3649 3650 SIGN_MEMCCOP $T=88010 509800 1 180 $X=85810 $Y=508800
X3653 VDD VSS 3651 3652 SIGN_MEMCCOP $T=86810 513200 1 0 $X=85810 $Y=510500
X3654 VDD VSS 3653 3654 SIGN_MEMCCOP $T=94010 509800 1 180 $X=91810 $Y=508800
X3655 VDD VSS 3655 3656 SIGN_MEMCCOP $T=92810 513200 1 0 $X=91810 $Y=510500
X3656 VDD VSS 3657 3658 SIGN_MEMCCOP $T=98810 509800 1 180 $X=96610 $Y=508800
X3657 VDD VSS 3659 3660 SIGN_MEMCCOP $T=97610 513200 1 0 $X=96610 $Y=510500
X3658 VDD VSS 3661 3662 SIGN_MEMCCOP $T=103610 509800 1 180 $X=101410 $Y=508800
X3659 VDD VSS 3663 3664 SIGN_MEMCCOP $T=102410 513200 1 0 $X=101410 $Y=510500
X3660 VDD VSS 3665 3666 SIGN_MEMCCOP $T=108410 509800 1 180 $X=106210 $Y=508800
X3661 VDD VSS 3667 3668 SIGN_MEMCCOP $T=107210 513200 1 0 $X=106210 $Y=510500
X3662 VDD VSS 3669 3670 SIGN_MEMCCOP $T=113210 509800 1 180 $X=111010 $Y=508800
X3663 VDD VSS 3671 3672 SIGN_MEMCCOP $T=112010 513200 1 0 $X=111010 $Y=510500
X3664 VDD VSS 3673 3674 SIGN_MEMCCOP $T=118010 509800 1 180 $X=115810 $Y=508800
X3665 VDD VSS 3675 3676 SIGN_MEMCCOP $T=116810 513200 1 0 $X=115810 $Y=510500
X3666 VDD VSS 3677 3678 SIGN_MEMCCOP $T=122810 509800 1 180 $X=120610 $Y=508800
X3667 VDD VSS 3679 3680 SIGN_MEMCCOP $T=121610 513200 1 0 $X=120610 $Y=510500
X3668 VDD VSS 3681 3682 SIGN_MEMCCOP $T=127610 509800 1 180 $X=125410 $Y=508800
X3669 VDD VSS 3683 3684 SIGN_MEMCCOP $T=126410 513200 1 0 $X=125410 $Y=510500
X3670 VDD VSS 3685 3686 SIGN_MEMCCOP $T=133610 509800 1 180 $X=131410 $Y=508800
X3671 VDD VSS 3687 3688 SIGN_MEMCCOP $T=132410 513200 1 0 $X=131410 $Y=510500
X3672 VDD VSS 3689 3690 SIGN_MEMCCOP $T=138410 509800 1 180 $X=136210 $Y=508800
X3673 VDD VSS 3691 3692 SIGN_MEMCCOP $T=137210 513200 1 0 $X=136210 $Y=510500
X3674 VDD VSS 3693 3694 SIGN_MEMCCOP $T=143210 509800 1 180 $X=141010 $Y=508800
X3675 VDD VSS 3695 3696 SIGN_MEMCCOP $T=142010 513200 1 0 $X=141010 $Y=510500
X3676 VDD VSS 3697 3698 SIGN_MEMCCOP $T=148010 509800 1 180 $X=145810 $Y=508800
X3677 VDD VSS 3699 3700 SIGN_MEMCCOP $T=146810 513200 1 0 $X=145810 $Y=510500
X3678 VDD VSS 3701 3702 SIGN_MEMCCOP $T=152810 509800 1 180 $X=150610 $Y=508800
X3679 VDD VSS 3703 3704 SIGN_MEMCCOP $T=151610 513200 1 0 $X=150610 $Y=510500
X3680 VDD VSS 3705 3706 SIGN_MEMCCOP $T=157610 509800 1 180 $X=155410 $Y=508800
X3681 VDD VSS 3707 3708 SIGN_MEMCCOP $T=156410 513200 1 0 $X=155410 $Y=510500
X3682 VDD VSS 3709 3710 SIGN_MEMCCOP $T=162410 509800 1 180 $X=160210 $Y=508800
X3683 VDD VSS 3711 3712 SIGN_MEMCCOP $T=161210 513200 1 0 $X=160210 $Y=510500
X3684 VDD VSS 3713 3714 SIGN_MEMCCOP $T=167210 509800 1 180 $X=165010 $Y=508800
X3685 VDD VSS 3715 3716 SIGN_MEMCCOP $T=166010 513200 1 0 $X=165010 $Y=510500
X3686 VDD VSS 3717 3718 SIGN_MEMCCOP $T=236190 73560 1 180 $X=233990 $Y=72560
X3687 VDD VSS 3719 3720 SIGN_MEMCCOP $T=234990 76960 1 0 $X=233990 $Y=74260
X3688 VDD VSS 3721 3722 SIGN_MEMCCOP $T=234990 76960 0 0 $X=233990 $Y=75960
X3689 VDD VSS 3723 3724 SIGN_MEMCCOP $T=236190 80360 0 180 $X=233990 $Y=77660
X3690 VDD VSS 3725 3726 SIGN_MEMCCOP $T=236190 80360 1 180 $X=233990 $Y=79360
X3691 VDD VSS 3727 3728 SIGN_MEMCCOP $T=234990 83760 1 0 $X=233990 $Y=81060
X3692 VDD VSS 3729 3730 SIGN_MEMCCOP $T=234990 83760 0 0 $X=233990 $Y=82760
X3693 VDD VSS 3731 3732 SIGN_MEMCCOP $T=236190 87160 0 180 $X=233990 $Y=84460
X3694 VDD VSS 3733 3734 SIGN_MEMCCOP $T=236190 87160 1 180 $X=233990 $Y=86160
X3695 VDD VSS 3735 3736 SIGN_MEMCCOP $T=234990 90560 1 0 $X=233990 $Y=87860
X3696 VDD VSS 3737 3738 SIGN_MEMCCOP $T=234990 90560 0 0 $X=233990 $Y=89560
X3697 VDD VSS 3739 3740 SIGN_MEMCCOP $T=236190 93960 0 180 $X=233990 $Y=91260
X3698 VDD VSS 3741 3742 SIGN_MEMCCOP $T=236190 93960 1 180 $X=233990 $Y=92960
X3699 VDD VSS 3743 3744 SIGN_MEMCCOP $T=234990 97360 1 0 $X=233990 $Y=94660
X3700 VDD VSS 3745 3746 SIGN_MEMCCOP $T=234990 97360 0 0 $X=233990 $Y=96360
X3701 VDD VSS 3747 3748 SIGN_MEMCCOP $T=236190 100760 0 180 $X=233990 $Y=98060
X3702 VDD VSS 3749 3750 SIGN_MEMCCOP $T=236190 100760 1 180 $X=233990 $Y=99760
X3703 VDD VSS 3751 3752 SIGN_MEMCCOP $T=234990 104160 1 0 $X=233990 $Y=101460
X3704 VDD VSS 3753 3754 SIGN_MEMCCOP $T=234990 104160 0 0 $X=233990 $Y=103160
X3705 VDD VSS 3755 3756 SIGN_MEMCCOP $T=236190 107560 0 180 $X=233990 $Y=104860
X3706 VDD VSS 3757 3758 SIGN_MEMCCOP $T=236190 107560 1 180 $X=233990 $Y=106560
X3707 VDD VSS 3759 3760 SIGN_MEMCCOP $T=234990 110960 1 0 $X=233990 $Y=108260
X3708 VDD VSS 3761 3762 SIGN_MEMCCOP $T=234990 110960 0 0 $X=233990 $Y=109960
X3709 VDD VSS 3763 3764 SIGN_MEMCCOP $T=236190 114360 0 180 $X=233990 $Y=111660
X3710 VDD VSS 3765 3766 SIGN_MEMCCOP $T=236190 114360 1 180 $X=233990 $Y=113360
X3711 VDD VSS 3767 3768 SIGN_MEMCCOP $T=234990 117760 1 0 $X=233990 $Y=115060
X3712 VDD VSS 3769 3770 SIGN_MEMCCOP $T=234990 117760 0 0 $X=233990 $Y=116760
X3713 VDD VSS 3771 3772 SIGN_MEMCCOP $T=236190 121160 0 180 $X=233990 $Y=118460
X3714 VDD VSS 3773 3774 SIGN_MEMCCOP $T=236190 121160 1 180 $X=233990 $Y=120160
X3715 VDD VSS 3775 3776 SIGN_MEMCCOP $T=234990 124560 1 0 $X=233990 $Y=121860
X3716 VDD VSS 3777 3778 SIGN_MEMCCOP $T=234990 124560 0 0 $X=233990 $Y=123560
X3717 VDD VSS 3779 3780 SIGN_MEMCCOP $T=236190 127960 0 180 $X=233990 $Y=125260
X3718 VDD VSS 3781 3782 SIGN_MEMCCOP $T=236190 127960 1 180 $X=233990 $Y=126960
X3719 VDD VSS 3783 3784 SIGN_MEMCCOP $T=234990 131360 1 0 $X=233990 $Y=128660
X3720 VDD VSS 3785 3786 SIGN_MEMCCOP $T=234990 131360 0 0 $X=233990 $Y=130360
X3721 VDD VSS 3787 3788 SIGN_MEMCCOP $T=236190 134760 0 180 $X=233990 $Y=132060
X3722 VDD VSS 3789 3790 SIGN_MEMCCOP $T=236190 134760 1 180 $X=233990 $Y=133760
X3723 VDD VSS 3791 3792 SIGN_MEMCCOP $T=234990 138160 1 0 $X=233990 $Y=135460
X3724 VDD VSS 3793 3794 SIGN_MEMCCOP $T=234990 138160 0 0 $X=233990 $Y=137160
X3725 VDD VSS 3795 3796 SIGN_MEMCCOP $T=236190 141560 0 180 $X=233990 $Y=138860
X3726 VDD VSS 3797 3798 SIGN_MEMCCOP $T=236190 141560 1 180 $X=233990 $Y=140560
X3727 VDD VSS 3799 3800 SIGN_MEMCCOP $T=234990 144960 1 0 $X=233990 $Y=142260
X3728 VDD VSS 3801 3802 SIGN_MEMCCOP $T=234990 144960 0 0 $X=233990 $Y=143960
X3729 VDD VSS 3803 3804 SIGN_MEMCCOP $T=236190 148360 0 180 $X=233990 $Y=145660
X3730 VDD VSS 3805 3806 SIGN_MEMCCOP $T=236190 148360 1 180 $X=233990 $Y=147360
X3731 VDD VSS 3807 3808 SIGN_MEMCCOP $T=234990 151760 1 0 $X=233990 $Y=149060
X3732 VDD VSS 3809 3810 SIGN_MEMCCOP $T=234990 151760 0 0 $X=233990 $Y=150760
X3733 VDD VSS 3811 3812 SIGN_MEMCCOP $T=236190 155160 0 180 $X=233990 $Y=152460
X3734 VDD VSS 3813 3814 SIGN_MEMCCOP $T=236190 155160 1 180 $X=233990 $Y=154160
X3735 VDD VSS 3815 3816 SIGN_MEMCCOP $T=234990 158560 1 0 $X=233990 $Y=155860
X3736 VDD VSS 3817 3818 SIGN_MEMCCOP $T=234990 158560 0 0 $X=233990 $Y=157560
X3737 VDD VSS 3819 3820 SIGN_MEMCCOP $T=236190 161960 0 180 $X=233990 $Y=159260
X3738 VDD VSS 3821 3822 SIGN_MEMCCOP $T=236190 161960 1 180 $X=233990 $Y=160960
X3739 VDD VSS 3823 3824 SIGN_MEMCCOP $T=234990 165360 1 0 $X=233990 $Y=162660
X3740 VDD VSS 3825 3826 SIGN_MEMCCOP $T=234990 165360 0 0 $X=233990 $Y=164360
X3741 VDD VSS 3827 3828 SIGN_MEMCCOP $T=236190 168760 0 180 $X=233990 $Y=166060
X3742 VDD VSS 3829 3830 SIGN_MEMCCOP $T=236190 168760 1 180 $X=233990 $Y=167760
X3743 VDD VSS 3831 3832 SIGN_MEMCCOP $T=234990 172160 1 0 $X=233990 $Y=169460
X3744 VDD VSS 3833 3834 SIGN_MEMCCOP $T=234990 172160 0 0 $X=233990 $Y=171160
X3745 VDD VSS 3835 3836 SIGN_MEMCCOP $T=236190 175560 0 180 $X=233990 $Y=172860
X3746 VDD VSS 3837 3838 SIGN_MEMCCOP $T=236190 175560 1 180 $X=233990 $Y=174560
X3747 VDD VSS 3839 3840 SIGN_MEMCCOP $T=234990 178960 1 0 $X=233990 $Y=176260
X3748 VDD VSS 3841 3842 SIGN_MEMCCOP $T=234990 178960 0 0 $X=233990 $Y=177960
X3749 VDD VSS 3843 3844 SIGN_MEMCCOP $T=236190 182360 0 180 $X=233990 $Y=179660
X3750 VDD VSS 3845 3846 SIGN_MEMCCOP $T=236190 182360 1 180 $X=233990 $Y=181360
X3751 VDD VSS 3847 3848 SIGN_MEMCCOP $T=234990 185760 1 0 $X=233990 $Y=183060
X3752 VDD VSS 3849 3850 SIGN_MEMCCOP $T=234990 185760 0 0 $X=233990 $Y=184760
X3753 VDD VSS 3851 3852 SIGN_MEMCCOP $T=236190 189160 0 180 $X=233990 $Y=186460
X3754 VDD VSS 3853 3854 SIGN_MEMCCOP $T=236190 189160 1 180 $X=233990 $Y=188160
X3755 VDD VSS 3855 3856 SIGN_MEMCCOP $T=234990 192560 1 0 $X=233990 $Y=189860
X3756 VDD VSS 3857 3858 SIGN_MEMCCOP $T=234990 192560 0 0 $X=233990 $Y=191560
X3757 VDD VSS 3859 3860 SIGN_MEMCCOP $T=236190 195960 0 180 $X=233990 $Y=193260
X3758 VDD VSS 3861 3862 SIGN_MEMCCOP $T=236190 195960 1 180 $X=233990 $Y=194960
X3759 VDD VSS 3863 3864 SIGN_MEMCCOP $T=234990 199360 1 0 $X=233990 $Y=196660
X3760 VDD VSS 3865 3866 SIGN_MEMCCOP $T=234990 199360 0 0 $X=233990 $Y=198360
X3761 VDD VSS 3867 3868 SIGN_MEMCCOP $T=236190 202760 0 180 $X=233990 $Y=200060
X3762 VDD VSS 3869 3870 SIGN_MEMCCOP $T=236190 202760 1 180 $X=233990 $Y=201760
X3763 VDD VSS 3871 3872 SIGN_MEMCCOP $T=234990 206160 1 0 $X=233990 $Y=203460
X3764 VDD VSS 3873 3874 SIGN_MEMCCOP $T=234990 206160 0 0 $X=233990 $Y=205160
X3765 VDD VSS 3875 3876 SIGN_MEMCCOP $T=236190 209560 0 180 $X=233990 $Y=206860
X3766 VDD VSS 3877 3878 SIGN_MEMCCOP $T=236190 209560 1 180 $X=233990 $Y=208560
X3767 VDD VSS 3879 3880 SIGN_MEMCCOP $T=234990 212960 1 0 $X=233990 $Y=210260
X3768 VDD VSS 3881 3882 SIGN_MEMCCOP $T=234990 212960 0 0 $X=233990 $Y=211960
X3769 VDD VSS 3883 3884 SIGN_MEMCCOP $T=236190 216360 0 180 $X=233990 $Y=213660
X3770 VDD VSS 3885 3886 SIGN_MEMCCOP $T=236190 216360 1 180 $X=233990 $Y=215360
X3771 VDD VSS 3887 3888 SIGN_MEMCCOP $T=234990 219760 1 0 $X=233990 $Y=217060
X3772 VDD VSS 3889 3890 SIGN_MEMCCOP $T=234990 219760 0 0 $X=233990 $Y=218760
X3773 VDD VSS 3891 3892 SIGN_MEMCCOP $T=236190 223160 0 180 $X=233990 $Y=220460
X3774 VDD VSS 3893 3894 SIGN_MEMCCOP $T=236190 223160 1 180 $X=233990 $Y=222160
X3775 VDD VSS 3895 3896 SIGN_MEMCCOP $T=234990 226560 1 0 $X=233990 $Y=223860
X3776 VDD VSS 3897 3898 SIGN_MEMCCOP $T=234990 226560 0 0 $X=233990 $Y=225560
X3777 VDD VSS 3899 3900 SIGN_MEMCCOP $T=236190 229960 0 180 $X=233990 $Y=227260
X3778 VDD VSS 3901 3902 SIGN_MEMCCOP $T=236190 229960 1 180 $X=233990 $Y=228960
X3779 VDD VSS 3903 3904 SIGN_MEMCCOP $T=234990 233360 1 0 $X=233990 $Y=230660
X3780 VDD VSS 3905 3906 SIGN_MEMCCOP $T=234990 233360 0 0 $X=233990 $Y=232360
X3781 VDD VSS 3907 3908 SIGN_MEMCCOP $T=236190 236760 0 180 $X=233990 $Y=234060
X3782 VDD VSS 3909 3910 SIGN_MEMCCOP $T=236190 236760 1 180 $X=233990 $Y=235760
X3783 VDD VSS 3911 3912 SIGN_MEMCCOP $T=234990 240160 1 0 $X=233990 $Y=237460
X3784 VDD VSS 3913 3914 SIGN_MEMCCOP $T=234990 240160 0 0 $X=233990 $Y=239160
X3785 VDD VSS 3915 3916 SIGN_MEMCCOP $T=236190 243560 0 180 $X=233990 $Y=240860
X3786 VDD VSS 3917 3918 SIGN_MEMCCOP $T=236190 243560 1 180 $X=233990 $Y=242560
X3787 VDD VSS 3919 3920 SIGN_MEMCCOP $T=234990 246960 1 0 $X=233990 $Y=244260
X3788 VDD VSS 3921 3922 SIGN_MEMCCOP $T=234990 246960 0 0 $X=233990 $Y=245960
X3789 VDD VSS 3923 3924 SIGN_MEMCCOP $T=236190 250360 0 180 $X=233990 $Y=247660
X3790 VDD VSS 3925 3926 SIGN_MEMCCOP $T=236190 250360 1 180 $X=233990 $Y=249360
X3791 VDD VSS 3927 3928 SIGN_MEMCCOP $T=234990 253760 1 0 $X=233990 $Y=251060
X3792 VDD VSS 3929 3930 SIGN_MEMCCOP $T=234990 253760 0 0 $X=233990 $Y=252760
X3793 VDD VSS 3931 3932 SIGN_MEMCCOP $T=236190 257160 0 180 $X=233990 $Y=254460
X3794 VDD VSS 3933 3934 SIGN_MEMCCOP $T=236190 257160 1 180 $X=233990 $Y=256160
X3795 VDD VSS 3935 3936 SIGN_MEMCCOP $T=234990 260560 1 0 $X=233990 $Y=257860
X3796 VDD VSS 3937 3938 SIGN_MEMCCOP $T=234990 260560 0 0 $X=233990 $Y=259560
X3797 VDD VSS 3939 3940 SIGN_MEMCCOP $T=236190 263960 0 180 $X=233990 $Y=261260
X3798 VDD VSS 3941 3942 SIGN_MEMCCOP $T=236190 263960 1 180 $X=233990 $Y=262960
X3799 VDD VSS 3943 3944 SIGN_MEMCCOP $T=234990 267360 1 0 $X=233990 $Y=264660
X3800 VDD VSS 3945 3946 SIGN_MEMCCOP $T=234990 267360 0 0 $X=233990 $Y=266360
X3801 VDD VSS 3947 3948 SIGN_MEMCCOP $T=236190 270760 0 180 $X=233990 $Y=268060
X3802 VDD VSS 3949 3950 SIGN_MEMCCOP $T=236190 270760 1 180 $X=233990 $Y=269760
X3803 VDD VSS 3951 3952 SIGN_MEMCCOP $T=234990 274160 1 0 $X=233990 $Y=271460
X3804 VDD VSS 3953 3954 SIGN_MEMCCOP $T=234990 274160 0 0 $X=233990 $Y=273160
X3805 VDD VSS 3955 3956 SIGN_MEMCCOP $T=236190 277560 0 180 $X=233990 $Y=274860
X3806 VDD VSS 3957 3958 SIGN_MEMCCOP $T=236190 277560 1 180 $X=233990 $Y=276560
X3807 VDD VSS 3959 3960 SIGN_MEMCCOP $T=234990 280960 1 0 $X=233990 $Y=278260
X3808 VDD VSS 3961 3962 SIGN_MEMCCOP $T=234990 280960 0 0 $X=233990 $Y=279960
X3809 VDD VSS 3963 3964 SIGN_MEMCCOP $T=236190 284360 0 180 $X=233990 $Y=281660
X3810 VDD VSS 3965 3966 SIGN_MEMCCOP $T=236190 284360 1 180 $X=233990 $Y=283360
X3811 VDD VSS 3967 3968 SIGN_MEMCCOP $T=234990 287760 1 0 $X=233990 $Y=285060
X3812 VDD VSS 3969 3970 SIGN_MEMCCOP $T=234990 287760 0 0 $X=233990 $Y=286760
X3813 VDD VSS 3971 3972 SIGN_MEMCCOP $T=236190 291160 0 180 $X=233990 $Y=288460
X3814 VDD VSS 3973 3974 SIGN_MEMCCOP $T=236190 291160 1 180 $X=233990 $Y=290160
X3815 VDD VSS 3975 3976 SIGN_MEMCCOP $T=234990 294560 1 0 $X=233990 $Y=291860
X3816 VDD VSS 3977 3978 SIGN_MEMCCOP $T=234990 294560 0 0 $X=233990 $Y=293560
X3817 VDD VSS 3979 3980 SIGN_MEMCCOP $T=236190 297960 0 180 $X=233990 $Y=295260
X3818 VDD VSS 3981 3982 SIGN_MEMCCOP $T=236190 297960 1 180 $X=233990 $Y=296960
X3819 VDD VSS 3983 3984 SIGN_MEMCCOP $T=234990 301360 1 0 $X=233990 $Y=298660
X3820 VDD VSS 3985 3986 SIGN_MEMCCOP $T=234990 301360 0 0 $X=233990 $Y=300360
X3821 VDD VSS 3987 3988 SIGN_MEMCCOP $T=236190 304760 0 180 $X=233990 $Y=302060
X3822 VDD VSS 3989 3990 SIGN_MEMCCOP $T=236190 304760 1 180 $X=233990 $Y=303760
X3823 VDD VSS 3991 3992 SIGN_MEMCCOP $T=234990 308160 1 0 $X=233990 $Y=305460
X3824 VDD VSS 3993 3994 SIGN_MEMCCOP $T=234990 308160 0 0 $X=233990 $Y=307160
X3825 VDD VSS 3995 3996 SIGN_MEMCCOP $T=236190 311560 0 180 $X=233990 $Y=308860
X3826 VDD VSS 3997 3998 SIGN_MEMCCOP $T=236190 311560 1 180 $X=233990 $Y=310560
X3827 VDD VSS 3999 4000 SIGN_MEMCCOP $T=234990 314960 1 0 $X=233990 $Y=312260
X3828 VDD VSS 4001 4002 SIGN_MEMCCOP $T=234990 314960 0 0 $X=233990 $Y=313960
X3829 VDD VSS 4003 4004 SIGN_MEMCCOP $T=236190 318360 0 180 $X=233990 $Y=315660
X3830 VDD VSS 4005 4006 SIGN_MEMCCOP $T=236190 318360 1 180 $X=233990 $Y=317360
X3831 VDD VSS 4007 4008 SIGN_MEMCCOP $T=234990 321760 1 0 $X=233990 $Y=319060
X3832 VDD VSS 4009 4010 SIGN_MEMCCOP $T=234990 321760 0 0 $X=233990 $Y=320760
X3833 VDD VSS 4011 4012 SIGN_MEMCCOP $T=236190 325160 0 180 $X=233990 $Y=322460
X3834 VDD VSS 4013 4014 SIGN_MEMCCOP $T=236190 325160 1 180 $X=233990 $Y=324160
X3835 VDD VSS 4015 4016 SIGN_MEMCCOP $T=234990 328560 1 0 $X=233990 $Y=325860
X3836 VDD VSS 4017 4018 SIGN_MEMCCOP $T=234990 328560 0 0 $X=233990 $Y=327560
X3837 VDD VSS 4019 4020 SIGN_MEMCCOP $T=236190 331960 0 180 $X=233990 $Y=329260
X3838 VDD VSS 4021 4022 SIGN_MEMCCOP $T=236190 331960 1 180 $X=233990 $Y=330960
X3839 VDD VSS 4023 4024 SIGN_MEMCCOP $T=234990 335360 1 0 $X=233990 $Y=332660
X3840 VDD VSS 4025 4026 SIGN_MEMCCOP $T=234990 335360 0 0 $X=233990 $Y=334360
X3841 VDD VSS 4027 4028 SIGN_MEMCCOP $T=236190 338760 0 180 $X=233990 $Y=336060
X3842 VDD VSS 4029 4030 SIGN_MEMCCOP $T=236190 338760 1 180 $X=233990 $Y=337760
X3843 VDD VSS 4031 4032 SIGN_MEMCCOP $T=234990 342160 1 0 $X=233990 $Y=339460
X3844 VDD VSS 4033 4034 SIGN_MEMCCOP $T=234990 342160 0 0 $X=233990 $Y=341160
X3845 VDD VSS 4035 4036 SIGN_MEMCCOP $T=236190 345560 0 180 $X=233990 $Y=342860
X3846 VDD VSS 4037 4038 SIGN_MEMCCOP $T=236190 345560 1 180 $X=233990 $Y=344560
X3847 VDD VSS 4039 4040 SIGN_MEMCCOP $T=234990 348960 1 0 $X=233990 $Y=346260
X3848 VDD VSS 4041 4042 SIGN_MEMCCOP $T=234990 348960 0 0 $X=233990 $Y=347960
X3849 VDD VSS 4043 4044 SIGN_MEMCCOP $T=236190 352360 0 180 $X=233990 $Y=349660
X3850 VDD VSS 4045 4046 SIGN_MEMCCOP $T=236190 352360 1 180 $X=233990 $Y=351360
X3851 VDD VSS 4047 4048 SIGN_MEMCCOP $T=234990 355760 1 0 $X=233990 $Y=353060
X3852 VDD VSS 4049 4050 SIGN_MEMCCOP $T=234990 355760 0 0 $X=233990 $Y=354760
X3853 VDD VSS 4051 4052 SIGN_MEMCCOP $T=236190 359160 0 180 $X=233990 $Y=356460
X3854 VDD VSS 4053 4054 SIGN_MEMCCOP $T=236190 359160 1 180 $X=233990 $Y=358160
X3855 VDD VSS 4055 4056 SIGN_MEMCCOP $T=234990 362560 1 0 $X=233990 $Y=359860
X3856 VDD VSS 4057 4058 SIGN_MEMCCOP $T=234990 362560 0 0 $X=233990 $Y=361560
X3857 VDD VSS 4059 4060 SIGN_MEMCCOP $T=236190 365960 0 180 $X=233990 $Y=363260
X3858 VDD VSS 4061 4062 SIGN_MEMCCOP $T=236190 365960 1 180 $X=233990 $Y=364960
X3859 VDD VSS 4063 4064 SIGN_MEMCCOP $T=234990 369360 1 0 $X=233990 $Y=366660
X3860 VDD VSS 4065 4066 SIGN_MEMCCOP $T=234990 369360 0 0 $X=233990 $Y=368360
X3861 VDD VSS 4067 4068 SIGN_MEMCCOP $T=236190 372760 0 180 $X=233990 $Y=370060
X3862 VDD VSS 4069 4070 SIGN_MEMCCOP $T=236190 372760 1 180 $X=233990 $Y=371760
X3863 VDD VSS 4071 4072 SIGN_MEMCCOP $T=234990 376160 1 0 $X=233990 $Y=373460
X3864 VDD VSS 4073 4074 SIGN_MEMCCOP $T=234990 376160 0 0 $X=233990 $Y=375160
X3865 VDD VSS 4075 4076 SIGN_MEMCCOP $T=236190 379560 0 180 $X=233990 $Y=376860
X3866 VDD VSS 4077 4078 SIGN_MEMCCOP $T=236190 379560 1 180 $X=233990 $Y=378560
X3867 VDD VSS 4079 4080 SIGN_MEMCCOP $T=234990 382960 1 0 $X=233990 $Y=380260
X3868 VDD VSS 4081 4082 SIGN_MEMCCOP $T=234990 382960 0 0 $X=233990 $Y=381960
X3869 VDD VSS 4083 4084 SIGN_MEMCCOP $T=236190 386360 0 180 $X=233990 $Y=383660
X3870 VDD VSS 4085 4086 SIGN_MEMCCOP $T=236190 386360 1 180 $X=233990 $Y=385360
X3871 VDD VSS 4087 4088 SIGN_MEMCCOP $T=234990 389760 1 0 $X=233990 $Y=387060
X3872 VDD VSS 4089 4090 SIGN_MEMCCOP $T=234990 389760 0 0 $X=233990 $Y=388760
X3873 VDD VSS 4091 4092 SIGN_MEMCCOP $T=236190 393160 0 180 $X=233990 $Y=390460
X3874 VDD VSS 4093 4094 SIGN_MEMCCOP $T=236190 393160 1 180 $X=233990 $Y=392160
X3875 VDD VSS 4095 4096 SIGN_MEMCCOP $T=234990 396560 1 0 $X=233990 $Y=393860
X3876 VDD VSS 4097 4098 SIGN_MEMCCOP $T=234990 396560 0 0 $X=233990 $Y=395560
X3877 VDD VSS 4099 4100 SIGN_MEMCCOP $T=236190 399960 0 180 $X=233990 $Y=397260
X3878 VDD VSS 4101 4102 SIGN_MEMCCOP $T=236190 399960 1 180 $X=233990 $Y=398960
X3879 VDD VSS 4103 4104 SIGN_MEMCCOP $T=234990 403360 1 0 $X=233990 $Y=400660
X3880 VDD VSS 4105 4106 SIGN_MEMCCOP $T=234990 403360 0 0 $X=233990 $Y=402360
X3881 VDD VSS 4107 4108 SIGN_MEMCCOP $T=236190 406760 0 180 $X=233990 $Y=404060
X3882 VDD VSS 4109 4110 SIGN_MEMCCOP $T=236190 406760 1 180 $X=233990 $Y=405760
X3883 VDD VSS 4111 4112 SIGN_MEMCCOP $T=234990 410160 1 0 $X=233990 $Y=407460
X3884 VDD VSS 4113 4114 SIGN_MEMCCOP $T=234990 410160 0 0 $X=233990 $Y=409160
X3885 VDD VSS 4115 4116 SIGN_MEMCCOP $T=236190 413560 0 180 $X=233990 $Y=410860
X3886 VDD VSS 4117 4118 SIGN_MEMCCOP $T=236190 413560 1 180 $X=233990 $Y=412560
X3887 VDD VSS 4119 4120 SIGN_MEMCCOP $T=234990 416960 1 0 $X=233990 $Y=414260
X3888 VDD VSS 4121 4122 SIGN_MEMCCOP $T=234990 416960 0 0 $X=233990 $Y=415960
X3889 VDD VSS 4123 4124 SIGN_MEMCCOP $T=236190 420360 0 180 $X=233990 $Y=417660
X3890 VDD VSS 4125 4126 SIGN_MEMCCOP $T=236190 420360 1 180 $X=233990 $Y=419360
X3891 VDD VSS 4127 4128 SIGN_MEMCCOP $T=234990 423760 1 0 $X=233990 $Y=421060
X3892 VDD VSS 4129 4130 SIGN_MEMCCOP $T=234990 423760 0 0 $X=233990 $Y=422760
X3893 VDD VSS 4131 4132 SIGN_MEMCCOP $T=236190 427160 0 180 $X=233990 $Y=424460
X3894 VDD VSS 4133 4134 SIGN_MEMCCOP $T=236190 427160 1 180 $X=233990 $Y=426160
X3895 VDD VSS 4135 4136 SIGN_MEMCCOP $T=234990 430560 1 0 $X=233990 $Y=427860
X3896 VDD VSS 4137 4138 SIGN_MEMCCOP $T=234990 430560 0 0 $X=233990 $Y=429560
X3897 VDD VSS 4139 4140 SIGN_MEMCCOP $T=236190 433960 0 180 $X=233990 $Y=431260
X3898 VDD VSS 4141 4142 SIGN_MEMCCOP $T=236190 433960 1 180 $X=233990 $Y=432960
X3899 VDD VSS 4143 4144 SIGN_MEMCCOP $T=234990 437360 1 0 $X=233990 $Y=434660
X3900 VDD VSS 4145 4146 SIGN_MEMCCOP $T=234990 437360 0 0 $X=233990 $Y=436360
X3901 VDD VSS 4147 4148 SIGN_MEMCCOP $T=236190 440760 0 180 $X=233990 $Y=438060
X3902 VDD VSS 4149 4150 SIGN_MEMCCOP $T=236190 440760 1 180 $X=233990 $Y=439760
X3903 VDD VSS 4151 4152 SIGN_MEMCCOP $T=234990 444160 1 0 $X=233990 $Y=441460
X3904 VDD VSS 4153 4154 SIGN_MEMCCOP $T=234990 444160 0 0 $X=233990 $Y=443160
X3905 VDD VSS 4155 4156 SIGN_MEMCCOP $T=236190 447560 0 180 $X=233990 $Y=444860
X3906 VDD VSS 4157 4158 SIGN_MEMCCOP $T=236190 447560 1 180 $X=233990 $Y=446560
X3907 VDD VSS 4159 4160 SIGN_MEMCCOP $T=234990 450960 1 0 $X=233990 $Y=448260
X3908 VDD VSS 4161 4162 SIGN_MEMCCOP $T=234990 450960 0 0 $X=233990 $Y=449960
X3909 VDD VSS 4163 4164 SIGN_MEMCCOP $T=236190 454360 0 180 $X=233990 $Y=451660
X3910 VDD VSS 4165 4166 SIGN_MEMCCOP $T=236190 454360 1 180 $X=233990 $Y=453360
X3911 VDD VSS 4167 4168 SIGN_MEMCCOP $T=234990 457760 1 0 $X=233990 $Y=455060
X3912 VDD VSS 4169 4170 SIGN_MEMCCOP $T=234990 457760 0 0 $X=233990 $Y=456760
X3913 VDD VSS 4171 4172 SIGN_MEMCCOP $T=236190 461160 0 180 $X=233990 $Y=458460
X3914 VDD VSS 4173 4174 SIGN_MEMCCOP $T=236190 461160 1 180 $X=233990 $Y=460160
X3915 VDD VSS 4175 4176 SIGN_MEMCCOP $T=234990 464560 1 0 $X=233990 $Y=461860
X3916 VDD VSS 4177 4178 SIGN_MEMCCOP $T=234990 464560 0 0 $X=233990 $Y=463560
X3917 VDD VSS 4179 4180 SIGN_MEMCCOP $T=236190 467960 0 180 $X=233990 $Y=465260
X3918 VDD VSS 4181 4182 SIGN_MEMCCOP $T=236190 467960 1 180 $X=233990 $Y=466960
X3919 VDD VSS 4183 4184 SIGN_MEMCCOP $T=234990 471360 1 0 $X=233990 $Y=468660
X3920 VDD VSS 4185 4186 SIGN_MEMCCOP $T=234990 471360 0 0 $X=233990 $Y=470360
X3921 VDD VSS 4187 4188 SIGN_MEMCCOP $T=236190 474760 0 180 $X=233990 $Y=472060
X3922 VDD VSS 4189 4190 SIGN_MEMCCOP $T=236190 474760 1 180 $X=233990 $Y=473760
X3923 VDD VSS 4191 4192 SIGN_MEMCCOP $T=234990 478160 1 0 $X=233990 $Y=475460
X3924 VDD VSS 4193 4194 SIGN_MEMCCOP $T=234990 478160 0 0 $X=233990 $Y=477160
X3925 VDD VSS 4195 4196 SIGN_MEMCCOP $T=236190 481560 0 180 $X=233990 $Y=478860
X3926 VDD VSS 4197 4198 SIGN_MEMCCOP $T=236190 481560 1 180 $X=233990 $Y=480560
X3927 VDD VSS 4199 4200 SIGN_MEMCCOP $T=234990 484960 1 0 $X=233990 $Y=482260
X3928 VDD VSS 4201 4202 SIGN_MEMCCOP $T=234990 484960 0 0 $X=233990 $Y=483960
X3929 VDD VSS 4203 4204 SIGN_MEMCCOP $T=236190 488360 0 180 $X=233990 $Y=485660
X3930 VDD VSS 4205 4206 SIGN_MEMCCOP $T=236190 488360 1 180 $X=233990 $Y=487360
X3931 VDD VSS 4207 4208 SIGN_MEMCCOP $T=234990 491760 1 0 $X=233990 $Y=489060
X3932 VDD VSS 4209 4210 SIGN_MEMCCOP $T=234990 491760 0 0 $X=233990 $Y=490760
X3933 VDD VSS 4211 4212 SIGN_MEMCCOP $T=236190 495160 0 180 $X=233990 $Y=492460
X3934 VDD VSS 4213 4214 SIGN_MEMCCOP $T=236190 495160 1 180 $X=233990 $Y=494160
X3935 VDD VSS 4215 4216 SIGN_MEMCCOP $T=234990 498560 1 0 $X=233990 $Y=495860
X3936 VDD VSS 4217 4218 SIGN_MEMCCOP $T=234990 498560 0 0 $X=233990 $Y=497560
X3937 VDD VSS 4219 4220 SIGN_MEMCCOP $T=236190 501960 0 180 $X=233990 $Y=499260
X3938 VDD VSS 4221 4222 SIGN_MEMCCOP $T=236190 501960 1 180 $X=233990 $Y=500960
X3939 VDD VSS 4223 4224 SIGN_MEMCCOP $T=234990 505360 1 0 $X=233990 $Y=502660
X3940 VDD VSS 4225 4226 SIGN_MEMCCOP $T=234990 505360 0 0 $X=233990 $Y=504360
X3941 VDD VSS 4227 4228 SIGN_MEMCCOP $T=236190 508760 0 180 $X=233990 $Y=506060
X3942 VDD VSS 4229 4230 SIGN_MEMCCOP $T=239790 509800 1 180 $X=237590 $Y=508800
X3943 VDD VSS 4231 4232 SIGN_MEMCCOP $T=238590 513200 1 0 $X=237590 $Y=510500
X3944 VDD VSS 4233 4234 SIGN_MEMCCOP $T=244590 509800 1 180 $X=242390 $Y=508800
X3945 VDD VSS 4235 4236 SIGN_MEMCCOP $T=243390 513200 1 0 $X=242390 $Y=510500
X3946 VDD VSS 4237 4238 SIGN_MEMCCOP $T=249390 509800 1 180 $X=247190 $Y=508800
X3947 VDD VSS 4239 4240 SIGN_MEMCCOP $T=248190 513200 1 0 $X=247190 $Y=510500
X3948 VDD VSS 4241 4242 SIGN_MEMCCOP $T=254190 509800 1 180 $X=251990 $Y=508800
X3949 VDD VSS 4243 4244 SIGN_MEMCCOP $T=252990 513200 1 0 $X=251990 $Y=510500
X3950 VDD VSS 4245 4246 SIGN_MEMCCOP $T=258990 509800 1 180 $X=256790 $Y=508800
X3951 VDD VSS 4247 4248 SIGN_MEMCCOP $T=257790 513200 1 0 $X=256790 $Y=510500
X3952 VDD VSS 4249 4250 SIGN_MEMCCOP $T=263790 509800 1 180 $X=261590 $Y=508800
X3953 VDD VSS 4251 4252 SIGN_MEMCCOP $T=262590 513200 1 0 $X=261590 $Y=510500
X3954 VDD VSS 4253 4254 SIGN_MEMCCOP $T=268590 509800 1 180 $X=266390 $Y=508800
X3955 VDD VSS 4255 4256 SIGN_MEMCCOP $T=267390 513200 1 0 $X=266390 $Y=510500
X3956 VDD VSS 4257 4258 SIGN_MEMCCOP $T=273390 509800 1 180 $X=271190 $Y=508800
X3957 VDD VSS 4259 4260 SIGN_MEMCCOP $T=272190 513200 1 0 $X=271190 $Y=510500
X3958 VDD VSS 4261 4262 SIGN_MEMCCOP $T=279390 509800 1 180 $X=277190 $Y=508800
X3959 VDD VSS 4263 4264 SIGN_MEMCCOP $T=278190 513200 1 0 $X=277190 $Y=510500
X3960 VDD VSS 4265 4266 SIGN_MEMCCOP $T=284190 509800 1 180 $X=281990 $Y=508800
X3961 VDD VSS 4267 4268 SIGN_MEMCCOP $T=282990 513200 1 0 $X=281990 $Y=510500
X3962 VDD VSS 4269 4270 SIGN_MEMCCOP $T=288990 509800 1 180 $X=286790 $Y=508800
X3963 VDD VSS 4271 4272 SIGN_MEMCCOP $T=287790 513200 1 0 $X=286790 $Y=510500
X3964 VDD VSS 4273 4274 SIGN_MEMCCOP $T=293790 509800 1 180 $X=291590 $Y=508800
X3965 VDD VSS 4275 4276 SIGN_MEMCCOP $T=292590 513200 1 0 $X=291590 $Y=510500
X3966 VDD VSS 4277 4278 SIGN_MEMCCOP $T=298590 509800 1 180 $X=296390 $Y=508800
X3967 VDD VSS 4279 4280 SIGN_MEMCCOP $T=297390 513200 1 0 $X=296390 $Y=510500
X3968 VDD VSS 4281 4282 SIGN_MEMCCOP $T=303390 509800 1 180 $X=301190 $Y=508800
X3969 VDD VSS 4283 4284 SIGN_MEMCCOP $T=302190 513200 1 0 $X=301190 $Y=510500
X3970 VDD VSS 4285 4286 SIGN_MEMCCOP $T=308190 509800 1 180 $X=305990 $Y=508800
X3971 VDD VSS 4287 4288 SIGN_MEMCCOP $T=306990 513200 1 0 $X=305990 $Y=510500
X3972 VDD VSS 4289 4290 SIGN_MEMCCOP $T=312990 509800 1 180 $X=310790 $Y=508800
X3973 VDD VSS 4291 4292 SIGN_MEMCCOP $T=311790 513200 1 0 $X=310790 $Y=510500
X3974 VDD VSS 4293 4294 SIGN_MEMCCOP $T=323790 509800 1 180 $X=321590 $Y=508800
X3975 VDD VSS 4295 4296 SIGN_MEMCCOP $T=322590 513200 1 0 $X=321590 $Y=510500
X3976 VDD VSS 4297 4298 SIGN_MEMCCOP $T=328590 509800 1 180 $X=326390 $Y=508800
X3977 VDD VSS 4299 4300 SIGN_MEMCCOP $T=327390 513200 1 0 $X=326390 $Y=510500
X3978 VDD VSS 4301 4302 SIGN_MEMCCOP $T=333390 509800 1 180 $X=331190 $Y=508800
X3979 VDD VSS 4303 4304 SIGN_MEMCCOP $T=332190 513200 1 0 $X=331190 $Y=510500
X3980 VDD VSS 4305 4306 SIGN_MEMCCOP $T=338190 509800 1 180 $X=335990 $Y=508800
X3981 VDD VSS 4307 4308 SIGN_MEMCCOP $T=336990 513200 1 0 $X=335990 $Y=510500
X3982 VDD VSS 4309 4310 SIGN_MEMCCOP $T=342990 509800 1 180 $X=340790 $Y=508800
X3983 VDD VSS 4311 4312 SIGN_MEMCCOP $T=341790 513200 1 0 $X=340790 $Y=510500
X3984 VDD VSS 4313 4314 SIGN_MEMCCOP $T=347790 509800 1 180 $X=345590 $Y=508800
X3985 VDD VSS 4315 4316 SIGN_MEMCCOP $T=346590 513200 1 0 $X=345590 $Y=510500
X3986 VDD VSS 4317 4318 SIGN_MEMCCOP $T=352590 509800 1 180 $X=350390 $Y=508800
X3987 VDD VSS 4319 4320 SIGN_MEMCCOP $T=351390 513200 1 0 $X=350390 $Y=510500
X3988 VDD VSS 4321 4322 SIGN_MEMCCOP $T=358590 509800 1 180 $X=356390 $Y=508800
X3989 VDD VSS 4323 4324 SIGN_MEMCCOP $T=357390 513200 1 0 $X=356390 $Y=510500
X3990 VDD VSS 4325 4326 SIGN_MEMCCOP $T=363390 509800 1 180 $X=361190 $Y=508800
X3991 VDD VSS 4327 4328 SIGN_MEMCCOP $T=362190 513200 1 0 $X=361190 $Y=510500
X3992 VDD VSS 4329 4330 SIGN_MEMCCOP $T=368190 509800 1 180 $X=365990 $Y=508800
X3993 VDD VSS 4331 4332 SIGN_MEMCCOP $T=366990 513200 1 0 $X=365990 $Y=510500
X3994 VDD VSS 4333 4334 SIGN_MEMCCOP $T=372990 509800 1 180 $X=370790 $Y=508800
X3995 VDD VSS 4335 4336 SIGN_MEMCCOP $T=371790 513200 1 0 $X=370790 $Y=510500
X3996 VDD VSS 4337 4338 SIGN_MEMCCOP $T=377790 509800 1 180 $X=375590 $Y=508800
X3997 VDD VSS 4339 4340 SIGN_MEMCCOP $T=376590 513200 1 0 $X=375590 $Y=510500
X3998 VDD VSS 4341 4342 SIGN_MEMCCOP $T=382590 509800 1 180 $X=380390 $Y=508800
X3999 VDD VSS 4343 4344 SIGN_MEMCCOP $T=381390 513200 1 0 $X=380390 $Y=510500
X4000 VDD VSS 4345 4346 SIGN_MEMCCOP $T=387390 509800 1 180 $X=385190 $Y=508800
X4001 VDD VSS 4347 4348 SIGN_MEMCCOP $T=386190 513200 1 0 $X=385190 $Y=510500
X4002 VDD VSS 4349 4350 SIGN_MEMCCOP $T=392190 509800 1 180 $X=389990 $Y=508800
X4003 VDD VSS 4351 4352 SIGN_MEMCCOP $T=390990 513200 1 0 $X=389990 $Y=510500
X4004 VDD VSS 4353 4354 SIGN_MEMCCEP $T=14810 509800 0 0 $X=13810 $Y=508800
X4005 VDD VSS 4355 4356 SIGN_MEMCCEP $T=16010 513200 0 180 $X=13810 $Y=510500
X4006 VDD VSS 4357 4358 SIGN_MEMCCEP $T=19610 509800 0 0 $X=18610 $Y=508800
X4007 VDD VSS 4359 4360 SIGN_MEMCCEP $T=20810 513200 0 180 $X=18610 $Y=510500
X4008 VDD VSS 4361 4362 SIGN_MEMCCEP $T=24410 509800 0 0 $X=23410 $Y=508800
X4009 VDD VSS 4363 4364 SIGN_MEMCCEP $T=25610 513200 0 180 $X=23410 $Y=510500
X4010 VDD VSS 4365 4366 SIGN_MEMCCEP $T=29210 509800 0 0 $X=28210 $Y=508800
X4011 VDD VSS 4367 4368 SIGN_MEMCCEP $T=30410 513200 0 180 $X=28210 $Y=510500
X4012 VDD VSS 4369 4370 SIGN_MEMCCEP $T=34010 509800 0 0 $X=33010 $Y=508800
X4013 VDD VSS 4371 4372 SIGN_MEMCCEP $T=35210 513200 0 180 $X=33010 $Y=510500
X4014 VDD VSS 4373 4374 SIGN_MEMCCEP $T=38810 509800 0 0 $X=37810 $Y=508800
X4015 VDD VSS 4375 4376 SIGN_MEMCCEP $T=40010 513200 0 180 $X=37810 $Y=510500
X4016 VDD VSS 4377 4378 SIGN_MEMCCEP $T=43610 509800 0 0 $X=42610 $Y=508800
X4017 VDD VSS 4379 4380 SIGN_MEMCCEP $T=44810 513200 0 180 $X=42610 $Y=510500
X4018 VDD VSS 4381 4382 SIGN_MEMCCEP $T=48410 509800 0 0 $X=47410 $Y=508800
X4019 VDD VSS 4383 4384 SIGN_MEMCCEP $T=49610 513200 0 180 $X=47410 $Y=510500
X4020 VDD VSS 4385 4386 SIGN_MEMCCEP $T=54410 509800 0 0 $X=53410 $Y=508800
X4021 VDD VSS 4387 4388 SIGN_MEMCCEP $T=55610 513200 0 180 $X=53410 $Y=510500
X4022 VDD VSS 4389 4390 SIGN_MEMCCEP $T=59210 509800 0 0 $X=58210 $Y=508800
X4023 VDD VSS 4391 4392 SIGN_MEMCCEP $T=60410 513200 0 180 $X=58210 $Y=510500
X4024 VDD VSS 4393 4394 SIGN_MEMCCEP $T=64010 509800 0 0 $X=63010 $Y=508800
X4025 VDD VSS 4395 4396 SIGN_MEMCCEP $T=65210 513200 0 180 $X=63010 $Y=510500
X4026 VDD VSS 4397 4398 SIGN_MEMCCEP $T=68810 509800 0 0 $X=67810 $Y=508800
X4027 VDD VSS 4399 4400 SIGN_MEMCCEP $T=70010 513200 0 180 $X=67810 $Y=510500
X4028 VDD VSS 4401 4402 SIGN_MEMCCEP $T=73610 509800 0 0 $X=72610 $Y=508800
X4029 VDD VSS 4403 4404 SIGN_MEMCCEP $T=74810 513200 0 180 $X=72610 $Y=510500
X4030 VDD VSS 4405 4406 SIGN_MEMCCEP $T=78410 509800 0 0 $X=77410 $Y=508800
X4031 VDD VSS 4407 4408 SIGN_MEMCCEP $T=79610 513200 0 180 $X=77410 $Y=510500
X4032 VDD VSS 4409 4410 SIGN_MEMCCEP $T=83210 509800 0 0 $X=82210 $Y=508800
X4033 VDD VSS 4411 4412 SIGN_MEMCCEP $T=84410 513200 0 180 $X=82210 $Y=510500
X4034 VDD VSS 4413 4414 SIGN_MEMCCEP $T=94010 509800 0 0 $X=93010 $Y=508800
X4035 VDD VSS 4415 4416 SIGN_MEMCCEP $T=95210 513200 0 180 $X=93010 $Y=510500
X4036 VDD VSS 4417 4418 SIGN_MEMCCEP $T=98810 509800 0 0 $X=97810 $Y=508800
X4037 VDD VSS 4419 4420 SIGN_MEMCCEP $T=100010 513200 0 180 $X=97810 $Y=510500
X4038 VDD VSS 4421 4422 SIGN_MEMCCEP $T=103610 509800 0 0 $X=102610 $Y=508800
X4039 VDD VSS 4423 4424 SIGN_MEMCCEP $T=104810 513200 0 180 $X=102610 $Y=510500
X4040 VDD VSS 4425 4426 SIGN_MEMCCEP $T=108410 509800 0 0 $X=107410 $Y=508800
X4041 VDD VSS 4427 4428 SIGN_MEMCCEP $T=109610 513200 0 180 $X=107410 $Y=510500
X4042 VDD VSS 4429 4430 SIGN_MEMCCEP $T=113210 509800 0 0 $X=112210 $Y=508800
X4043 VDD VSS 4431 4432 SIGN_MEMCCEP $T=114410 513200 0 180 $X=112210 $Y=510500
X4044 VDD VSS 4433 4434 SIGN_MEMCCEP $T=118010 509800 0 0 $X=117010 $Y=508800
X4045 VDD VSS 4435 4436 SIGN_MEMCCEP $T=119210 513200 0 180 $X=117010 $Y=510500
X4046 VDD VSS 4437 4438 SIGN_MEMCCEP $T=122810 509800 0 0 $X=121810 $Y=508800
X4047 VDD VSS 4439 4440 SIGN_MEMCCEP $T=124010 513200 0 180 $X=121810 $Y=510500
X4048 VDD VSS 4441 4442 SIGN_MEMCCEP $T=127610 509800 0 0 $X=126610 $Y=508800
X4049 VDD VSS 4443 4444 SIGN_MEMCCEP $T=128810 513200 0 180 $X=126610 $Y=510500
X4050 VDD VSS 4445 4446 SIGN_MEMCCEP $T=133610 509800 0 0 $X=132610 $Y=508800
X4051 VDD VSS 4447 4448 SIGN_MEMCCEP $T=134810 513200 0 180 $X=132610 $Y=510500
X4052 VDD VSS 4449 4450 SIGN_MEMCCEP $T=138410 509800 0 0 $X=137410 $Y=508800
X4053 VDD VSS 4451 4452 SIGN_MEMCCEP $T=139610 513200 0 180 $X=137410 $Y=510500
X4054 VDD VSS 4453 4454 SIGN_MEMCCEP $T=143210 509800 0 0 $X=142210 $Y=508800
X4055 VDD VSS 4455 4456 SIGN_MEMCCEP $T=144410 513200 0 180 $X=142210 $Y=510500
X4056 VDD VSS 4457 4458 SIGN_MEMCCEP $T=148010 509800 0 0 $X=147010 $Y=508800
X4057 VDD VSS 4459 4460 SIGN_MEMCCEP $T=149210 513200 0 180 $X=147010 $Y=510500
X4058 VDD VSS 4461 4462 SIGN_MEMCCEP $T=152810 509800 0 0 $X=151810 $Y=508800
X4059 VDD VSS 4463 4464 SIGN_MEMCCEP $T=154010 513200 0 180 $X=151810 $Y=510500
X4060 VDD VSS 4465 4466 SIGN_MEMCCEP $T=157610 509800 0 0 $X=156610 $Y=508800
X4061 VDD VSS 4467 4468 SIGN_MEMCCEP $T=158810 513200 0 180 $X=156610 $Y=510500
X4062 VDD VSS 4469 4470 SIGN_MEMCCEP $T=162410 509800 0 0 $X=161410 $Y=508800
X4063 VDD VSS 4471 4472 SIGN_MEMCCEP $T=163610 513200 0 180 $X=161410 $Y=510500
X4064 VDD VSS 4473 4474 SIGN_MEMCCEP $T=167210 509800 0 0 $X=166210 $Y=508800
X4065 VDD VSS 4475 4476 SIGN_MEMCCEP $T=168410 513200 0 180 $X=166210 $Y=510500
X4066 VDD VSS 4477 4478 SIGN_MEMCCEP $T=239790 509800 0 0 $X=238790 $Y=508800
X4067 VDD VSS 4479 4480 SIGN_MEMCCEP $T=240990 513200 0 180 $X=238790 $Y=510500
X4068 VDD VSS 4481 4482 SIGN_MEMCCEP $T=244590 509800 0 0 $X=243590 $Y=508800
X4069 VDD VSS 4483 4484 SIGN_MEMCCEP $T=245790 513200 0 180 $X=243590 $Y=510500
X4070 VDD VSS 4485 4486 SIGN_MEMCCEP $T=249390 509800 0 0 $X=248390 $Y=508800
X4071 VDD VSS 4487 4488 SIGN_MEMCCEP $T=250590 513200 0 180 $X=248390 $Y=510500
X4072 VDD VSS 4489 4490 SIGN_MEMCCEP $T=254190 509800 0 0 $X=253190 $Y=508800
X4073 VDD VSS 4491 4492 SIGN_MEMCCEP $T=255390 513200 0 180 $X=253190 $Y=510500
X4074 VDD VSS 4493 4494 SIGN_MEMCCEP $T=258990 509800 0 0 $X=257990 $Y=508800
X4075 VDD VSS 4495 4496 SIGN_MEMCCEP $T=260190 513200 0 180 $X=257990 $Y=510500
X4076 VDD VSS 4497 4498 SIGN_MEMCCEP $T=263790 509800 0 0 $X=262790 $Y=508800
X4077 VDD VSS 4499 4500 SIGN_MEMCCEP $T=264990 513200 0 180 $X=262790 $Y=510500
X4078 VDD VSS 4501 4502 SIGN_MEMCCEP $T=268590 509800 0 0 $X=267590 $Y=508800
X4079 VDD VSS 4503 4504 SIGN_MEMCCEP $T=269790 513200 0 180 $X=267590 $Y=510500
X4080 VDD VSS 4505 4506 SIGN_MEMCCEP $T=273390 509800 0 0 $X=272390 $Y=508800
X4081 VDD VSS 4507 4508 SIGN_MEMCCEP $T=274590 513200 0 180 $X=272390 $Y=510500
X4082 VDD VSS 4509 4510 SIGN_MEMCCEP $T=279390 509800 0 0 $X=278390 $Y=508800
X4083 VDD VSS 4511 4512 SIGN_MEMCCEP $T=280590 513200 0 180 $X=278390 $Y=510500
X4084 VDD VSS 4513 4514 SIGN_MEMCCEP $T=284190 509800 0 0 $X=283190 $Y=508800
X4085 VDD VSS 4515 4516 SIGN_MEMCCEP $T=285390 513200 0 180 $X=283190 $Y=510500
X4086 VDD VSS 4517 4518 SIGN_MEMCCEP $T=288990 509800 0 0 $X=287990 $Y=508800
X4087 VDD VSS 4519 4520 SIGN_MEMCCEP $T=290190 513200 0 180 $X=287990 $Y=510500
X4088 VDD VSS 4521 4522 SIGN_MEMCCEP $T=293790 509800 0 0 $X=292790 $Y=508800
X4089 VDD VSS 4523 4524 SIGN_MEMCCEP $T=294990 513200 0 180 $X=292790 $Y=510500
X4090 VDD VSS 4525 4526 SIGN_MEMCCEP $T=298590 509800 0 0 $X=297590 $Y=508800
X4091 VDD VSS 4527 4528 SIGN_MEMCCEP $T=299790 513200 0 180 $X=297590 $Y=510500
X4092 VDD VSS 4529 4530 SIGN_MEMCCEP $T=303390 509800 0 0 $X=302390 $Y=508800
X4093 VDD VSS 4531 4532 SIGN_MEMCCEP $T=304590 513200 0 180 $X=302390 $Y=510500
X4094 VDD VSS 4533 4534 SIGN_MEMCCEP $T=308190 509800 0 0 $X=307190 $Y=508800
X4095 VDD VSS 4535 4536 SIGN_MEMCCEP $T=309390 513200 0 180 $X=307190 $Y=510500
X4096 VDD VSS 4537 4538 SIGN_MEMCCEP $T=312990 509800 0 0 $X=311990 $Y=508800
X4097 VDD VSS 4539 4540 SIGN_MEMCCEP $T=314190 513200 0 180 $X=311990 $Y=510500
X4098 VDD VSS 4541 4542 SIGN_MEMCCEP $T=318990 509800 0 0 $X=317990 $Y=508800
X4099 VDD VSS 4543 4544 SIGN_MEMCCEP $T=320190 513200 0 180 $X=317990 $Y=510500
X4100 VDD VSS 4545 4546 SIGN_MEMCCEP $T=323790 509800 0 0 $X=322790 $Y=508800
X4101 VDD VSS 4547 4548 SIGN_MEMCCEP $T=324990 513200 0 180 $X=322790 $Y=510500
X4102 VDD VSS 4549 4550 SIGN_MEMCCEP $T=328590 509800 0 0 $X=327590 $Y=508800
X4103 VDD VSS 4551 4552 SIGN_MEMCCEP $T=329790 513200 0 180 $X=327590 $Y=510500
X4104 VDD VSS 4553 4554 SIGN_MEMCCEP $T=333390 509800 0 0 $X=332390 $Y=508800
X4105 VDD VSS 4555 4556 SIGN_MEMCCEP $T=334590 513200 0 180 $X=332390 $Y=510500
X4106 VDD VSS 4557 4558 SIGN_MEMCCEP $T=338190 509800 0 0 $X=337190 $Y=508800
X4107 VDD VSS 4559 4560 SIGN_MEMCCEP $T=339390 513200 0 180 $X=337190 $Y=510500
X4108 VDD VSS 4561 4562 SIGN_MEMCCEP $T=342990 509800 0 0 $X=341990 $Y=508800
X4109 VDD VSS 4563 4564 SIGN_MEMCCEP $T=344190 513200 0 180 $X=341990 $Y=510500
X4110 VDD VSS 4565 4566 SIGN_MEMCCEP $T=347790 509800 0 0 $X=346790 $Y=508800
X4111 VDD VSS 4567 4568 SIGN_MEMCCEP $T=348990 513200 0 180 $X=346790 $Y=510500
X4112 VDD VSS 4569 4570 SIGN_MEMCCEP $T=352590 509800 0 0 $X=351590 $Y=508800
X4113 VDD VSS 4571 4572 SIGN_MEMCCEP $T=353790 513200 0 180 $X=351590 $Y=510500
X4114 VDD VSS 4573 4574 SIGN_MEMCCEP $T=358590 509800 0 0 $X=357590 $Y=508800
X4115 VDD VSS 4575 4576 SIGN_MEMCCEP $T=359790 513200 0 180 $X=357590 $Y=510500
X4116 VDD VSS 4577 4578 SIGN_MEMCCEP $T=363390 509800 0 0 $X=362390 $Y=508800
X4117 VDD VSS 4579 4580 SIGN_MEMCCEP $T=364590 513200 0 180 $X=362390 $Y=510500
X4118 VDD VSS 4581 4582 SIGN_MEMCCEP $T=368190 509800 0 0 $X=367190 $Y=508800
X4119 VDD VSS 4583 4584 SIGN_MEMCCEP $T=369390 513200 0 180 $X=367190 $Y=510500
X4120 VDD VSS 4585 4586 SIGN_MEMCCEP $T=372990 509800 0 0 $X=371990 $Y=508800
X4121 VDD VSS 4587 4588 SIGN_MEMCCEP $T=374190 513200 0 180 $X=371990 $Y=510500
X4122 VDD VSS 4589 4590 SIGN_MEMCCEP $T=377790 509800 0 0 $X=376790 $Y=508800
X4123 VDD VSS 4591 4592 SIGN_MEMCCEP $T=378990 513200 0 180 $X=376790 $Y=510500
X4124 VDD VSS 4593 4594 SIGN_MEMCCEP $T=382590 509800 0 0 $X=381590 $Y=508800
X4125 VDD VSS 4595 4596 SIGN_MEMCCEP $T=383790 513200 0 180 $X=381590 $Y=510500
X4126 VDD VSS 4597 4598 SIGN_MEMCCEP $T=387390 509800 0 0 $X=386390 $Y=508800
X4127 VDD VSS 4599 4600 SIGN_MEMCCEP $T=388590 513200 0 180 $X=386390 $Y=510500
X4128 VDD VSS 4601 4602 SIGN_MEMCCEP $T=392190 509800 0 0 $X=391190 $Y=508800
X4129 VDD VSS 4603 4604 SIGN_MEMCCEP $T=393390 513200 0 180 $X=391190 $Y=510500
X4130 VSS VDD 4605 4606 SIGN_MEMCCOG $T=17210 509800 1 180 $X=15010 $Y=508800
X4131 VSS VDD 4607 4608 SIGN_MEMCCOG $T=16010 513200 1 0 $X=15010 $Y=510500
X4132 VSS VDD 4609 4610 SIGN_MEMCCOG $T=22010 509800 1 180 $X=19810 $Y=508800
X4133 VSS VDD 4611 4612 SIGN_MEMCCOG $T=20810 513200 1 0 $X=19810 $Y=510500
X4134 VSS VDD 4613 4614 SIGN_MEMCCOG $T=26810 509800 1 180 $X=24610 $Y=508800
X4135 VSS VDD 4615 4616 SIGN_MEMCCOG $T=25610 513200 1 0 $X=24610 $Y=510500
X4136 VSS VDD 4617 4618 SIGN_MEMCCOG $T=31610 509800 1 180 $X=29410 $Y=508800
X4137 VSS VDD 4619 4620 SIGN_MEMCCOG $T=30410 513200 1 0 $X=29410 $Y=510500
X4138 VSS VDD 4621 4622 SIGN_MEMCCOG $T=36410 509800 1 180 $X=34210 $Y=508800
X4139 VSS VDD 4623 4624 SIGN_MEMCCOG $T=35210 513200 1 0 $X=34210 $Y=510500
X4140 VSS VDD 4625 4626 SIGN_MEMCCOG $T=41210 509800 1 180 $X=39010 $Y=508800
X4141 VSS VDD 4627 4628 SIGN_MEMCCOG $T=40010 513200 1 0 $X=39010 $Y=510500
X4142 VSS VDD 4629 4630 SIGN_MEMCCOG $T=46010 509800 1 180 $X=43810 $Y=508800
X4143 VSS VDD 4631 4632 SIGN_MEMCCOG $T=44810 513200 1 0 $X=43810 $Y=510500
X4144 VSS VDD 4633 4634 SIGN_MEMCCOG $T=50810 509800 1 180 $X=48610 $Y=508800
X4145 VSS VDD 4635 4636 SIGN_MEMCCOG $T=49610 513200 1 0 $X=48610 $Y=510500
X4146 VSS VDD 4637 4638 SIGN_MEMCCOG $T=56810 509800 1 180 $X=54610 $Y=508800
X4147 VSS VDD 4639 4640 SIGN_MEMCCOG $T=55610 513200 1 0 $X=54610 $Y=510500
X4148 VSS VDD 4641 4642 SIGN_MEMCCOG $T=61610 509800 1 180 $X=59410 $Y=508800
X4149 VSS VDD 4643 4644 SIGN_MEMCCOG $T=60410 513200 1 0 $X=59410 $Y=510500
X4150 VSS VDD 4645 4646 SIGN_MEMCCOG $T=66410 509800 1 180 $X=64210 $Y=508800
X4151 VSS VDD 4647 4648 SIGN_MEMCCOG $T=65210 513200 1 0 $X=64210 $Y=510500
X4152 VSS VDD 4649 4650 SIGN_MEMCCOG $T=71210 509800 1 180 $X=69010 $Y=508800
X4153 VSS VDD 4651 4652 SIGN_MEMCCOG $T=70010 513200 1 0 $X=69010 $Y=510500
X4154 VSS VDD 4653 4654 SIGN_MEMCCOG $T=76010 509800 1 180 $X=73810 $Y=508800
X4155 VSS VDD 4655 4656 SIGN_MEMCCOG $T=74810 513200 1 0 $X=73810 $Y=510500
X4156 VSS VDD 4657 4658 SIGN_MEMCCOG $T=80810 509800 1 180 $X=78610 $Y=508800
X4157 VSS VDD 4659 4660 SIGN_MEMCCOG $T=79610 513200 1 0 $X=78610 $Y=510500
X4158 VSS VDD 4661 4662 SIGN_MEMCCOG $T=85610 509800 1 180 $X=83410 $Y=508800
X4159 VSS VDD 4663 4664 SIGN_MEMCCOG $T=84410 513200 1 0 $X=83410 $Y=510500
X4160 VSS VDD 4665 4666 SIGN_MEMCCOG $T=96410 509800 1 180 $X=94210 $Y=508800
X4161 VSS VDD 4667 4668 SIGN_MEMCCOG $T=95210 513200 1 0 $X=94210 $Y=510500
X4162 VSS VDD 4669 4670 SIGN_MEMCCOG $T=101210 509800 1 180 $X=99010 $Y=508800
X4163 VSS VDD 4671 4672 SIGN_MEMCCOG $T=100010 513200 1 0 $X=99010 $Y=510500
X4164 VSS VDD 4673 4674 SIGN_MEMCCOG $T=106010 509800 1 180 $X=103810 $Y=508800
X4165 VSS VDD 4675 4676 SIGN_MEMCCOG $T=104810 513200 1 0 $X=103810 $Y=510500
X4166 VSS VDD 4677 4678 SIGN_MEMCCOG $T=110810 509800 1 180 $X=108610 $Y=508800
X4167 VSS VDD 4679 4680 SIGN_MEMCCOG $T=109610 513200 1 0 $X=108610 $Y=510500
X4168 VSS VDD 4681 4682 SIGN_MEMCCOG $T=115610 509800 1 180 $X=113410 $Y=508800
X4169 VSS VDD 4683 4684 SIGN_MEMCCOG $T=114410 513200 1 0 $X=113410 $Y=510500
X4170 VSS VDD 4685 4686 SIGN_MEMCCOG $T=120410 509800 1 180 $X=118210 $Y=508800
X4171 VSS VDD 4687 4688 SIGN_MEMCCOG $T=119210 513200 1 0 $X=118210 $Y=510500
X4172 VSS VDD 4689 4690 SIGN_MEMCCOG $T=125210 509800 1 180 $X=123010 $Y=508800
X4173 VSS VDD 4691 4692 SIGN_MEMCCOG $T=124010 513200 1 0 $X=123010 $Y=510500
X4174 VSS VDD 4693 4694 SIGN_MEMCCOG $T=130010 509800 1 180 $X=127810 $Y=508800
X4175 VSS VDD 4695 4696 SIGN_MEMCCOG $T=128810 513200 1 0 $X=127810 $Y=510500
X4176 VSS VDD 4697 4698 SIGN_MEMCCOG $T=136010 509800 1 180 $X=133810 $Y=508800
X4177 VSS VDD 4699 4700 SIGN_MEMCCOG $T=134810 513200 1 0 $X=133810 $Y=510500
X4178 VSS VDD 4701 4702 SIGN_MEMCCOG $T=140810 509800 1 180 $X=138610 $Y=508800
X4179 VSS VDD 4703 4704 SIGN_MEMCCOG $T=139610 513200 1 0 $X=138610 $Y=510500
X4180 VSS VDD 4705 4706 SIGN_MEMCCOG $T=145610 509800 1 180 $X=143410 $Y=508800
X4181 VSS VDD 4707 4708 SIGN_MEMCCOG $T=144410 513200 1 0 $X=143410 $Y=510500
X4182 VSS VDD 4709 4710 SIGN_MEMCCOG $T=150410 509800 1 180 $X=148210 $Y=508800
X4183 VSS VDD 4711 4712 SIGN_MEMCCOG $T=149210 513200 1 0 $X=148210 $Y=510500
X4184 VSS VDD 4713 4714 SIGN_MEMCCOG $T=155210 509800 1 180 $X=153010 $Y=508800
X4185 VSS VDD 4715 4716 SIGN_MEMCCOG $T=154010 513200 1 0 $X=153010 $Y=510500
X4186 VSS VDD 4717 4718 SIGN_MEMCCOG $T=160010 509800 1 180 $X=157810 $Y=508800
X4187 VSS VDD 4719 4720 SIGN_MEMCCOG $T=158810 513200 1 0 $X=157810 $Y=510500
X4188 VSS VDD 4721 4722 SIGN_MEMCCOG $T=164810 509800 1 180 $X=162610 $Y=508800
X4189 VSS VDD 4723 4724 SIGN_MEMCCOG $T=163610 513200 1 0 $X=162610 $Y=510500
X4190 VSS VDD 4725 4726 SIGN_MEMCCOG $T=169610 509800 1 180 $X=167410 $Y=508800
X4191 VSS VDD 4727 4728 SIGN_MEMCCOG $T=168410 513200 1 0 $X=167410 $Y=510500
X4192 VSS VDD 4729 4730 SIGN_MEMCCOG $T=242190 509800 1 180 $X=239990 $Y=508800
X4193 VSS VDD 4731 4732 SIGN_MEMCCOG $T=240990 513200 1 0 $X=239990 $Y=510500
X4194 VSS VDD 4733 4734 SIGN_MEMCCOG $T=246990 509800 1 180 $X=244790 $Y=508800
X4195 VSS VDD 4735 4736 SIGN_MEMCCOG $T=245790 513200 1 0 $X=244790 $Y=510500
X4196 VSS VDD 4737 4738 SIGN_MEMCCOG $T=251790 509800 1 180 $X=249590 $Y=508800
X4197 VSS VDD 4739 4740 SIGN_MEMCCOG $T=250590 513200 1 0 $X=249590 $Y=510500
X4198 VSS VDD 4741 4742 SIGN_MEMCCOG $T=256590 509800 1 180 $X=254390 $Y=508800
X4199 VSS VDD 4743 4744 SIGN_MEMCCOG $T=255390 513200 1 0 $X=254390 $Y=510500
X4200 VSS VDD 4745 4746 SIGN_MEMCCOG $T=261390 509800 1 180 $X=259190 $Y=508800
X4201 VSS VDD 4747 4748 SIGN_MEMCCOG $T=260190 513200 1 0 $X=259190 $Y=510500
X4202 VSS VDD 4749 4750 SIGN_MEMCCOG $T=266190 509800 1 180 $X=263990 $Y=508800
X4203 VSS VDD 4751 4752 SIGN_MEMCCOG $T=264990 513200 1 0 $X=263990 $Y=510500
X4204 VSS VDD 4753 4754 SIGN_MEMCCOG $T=270990 509800 1 180 $X=268790 $Y=508800
X4205 VSS VDD 4755 4756 SIGN_MEMCCOG $T=269790 513200 1 0 $X=268790 $Y=510500
X4206 VSS VDD 4757 4758 SIGN_MEMCCOG $T=275790 509800 1 180 $X=273590 $Y=508800
X4207 VSS VDD 4759 4760 SIGN_MEMCCOG $T=274590 513200 1 0 $X=273590 $Y=510500
X4208 VSS VDD 4761 4762 SIGN_MEMCCOG $T=281790 509800 1 180 $X=279590 $Y=508800
X4209 VSS VDD 4763 4764 SIGN_MEMCCOG $T=280590 513200 1 0 $X=279590 $Y=510500
X4210 VSS VDD 4765 4766 SIGN_MEMCCOG $T=286590 509800 1 180 $X=284390 $Y=508800
X4211 VSS VDD 4767 4768 SIGN_MEMCCOG $T=285390 513200 1 0 $X=284390 $Y=510500
X4212 VSS VDD 4769 4770 SIGN_MEMCCOG $T=291390 509800 1 180 $X=289190 $Y=508800
X4213 VSS VDD 4771 4772 SIGN_MEMCCOG $T=290190 513200 1 0 $X=289190 $Y=510500
X4214 VSS VDD 4773 4774 SIGN_MEMCCOG $T=296190 509800 1 180 $X=293990 $Y=508800
X4215 VSS VDD 4775 4776 SIGN_MEMCCOG $T=294990 513200 1 0 $X=293990 $Y=510500
X4216 VSS VDD 4777 4778 SIGN_MEMCCOG $T=300990 509800 1 180 $X=298790 $Y=508800
X4217 VSS VDD 4779 4780 SIGN_MEMCCOG $T=299790 513200 1 0 $X=298790 $Y=510500
X4218 VSS VDD 4781 4782 SIGN_MEMCCOG $T=305790 509800 1 180 $X=303590 $Y=508800
X4219 VSS VDD 4783 4784 SIGN_MEMCCOG $T=304590 513200 1 0 $X=303590 $Y=510500
X4220 VSS VDD 4785 4786 SIGN_MEMCCOG $T=310590 509800 1 180 $X=308390 $Y=508800
X4221 VSS VDD 4787 4788 SIGN_MEMCCOG $T=309390 513200 1 0 $X=308390 $Y=510500
X4222 VSS VDD 4789 4790 SIGN_MEMCCOG $T=315390 509800 1 180 $X=313190 $Y=508800
X4223 VSS VDD 4791 4792 SIGN_MEMCCOG $T=314190 513200 1 0 $X=313190 $Y=510500
X4224 VSS VDD 4793 4794 SIGN_MEMCCOG $T=321390 509800 1 180 $X=319190 $Y=508800
X4225 VSS VDD 4795 4796 SIGN_MEMCCOG $T=320190 513200 1 0 $X=319190 $Y=510500
X4226 VSS VDD 4797 4798 SIGN_MEMCCOG $T=326190 509800 1 180 $X=323990 $Y=508800
X4227 VSS VDD 4799 4800 SIGN_MEMCCOG $T=324990 513200 1 0 $X=323990 $Y=510500
X4228 VSS VDD 4801 4802 SIGN_MEMCCOG $T=330990 509800 1 180 $X=328790 $Y=508800
X4229 VSS VDD 4803 4804 SIGN_MEMCCOG $T=329790 513200 1 0 $X=328790 $Y=510500
X4230 VSS VDD 4805 4806 SIGN_MEMCCOG $T=335790 509800 1 180 $X=333590 $Y=508800
X4231 VSS VDD 4807 4808 SIGN_MEMCCOG $T=334590 513200 1 0 $X=333590 $Y=510500
X4232 VSS VDD 4809 4810 SIGN_MEMCCOG $T=340590 509800 1 180 $X=338390 $Y=508800
X4233 VSS VDD 4811 4812 SIGN_MEMCCOG $T=339390 513200 1 0 $X=338390 $Y=510500
X4234 VSS VDD 4813 4814 SIGN_MEMCCOG $T=345390 509800 1 180 $X=343190 $Y=508800
X4235 VSS VDD 4815 4816 SIGN_MEMCCOG $T=344190 513200 1 0 $X=343190 $Y=510500
X4236 VSS VDD 4817 4818 SIGN_MEMCCOG $T=350190 509800 1 180 $X=347990 $Y=508800
X4237 VSS VDD 4819 4820 SIGN_MEMCCOG $T=348990 513200 1 0 $X=347990 $Y=510500
X4238 VSS VDD 4821 4822 SIGN_MEMCCOG $T=354990 509800 1 180 $X=352790 $Y=508800
X4239 VSS VDD 4823 4824 SIGN_MEMCCOG $T=353790 513200 1 0 $X=352790 $Y=510500
X4240 VSS VDD 4825 4826 SIGN_MEMCCOG $T=360990 509800 1 180 $X=358790 $Y=508800
X4241 VSS VDD 4827 4828 SIGN_MEMCCOG $T=359790 513200 1 0 $X=358790 $Y=510500
X4242 VSS VDD 4829 4830 SIGN_MEMCCOG $T=365790 509800 1 180 $X=363590 $Y=508800
X4243 VSS VDD 4831 4832 SIGN_MEMCCOG $T=364590 513200 1 0 $X=363590 $Y=510500
X4244 VSS VDD 4833 4834 SIGN_MEMCCOG $T=370590 509800 1 180 $X=368390 $Y=508800
X4245 VSS VDD 4835 4836 SIGN_MEMCCOG $T=369390 513200 1 0 $X=368390 $Y=510500
X4246 VSS VDD 4837 4838 SIGN_MEMCCOG $T=375390 509800 1 180 $X=373190 $Y=508800
X4247 VSS VDD 4839 4840 SIGN_MEMCCOG $T=374190 513200 1 0 $X=373190 $Y=510500
X4248 VSS VDD 4841 4842 SIGN_MEMCCOG $T=380190 509800 1 180 $X=377990 $Y=508800
X4249 VSS VDD 4843 4844 SIGN_MEMCCOG $T=378990 513200 1 0 $X=377990 $Y=510500
X4250 VSS VDD 4845 4846 SIGN_MEMCCOG $T=384990 509800 1 180 $X=382790 $Y=508800
X4251 VSS VDD 4847 4848 SIGN_MEMCCOG $T=383790 513200 1 0 $X=382790 $Y=510500
X4252 VSS VDD 4849 4850 SIGN_MEMCCOG $T=389790 509800 1 180 $X=387590 $Y=508800
X4253 VSS VDD 4851 4852 SIGN_MEMCCOG $T=388590 513200 1 0 $X=387590 $Y=510500
X4254 VSS VDD 4853 4854 SIGN_MEMCCOG $T=394590 509800 1 180 $X=392390 $Y=508800
X4255 VSS VDD 4855 4856 SIGN_MEMCCOG $T=393390 513200 1 0 $X=392390 $Y=510500
X4256 VSS VSS 864 865 SIGN_MEMFLCCSTRAP $T=52010 509800 1 180 $X=49810 $Y=508800
X4257 VSS VSS 864 865 SIGN_MEMFLCCSTRAP $T=52010 513200 0 180 $X=49810 $Y=510500
X4258 VSS 50 866 867 SIGN_MEMFLCCSTRAP $T=91610 509800 1 180 $X=89410 $Y=508800
X4259 VSS 50 866 867 SIGN_MEMFLCCSTRAP $T=91610 513200 0 180 $X=89410 $Y=510500
X4260 VSS 50 868 869 SIGN_MEMFLCCSTRAP $T=131210 509800 1 180 $X=129010 $Y=508800
X4261 VSS 50 868 869 SIGN_MEMFLCCSTRAP $T=131210 513200 0 180 $X=129010 $Y=510500
X4262 VSS 50 870 871 SIGN_MEMFLCCSTRAP $T=275790 509800 0 0 $X=274790 $Y=508800
X4263 VSS 50 870 871 SIGN_MEMFLCCSTRAP $T=275790 513200 1 0 $X=274790 $Y=510500
X4264 VSS 50 872 873 SIGN_MEMFLCCSTRAP $T=315390 509800 0 0 $X=314390 $Y=508800
X4265 VSS 50 872 873 SIGN_MEMFLCCSTRAP $T=315390 513200 1 0 $X=314390 $Y=510500
X4266 VSS VSS 874 875 SIGN_MEMFLCCSTRAP $T=354990 509800 0 0 $X=353990 $Y=508800
X4267 VSS VSS 874 875 SIGN_MEMFLCCSTRAP $T=354990 513200 1 0 $X=353990 $Y=510500
X4268 VDD VSS D<7> Q<7> D<6> Q<6> D<5> Q<5> D<4> Q<4> D<3> Q<3> D<2> Q<2> D<1> Q<1> D<0> Q<0> 51 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263
+ 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283
+ 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303
+ 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 323 VSS 324 325 326
+ 327 328 329 330 331 332 333 4857 4858 4859 4860 4861 4862 4863 4864 4865 4866 4867 4868 4869
+ 4870 4871 4872 4873 4874 4875 4876 4877 4878 4879 4880 4881 4882 4883 4884 4885 4886 4887 4888 4889
+ 4890 4891 4892 4893 4894 4895 4896 4897 4898 4899 4900 4901 4902 4903 4904 4905 4906 4907 4908 4909
+ 4910 4911 4912 4913 4914 4915 4916 4917 4918 4919 4920 4921 4922 4923 4924 4925 4926 4927 4928 4929
+ 4930 4931 4932 4933 4934 4935 4936 4937 4938 4939 4940 4941 4942 4943 4944 4945 4946 4947 4948 4949
+ 4950 4951 4952 4953 4954 4955 4956 4957 4958 4959 4960 4961 4962 4963 4964 4965 4966 4967 4968 4969
+ 4970 4971 4972 4973 4974 4975 4976 4977 4978 4979 4980 4981 4982 4983 4984 4985 4986 4987 4988 4989
+ 4990 4991 4992 4993 4994 4995 4996 4997 4998 4999 5000 5001 5002 5003 5004 5005 5006 5007 5008 5009
+ 5010 5011 5012 5013 5014 5015 5016 5017 5018 5019 5020 5021 5022 5023 5024 5025 5026 5027 5028 5029
+ 5030 5031 5032 5033 5034 5035 5036 5037 5038 5039 5040 5041 5042 5043 5044 5045 5046 5047 5048 5049
+ 5050 5051 5052 5053 5054 5055 5056 5057 5058 5059 5060 5061 5062 5063 5064 5065 5066 5067 5068 5069
+ 5070 5071 5072 5073 5074 5075 5076 5077 5078 5079 5080 5081 5082 5083 5084 5085 5086 5087 5088 5089
+ 5090 5091 5092 5093 5094 5095 5096 5097 5098 5099 5100 5101 5102 5103 5104 5105 5106 5107 5108 5109
+ 5110 5111 5112 5113 5114 5115 5116 5117 5118 5119 5120 5121 5122 5123 5124 5125 5126 5127 5128 5129
+ 5130 5131 5132 5133 5134 5135 5136 5137 5138 5139 5140 5141 5142 5143 5144 5145 5146 5147 5148 5149
+ 5150 5151 5152 5153 5154 5155 5156 5157 5158 5159 5160 5161 5162 5163 5164 5165 5166 5167 5168 5169
+ 5170 5171 5172 5173 5174 5175 5176 5177 5178 5179 5180 5181 5182 5183 5184 5185 5186 5187 5188 5189
+ 5190 5191 5192 5193 5194 5195 5196 5197 5198 5199 5200 5201 5202 5203 5204 5205 5206 5207 5208 5209
+ 5210 5211 5212 5213 5214 5215 5216 5217 5218 5219 5220 5221 5222 5223 5224 5225 5226 5227 5228 5229
+ 5230 5231 5232 5233 5234 5235 5236 5237 5238 5239 5240 5241 5242 5243 5244 5245 5246 5247 5248 5249
+ 5250 5251 5252 5253 5254 5255 5256 5257 5258 5259 5260 5261 5262 5263 5264 5265 5266 5267 5268 5269
+ 5270 5271 5272 5273 5274 5275 5276 5277 5278 5279 5280 5281 5282 5283 5284 5285 5286 5287 5288 5289
+ 5290 5291 5292 5293 5294 5295 5296 5297 5298 5299 5300 5301 5302 5303 5304 5305 5306 5307 5308 5309
+ 5310 5311 5312 5313 5314 5315 5316 5317 5318 5319 5320 5321 5322 5323 5324 5325 5326 5327 5328 5329
+ 5330 5331 5332 5333 5334 5335 5336 5337 5338 5339 5340 5341 5342 5343 5344 5345 5346 5347 5348 5349
+ 5350 5351 5352 5353 5354 5355 5356 5357 5358 5359 5360 5361 5362 5363 5364 5365 5366 5367 5368 5369
+ 5370
+ SIGN_MEMWING_8_LEFT $T=169610 10240 1 180 $X=11410 $Y=9240
X4333 VSS VDD 5371 5372 base_flmo_nvpv $T=90410 509800 1 180 $X=88210 $Y=508800
X4334 VSS VDD 5373 5374 base_flmo_nvpv $T=89210 513200 1 0 $X=88210 $Y=510500
X4466 VSS A<11> VDD 52 55 VSS ai $T=172010 10240 0 0 $X=171010 $Y=9240
X4467 VSS A<10> VDD 59 56 VSS ai $T=178810 10240 1 180 $X=174410 $Y=9240
X4468 VSS VDD 53 54 334 334 VSS 59 56 55 ap $T=172010 19280 0 0 $X=171010 $Y=18280
X4469 VSS VDD 57 58 334 334 VSS 59 56 52 ap $T=178810 19280 1 180 $X=174410 $Y=18280
X4470 VSS VDD 53 54 57 58 63 64 50 126 125 853 854 855 856 857 858 859 860 51
+ 190 189 254 253 318 317 124 123 122 121 188 187 186 185 252 251 250 249 316 315
+ 314 313 120 119 118 117 116 115 114 113 184 183 182 181 180 179 178 177 248 247
+ 246 245 244 243 242 241 312 311 310 309 308 307 306 305 112 111 110 109 108 107
+ 106 105 104 103 102 101 100 99 98 97 176 175 174 173 172 171 170 169 168 167
+ 166 165 164 163 162 161 240 239 238 237 236 235 234 233 232 231 230 229 228 227
+ 226 225 304 303 302 301 300 299 298 297 296 295 294 293 292 291 290 289 96 95
+ 94 93 92 91 90 89 88 87 86 85 84 83 82 81 80 79 78 77 76 75
+ 74 73 72 71 70 69 68 67 66 65 160 159 158 157 156 155 154 153 152 151
+ 150 149 148 147 146 145 144 143 142 141 140 139 138 137 136 135 134 133 132 131
+ 130 129 224 223 222 221 220 219 218 217 216 215 214 213 212 211 210 209 208 207
+ 206 205 204 203 202 201 200 199 198 197 196 195 194 193 288 287 286 285 284 283
+ 282 281 280 279 278 277 276 275 274 273 272 271 270 269 268 267 266 265 264 263
+ 262 261 260 259 258 257 127 128 191 192 255 256 61 50 60 845 846 847 848 849
+ 850 851 852
+ SIGN_MEMWORD_ROWS $T=172010 70630 0 0 $X=171010 $Y=69630
X4471 VSS VDD A<9> A<8> A<7> 845 846 847 848 849 850 851 852 VSS 334 334 SIGN_MEMHXP38X $T=178810 10240 0 0 $X=177810 $Y=9240
X4472 VSS VDD A<6> A<5> A<4> 853 854 855 856 857 858 859 860 VSS 334 334 SIGN_MEMHXP38X $T=192410 10240 0 0 $X=191410 $Y=9240
X4473 VSS VDD A<3> A<2> A<1> 326 327 328 329 330 331 332 333 VSS 334 334 SIGN_MEMHYP38X $T=206010 10240 0 0 $X=205010 $Y=9240
X4474 VSS VDD A<0> 324 325 334 VSS SIGN_MEMHYP12RX $T=219610 10240 0 0 $X=218610 $Y=9240
X4475 VDD VSS CEN WEN CLK 323 62 51 61 335 336 SIGN_MEMHBFX $T=224190 10240 0 0 $X=223190 $Y=9240
X4476 VDD VSS 336 335 CLK 62 334 51 51 51 51 SIGN_MEMCLK_DRVS $T=224190 37260 0 0 $X=223190 $Y=36260
X4477 VSS 876 SIGN_MEMFLCCMBLST2 $T=233790 73560 0 0 $X=232790 $Y=72560
X4478 VSS 876 SIGN_MEMFLCCMBLST2 $T=233790 76960 1 0 $X=232790 $Y=74260
X4479 VSS 877 SIGN_MEMFLCCMBLST2 $T=233790 76960 0 0 $X=232790 $Y=75960
X4480 VSS 877 SIGN_MEMFLCCMBLST2 $T=233790 80360 1 0 $X=232790 $Y=77660
X4481 VSS 878 SIGN_MEMFLCCMBLST2 $T=233790 80360 0 0 $X=232790 $Y=79360
X4482 VSS 878 SIGN_MEMFLCCMBLST2 $T=233790 83760 1 0 $X=232790 $Y=81060
X4483 VSS 879 SIGN_MEMFLCCMBLST2 $T=233790 83760 0 0 $X=232790 $Y=82760
X4484 VSS 879 SIGN_MEMFLCCMBLST2 $T=233790 87160 1 0 $X=232790 $Y=84460
X4485 VSS 880 SIGN_MEMFLCCMBLST2 $T=233790 87160 0 0 $X=232790 $Y=86160
X4486 VSS 880 SIGN_MEMFLCCMBLST2 $T=233790 90560 1 0 $X=232790 $Y=87860
X4487 VSS 881 SIGN_MEMFLCCMBLST2 $T=233790 90560 0 0 $X=232790 $Y=89560
X4488 VSS 881 SIGN_MEMFLCCMBLST2 $T=233790 93960 1 0 $X=232790 $Y=91260
X4489 VSS 882 SIGN_MEMFLCCMBLST2 $T=233790 93960 0 0 $X=232790 $Y=92960
X4490 VSS 882 SIGN_MEMFLCCMBLST2 $T=233790 97360 1 0 $X=232790 $Y=94660
X4491 VSS 883 SIGN_MEMFLCCMBLST2 $T=233790 97360 0 0 $X=232790 $Y=96360
X4492 VSS 883 SIGN_MEMFLCCMBLST2 $T=233790 100760 1 0 $X=232790 $Y=98060
X4493 VSS 884 SIGN_MEMFLCCMBLST2 $T=233790 100760 0 0 $X=232790 $Y=99760
X4494 VSS 884 SIGN_MEMFLCCMBLST2 $T=233790 104160 1 0 $X=232790 $Y=101460
X4495 VSS 885 SIGN_MEMFLCCMBLST2 $T=233790 104160 0 0 $X=232790 $Y=103160
X4496 VSS 885 SIGN_MEMFLCCMBLST2 $T=233790 107560 1 0 $X=232790 $Y=104860
X4497 VSS 886 SIGN_MEMFLCCMBLST2 $T=233790 107560 0 0 $X=232790 $Y=106560
X4498 VSS 886 SIGN_MEMFLCCMBLST2 $T=233790 110960 1 0 $X=232790 $Y=108260
X4499 VSS 887 SIGN_MEMFLCCMBLST2 $T=233790 110960 0 0 $X=232790 $Y=109960
X4500 VSS 887 SIGN_MEMFLCCMBLST2 $T=233790 114360 1 0 $X=232790 $Y=111660
X4501 VSS 888 SIGN_MEMFLCCMBLST2 $T=233790 114360 0 0 $X=232790 $Y=113360
X4502 VSS 888 SIGN_MEMFLCCMBLST2 $T=233790 117760 1 0 $X=232790 $Y=115060
X4503 VSS 889 SIGN_MEMFLCCMBLST2 $T=233790 117760 0 0 $X=232790 $Y=116760
X4504 VSS 889 SIGN_MEMFLCCMBLST2 $T=233790 121160 1 0 $X=232790 $Y=118460
X4505 VSS 890 SIGN_MEMFLCCMBLST2 $T=233790 121160 0 0 $X=232790 $Y=120160
X4506 VSS 890 SIGN_MEMFLCCMBLST2 $T=233790 124560 1 0 $X=232790 $Y=121860
X4507 VSS 891 SIGN_MEMFLCCMBLST2 $T=233790 124560 0 0 $X=232790 $Y=123560
X4508 VSS 891 SIGN_MEMFLCCMBLST2 $T=233790 127960 1 0 $X=232790 $Y=125260
X4509 VSS 892 SIGN_MEMFLCCMBLST2 $T=233790 127960 0 0 $X=232790 $Y=126960
X4510 VSS 892 SIGN_MEMFLCCMBLST2 $T=233790 131360 1 0 $X=232790 $Y=128660
X4511 VSS 893 SIGN_MEMFLCCMBLST2 $T=233790 131360 0 0 $X=232790 $Y=130360
X4512 VSS 893 SIGN_MEMFLCCMBLST2 $T=233790 134760 1 0 $X=232790 $Y=132060
X4513 VSS 894 SIGN_MEMFLCCMBLST2 $T=233790 134760 0 0 $X=232790 $Y=133760
X4514 VSS 894 SIGN_MEMFLCCMBLST2 $T=233790 138160 1 0 $X=232790 $Y=135460
X4515 VSS 895 SIGN_MEMFLCCMBLST2 $T=233790 138160 0 0 $X=232790 $Y=137160
X4516 VSS 895 SIGN_MEMFLCCMBLST2 $T=233790 141560 1 0 $X=232790 $Y=138860
X4517 VSS 896 SIGN_MEMFLCCMBLST2 $T=233790 141560 0 0 $X=232790 $Y=140560
X4518 VSS 896 SIGN_MEMFLCCMBLST2 $T=233790 144960 1 0 $X=232790 $Y=142260
X4519 VSS 897 SIGN_MEMFLCCMBLST2 $T=233790 144960 0 0 $X=232790 $Y=143960
X4520 VSS 897 SIGN_MEMFLCCMBLST2 $T=233790 148360 1 0 $X=232790 $Y=145660
X4521 VSS 898 SIGN_MEMFLCCMBLST2 $T=233790 148360 0 0 $X=232790 $Y=147360
X4522 VSS 898 SIGN_MEMFLCCMBLST2 $T=233790 151760 1 0 $X=232790 $Y=149060
X4523 VSS 899 SIGN_MEMFLCCMBLST2 $T=233790 151760 0 0 $X=232790 $Y=150760
X4524 VSS 899 SIGN_MEMFLCCMBLST2 $T=233790 155160 1 0 $X=232790 $Y=152460
X4525 VSS 900 SIGN_MEMFLCCMBLST2 $T=233790 155160 0 0 $X=232790 $Y=154160
X4526 VSS 900 SIGN_MEMFLCCMBLST2 $T=233790 158560 1 0 $X=232790 $Y=155860
X4527 VSS 901 SIGN_MEMFLCCMBLST2 $T=233790 158560 0 0 $X=232790 $Y=157560
X4528 VSS 901 SIGN_MEMFLCCMBLST2 $T=233790 161960 1 0 $X=232790 $Y=159260
X4529 VSS 902 SIGN_MEMFLCCMBLST2 $T=233790 161960 0 0 $X=232790 $Y=160960
X4530 VSS 902 SIGN_MEMFLCCMBLST2 $T=233790 165360 1 0 $X=232790 $Y=162660
X4531 VSS 903 SIGN_MEMFLCCMBLST2 $T=233790 165360 0 0 $X=232790 $Y=164360
X4532 VSS 903 SIGN_MEMFLCCMBLST2 $T=233790 168760 1 0 $X=232790 $Y=166060
X4533 VSS 904 SIGN_MEMFLCCMBLST2 $T=233790 168760 0 0 $X=232790 $Y=167760
X4534 VSS 904 SIGN_MEMFLCCMBLST2 $T=233790 172160 1 0 $X=232790 $Y=169460
X4535 VSS 905 SIGN_MEMFLCCMBLST2 $T=233790 172160 0 0 $X=232790 $Y=171160
X4536 VSS 905 SIGN_MEMFLCCMBLST2 $T=233790 175560 1 0 $X=232790 $Y=172860
X4537 VSS 906 SIGN_MEMFLCCMBLST2 $T=233790 175560 0 0 $X=232790 $Y=174560
X4538 VSS 906 SIGN_MEMFLCCMBLST2 $T=233790 178960 1 0 $X=232790 $Y=176260
X4539 VSS 907 SIGN_MEMFLCCMBLST2 $T=233790 178960 0 0 $X=232790 $Y=177960
X4540 VSS 907 SIGN_MEMFLCCMBLST2 $T=233790 182360 1 0 $X=232790 $Y=179660
X4541 VSS 908 SIGN_MEMFLCCMBLST2 $T=233790 182360 0 0 $X=232790 $Y=181360
X4542 VSS 908 SIGN_MEMFLCCMBLST2 $T=233790 185760 1 0 $X=232790 $Y=183060
X4543 VSS 909 SIGN_MEMFLCCMBLST2 $T=233790 185760 0 0 $X=232790 $Y=184760
X4544 VSS 909 SIGN_MEMFLCCMBLST2 $T=233790 189160 1 0 $X=232790 $Y=186460
X4545 VSS 910 SIGN_MEMFLCCMBLST2 $T=233790 189160 0 0 $X=232790 $Y=188160
X4546 VSS 910 SIGN_MEMFLCCMBLST2 $T=233790 192560 1 0 $X=232790 $Y=189860
X4547 VSS 911 SIGN_MEMFLCCMBLST2 $T=233790 192560 0 0 $X=232790 $Y=191560
X4548 VSS 911 SIGN_MEMFLCCMBLST2 $T=233790 195960 1 0 $X=232790 $Y=193260
X4549 VSS 912 SIGN_MEMFLCCMBLST2 $T=233790 195960 0 0 $X=232790 $Y=194960
X4550 VSS 912 SIGN_MEMFLCCMBLST2 $T=233790 199360 1 0 $X=232790 $Y=196660
X4551 VSS 913 SIGN_MEMFLCCMBLST2 $T=233790 199360 0 0 $X=232790 $Y=198360
X4552 VSS 913 SIGN_MEMFLCCMBLST2 $T=233790 202760 1 0 $X=232790 $Y=200060
X4553 VSS 914 SIGN_MEMFLCCMBLST2 $T=233790 202760 0 0 $X=232790 $Y=201760
X4554 VSS 914 SIGN_MEMFLCCMBLST2 $T=233790 206160 1 0 $X=232790 $Y=203460
X4555 VSS 915 SIGN_MEMFLCCMBLST2 $T=233790 206160 0 0 $X=232790 $Y=205160
X4556 VSS 915 SIGN_MEMFLCCMBLST2 $T=233790 209560 1 0 $X=232790 $Y=206860
X4557 VSS 916 SIGN_MEMFLCCMBLST2 $T=233790 209560 0 0 $X=232790 $Y=208560
X4558 VSS 916 SIGN_MEMFLCCMBLST2 $T=233790 212960 1 0 $X=232790 $Y=210260
X4559 VSS 917 SIGN_MEMFLCCMBLST2 $T=233790 212960 0 0 $X=232790 $Y=211960
X4560 VSS 917 SIGN_MEMFLCCMBLST2 $T=233790 216360 1 0 $X=232790 $Y=213660
X4561 VSS 918 SIGN_MEMFLCCMBLST2 $T=233790 216360 0 0 $X=232790 $Y=215360
X4562 VSS 918 SIGN_MEMFLCCMBLST2 $T=233790 219760 1 0 $X=232790 $Y=217060
X4563 VSS 919 SIGN_MEMFLCCMBLST2 $T=233790 219760 0 0 $X=232790 $Y=218760
X4564 VSS 919 SIGN_MEMFLCCMBLST2 $T=233790 223160 1 0 $X=232790 $Y=220460
X4565 VSS 920 SIGN_MEMFLCCMBLST2 $T=233790 223160 0 0 $X=232790 $Y=222160
X4566 VSS 920 SIGN_MEMFLCCMBLST2 $T=233790 226560 1 0 $X=232790 $Y=223860
X4567 VSS 921 SIGN_MEMFLCCMBLST2 $T=233790 226560 0 0 $X=232790 $Y=225560
X4568 VSS 921 SIGN_MEMFLCCMBLST2 $T=233790 229960 1 0 $X=232790 $Y=227260
X4569 VSS 922 SIGN_MEMFLCCMBLST2 $T=233790 229960 0 0 $X=232790 $Y=228960
X4570 VSS 922 SIGN_MEMFLCCMBLST2 $T=233790 233360 1 0 $X=232790 $Y=230660
X4571 VSS 923 SIGN_MEMFLCCMBLST2 $T=233790 233360 0 0 $X=232790 $Y=232360
X4572 VSS 923 SIGN_MEMFLCCMBLST2 $T=233790 236760 1 0 $X=232790 $Y=234060
X4573 VSS 924 SIGN_MEMFLCCMBLST2 $T=233790 236760 0 0 $X=232790 $Y=235760
X4574 VSS 924 SIGN_MEMFLCCMBLST2 $T=233790 240160 1 0 $X=232790 $Y=237460
X4575 VSS 925 SIGN_MEMFLCCMBLST2 $T=233790 240160 0 0 $X=232790 $Y=239160
X4576 VSS 925 SIGN_MEMFLCCMBLST2 $T=233790 243560 1 0 $X=232790 $Y=240860
X4577 VSS 926 SIGN_MEMFLCCMBLST2 $T=233790 243560 0 0 $X=232790 $Y=242560
X4578 VSS 926 SIGN_MEMFLCCMBLST2 $T=233790 246960 1 0 $X=232790 $Y=244260
X4579 VSS 927 SIGN_MEMFLCCMBLST2 $T=233790 246960 0 0 $X=232790 $Y=245960
X4580 VSS 927 SIGN_MEMFLCCMBLST2 $T=233790 250360 1 0 $X=232790 $Y=247660
X4581 VSS 928 SIGN_MEMFLCCMBLST2 $T=233790 250360 0 0 $X=232790 $Y=249360
X4582 VSS 928 SIGN_MEMFLCCMBLST2 $T=233790 253760 1 0 $X=232790 $Y=251060
X4583 VSS 929 SIGN_MEMFLCCMBLST2 $T=233790 253760 0 0 $X=232790 $Y=252760
X4584 VSS 929 SIGN_MEMFLCCMBLST2 $T=233790 257160 1 0 $X=232790 $Y=254460
X4585 VSS 930 SIGN_MEMFLCCMBLST2 $T=233790 257160 0 0 $X=232790 $Y=256160
X4586 VSS 930 SIGN_MEMFLCCMBLST2 $T=233790 260560 1 0 $X=232790 $Y=257860
X4587 VSS 931 SIGN_MEMFLCCMBLST2 $T=233790 260560 0 0 $X=232790 $Y=259560
X4588 VSS 931 SIGN_MEMFLCCMBLST2 $T=233790 263960 1 0 $X=232790 $Y=261260
X4589 VSS 932 SIGN_MEMFLCCMBLST2 $T=233790 263960 0 0 $X=232790 $Y=262960
X4590 VSS 932 SIGN_MEMFLCCMBLST2 $T=233790 267360 1 0 $X=232790 $Y=264660
X4591 VSS 933 SIGN_MEMFLCCMBLST2 $T=233790 267360 0 0 $X=232790 $Y=266360
X4592 VSS 933 SIGN_MEMFLCCMBLST2 $T=233790 270760 1 0 $X=232790 $Y=268060
X4593 VSS 934 SIGN_MEMFLCCMBLST2 $T=233790 270760 0 0 $X=232790 $Y=269760
X4594 VSS 934 SIGN_MEMFLCCMBLST2 $T=233790 274160 1 0 $X=232790 $Y=271460
X4595 VSS 935 SIGN_MEMFLCCMBLST2 $T=233790 274160 0 0 $X=232790 $Y=273160
X4596 VSS 935 SIGN_MEMFLCCMBLST2 $T=233790 277560 1 0 $X=232790 $Y=274860
X4597 VSS 936 SIGN_MEMFLCCMBLST2 $T=233790 277560 0 0 $X=232790 $Y=276560
X4598 VSS 936 SIGN_MEMFLCCMBLST2 $T=233790 280960 1 0 $X=232790 $Y=278260
X4599 VSS 937 SIGN_MEMFLCCMBLST2 $T=233790 280960 0 0 $X=232790 $Y=279960
X4600 VSS 937 SIGN_MEMFLCCMBLST2 $T=233790 284360 1 0 $X=232790 $Y=281660
X4601 VSS 938 SIGN_MEMFLCCMBLST2 $T=233790 284360 0 0 $X=232790 $Y=283360
X4602 VSS 938 SIGN_MEMFLCCMBLST2 $T=233790 287760 1 0 $X=232790 $Y=285060
X4603 VSS 939 SIGN_MEMFLCCMBLST2 $T=233790 287760 0 0 $X=232790 $Y=286760
X4604 VSS 939 SIGN_MEMFLCCMBLST2 $T=233790 291160 1 0 $X=232790 $Y=288460
X4605 VSS 940 SIGN_MEMFLCCMBLST2 $T=233790 291160 0 0 $X=232790 $Y=290160
X4606 VSS 940 SIGN_MEMFLCCMBLST2 $T=233790 294560 1 0 $X=232790 $Y=291860
X4607 VSS 941 SIGN_MEMFLCCMBLST2 $T=233790 294560 0 0 $X=232790 $Y=293560
X4608 VSS 941 SIGN_MEMFLCCMBLST2 $T=233790 297960 1 0 $X=232790 $Y=295260
X4609 VSS 942 SIGN_MEMFLCCMBLST2 $T=233790 297960 0 0 $X=232790 $Y=296960
X4610 VSS 942 SIGN_MEMFLCCMBLST2 $T=233790 301360 1 0 $X=232790 $Y=298660
X4611 VSS 943 SIGN_MEMFLCCMBLST2 $T=233790 301360 0 0 $X=232790 $Y=300360
X4612 VSS 943 SIGN_MEMFLCCMBLST2 $T=233790 304760 1 0 $X=232790 $Y=302060
X4613 VSS 944 SIGN_MEMFLCCMBLST2 $T=233790 304760 0 0 $X=232790 $Y=303760
X4614 VSS 944 SIGN_MEMFLCCMBLST2 $T=233790 308160 1 0 $X=232790 $Y=305460
X4615 VSS 945 SIGN_MEMFLCCMBLST2 $T=233790 308160 0 0 $X=232790 $Y=307160
X4616 VSS 945 SIGN_MEMFLCCMBLST2 $T=233790 311560 1 0 $X=232790 $Y=308860
X4617 VSS 946 SIGN_MEMFLCCMBLST2 $T=233790 311560 0 0 $X=232790 $Y=310560
X4618 VSS 946 SIGN_MEMFLCCMBLST2 $T=233790 314960 1 0 $X=232790 $Y=312260
X4619 VSS 947 SIGN_MEMFLCCMBLST2 $T=233790 314960 0 0 $X=232790 $Y=313960
X4620 VSS 947 SIGN_MEMFLCCMBLST2 $T=233790 318360 1 0 $X=232790 $Y=315660
X4621 VSS 948 SIGN_MEMFLCCMBLST2 $T=233790 318360 0 0 $X=232790 $Y=317360
X4622 VSS 948 SIGN_MEMFLCCMBLST2 $T=233790 321760 1 0 $X=232790 $Y=319060
X4623 VSS 949 SIGN_MEMFLCCMBLST2 $T=233790 321760 0 0 $X=232790 $Y=320760
X4624 VSS 949 SIGN_MEMFLCCMBLST2 $T=233790 325160 1 0 $X=232790 $Y=322460
X4625 VSS 950 SIGN_MEMFLCCMBLST2 $T=233790 325160 0 0 $X=232790 $Y=324160
X4626 VSS 950 SIGN_MEMFLCCMBLST2 $T=233790 328560 1 0 $X=232790 $Y=325860
X4627 VSS 951 SIGN_MEMFLCCMBLST2 $T=233790 328560 0 0 $X=232790 $Y=327560
X4628 VSS 951 SIGN_MEMFLCCMBLST2 $T=233790 331960 1 0 $X=232790 $Y=329260
X4629 VSS 952 SIGN_MEMFLCCMBLST2 $T=233790 331960 0 0 $X=232790 $Y=330960
X4630 VSS 952 SIGN_MEMFLCCMBLST2 $T=233790 335360 1 0 $X=232790 $Y=332660
X4631 VSS 953 SIGN_MEMFLCCMBLST2 $T=233790 335360 0 0 $X=232790 $Y=334360
X4632 VSS 953 SIGN_MEMFLCCMBLST2 $T=233790 338760 1 0 $X=232790 $Y=336060
X4633 VSS 954 SIGN_MEMFLCCMBLST2 $T=233790 338760 0 0 $X=232790 $Y=337760
X4634 VSS 954 SIGN_MEMFLCCMBLST2 $T=233790 342160 1 0 $X=232790 $Y=339460
X4635 VSS 955 SIGN_MEMFLCCMBLST2 $T=233790 342160 0 0 $X=232790 $Y=341160
X4636 VSS 955 SIGN_MEMFLCCMBLST2 $T=233790 345560 1 0 $X=232790 $Y=342860
X4637 VSS 956 SIGN_MEMFLCCMBLST2 $T=233790 345560 0 0 $X=232790 $Y=344560
X4638 VSS 956 SIGN_MEMFLCCMBLST2 $T=233790 348960 1 0 $X=232790 $Y=346260
X4639 VSS 957 SIGN_MEMFLCCMBLST2 $T=233790 348960 0 0 $X=232790 $Y=347960
X4640 VSS 957 SIGN_MEMFLCCMBLST2 $T=233790 352360 1 0 $X=232790 $Y=349660
X4641 VSS 958 SIGN_MEMFLCCMBLST2 $T=233790 352360 0 0 $X=232790 $Y=351360
X4642 VSS 958 SIGN_MEMFLCCMBLST2 $T=233790 355760 1 0 $X=232790 $Y=353060
X4643 VSS 959 SIGN_MEMFLCCMBLST2 $T=233790 355760 0 0 $X=232790 $Y=354760
X4644 VSS 959 SIGN_MEMFLCCMBLST2 $T=233790 359160 1 0 $X=232790 $Y=356460
X4645 VSS 960 SIGN_MEMFLCCMBLST2 $T=233790 359160 0 0 $X=232790 $Y=358160
X4646 VSS 960 SIGN_MEMFLCCMBLST2 $T=233790 362560 1 0 $X=232790 $Y=359860
X4647 VSS 961 SIGN_MEMFLCCMBLST2 $T=233790 362560 0 0 $X=232790 $Y=361560
X4648 VSS 961 SIGN_MEMFLCCMBLST2 $T=233790 365960 1 0 $X=232790 $Y=363260
X4649 VSS 962 SIGN_MEMFLCCMBLST2 $T=233790 365960 0 0 $X=232790 $Y=364960
X4650 VSS 962 SIGN_MEMFLCCMBLST2 $T=233790 369360 1 0 $X=232790 $Y=366660
X4651 VSS 963 SIGN_MEMFLCCMBLST2 $T=233790 369360 0 0 $X=232790 $Y=368360
X4652 VSS 963 SIGN_MEMFLCCMBLST2 $T=233790 372760 1 0 $X=232790 $Y=370060
X4653 VSS 964 SIGN_MEMFLCCMBLST2 $T=233790 372760 0 0 $X=232790 $Y=371760
X4654 VSS 964 SIGN_MEMFLCCMBLST2 $T=233790 376160 1 0 $X=232790 $Y=373460
X4655 VSS 965 SIGN_MEMFLCCMBLST2 $T=233790 376160 0 0 $X=232790 $Y=375160
X4656 VSS 965 SIGN_MEMFLCCMBLST2 $T=233790 379560 1 0 $X=232790 $Y=376860
X4657 VSS 966 SIGN_MEMFLCCMBLST2 $T=233790 379560 0 0 $X=232790 $Y=378560
X4658 VSS 966 SIGN_MEMFLCCMBLST2 $T=233790 382960 1 0 $X=232790 $Y=380260
X4659 VSS 967 SIGN_MEMFLCCMBLST2 $T=233790 382960 0 0 $X=232790 $Y=381960
X4660 VSS 967 SIGN_MEMFLCCMBLST2 $T=233790 386360 1 0 $X=232790 $Y=383660
X4661 VSS 968 SIGN_MEMFLCCMBLST2 $T=233790 386360 0 0 $X=232790 $Y=385360
X4662 VSS 968 SIGN_MEMFLCCMBLST2 $T=233790 389760 1 0 $X=232790 $Y=387060
X4663 VSS 969 SIGN_MEMFLCCMBLST2 $T=233790 389760 0 0 $X=232790 $Y=388760
X4664 VSS 969 SIGN_MEMFLCCMBLST2 $T=233790 393160 1 0 $X=232790 $Y=390460
X4665 VSS 970 SIGN_MEMFLCCMBLST2 $T=233790 393160 0 0 $X=232790 $Y=392160
X4666 VSS 970 SIGN_MEMFLCCMBLST2 $T=233790 396560 1 0 $X=232790 $Y=393860
X4667 VSS 971 SIGN_MEMFLCCMBLST2 $T=233790 396560 0 0 $X=232790 $Y=395560
X4668 VSS 971 SIGN_MEMFLCCMBLST2 $T=233790 399960 1 0 $X=232790 $Y=397260
X4669 VSS 972 SIGN_MEMFLCCMBLST2 $T=233790 399960 0 0 $X=232790 $Y=398960
X4670 VSS 972 SIGN_MEMFLCCMBLST2 $T=233790 403360 1 0 $X=232790 $Y=400660
X4671 VSS 973 SIGN_MEMFLCCMBLST2 $T=233790 403360 0 0 $X=232790 $Y=402360
X4672 VSS 973 SIGN_MEMFLCCMBLST2 $T=233790 406760 1 0 $X=232790 $Y=404060
X4673 VSS 974 SIGN_MEMFLCCMBLST2 $T=233790 406760 0 0 $X=232790 $Y=405760
X4674 VSS 974 SIGN_MEMFLCCMBLST2 $T=233790 410160 1 0 $X=232790 $Y=407460
X4675 VSS 975 SIGN_MEMFLCCMBLST2 $T=233790 410160 0 0 $X=232790 $Y=409160
X4676 VSS 975 SIGN_MEMFLCCMBLST2 $T=233790 413560 1 0 $X=232790 $Y=410860
X4677 VSS 976 SIGN_MEMFLCCMBLST2 $T=233790 413560 0 0 $X=232790 $Y=412560
X4678 VSS 976 SIGN_MEMFLCCMBLST2 $T=233790 416960 1 0 $X=232790 $Y=414260
X4679 VSS 977 SIGN_MEMFLCCMBLST2 $T=233790 416960 0 0 $X=232790 $Y=415960
X4680 VSS 977 SIGN_MEMFLCCMBLST2 $T=233790 420360 1 0 $X=232790 $Y=417660
X4681 VSS 978 SIGN_MEMFLCCMBLST2 $T=233790 420360 0 0 $X=232790 $Y=419360
X4682 VSS 978 SIGN_MEMFLCCMBLST2 $T=233790 423760 1 0 $X=232790 $Y=421060
X4683 VSS 979 SIGN_MEMFLCCMBLST2 $T=233790 423760 0 0 $X=232790 $Y=422760
X4684 VSS 979 SIGN_MEMFLCCMBLST2 $T=233790 427160 1 0 $X=232790 $Y=424460
X4685 VSS 980 SIGN_MEMFLCCMBLST2 $T=233790 427160 0 0 $X=232790 $Y=426160
X4686 VSS 980 SIGN_MEMFLCCMBLST2 $T=233790 430560 1 0 $X=232790 $Y=427860
X4687 VSS 981 SIGN_MEMFLCCMBLST2 $T=233790 430560 0 0 $X=232790 $Y=429560
X4688 VSS 981 SIGN_MEMFLCCMBLST2 $T=233790 433960 1 0 $X=232790 $Y=431260
X4689 VSS 982 SIGN_MEMFLCCMBLST2 $T=233790 433960 0 0 $X=232790 $Y=432960
X4690 VSS 982 SIGN_MEMFLCCMBLST2 $T=233790 437360 1 0 $X=232790 $Y=434660
X4691 VSS 983 SIGN_MEMFLCCMBLST2 $T=233790 437360 0 0 $X=232790 $Y=436360
X4692 VSS 983 SIGN_MEMFLCCMBLST2 $T=233790 440760 1 0 $X=232790 $Y=438060
X4693 VSS 984 SIGN_MEMFLCCMBLST2 $T=233790 440760 0 0 $X=232790 $Y=439760
X4694 VSS 984 SIGN_MEMFLCCMBLST2 $T=233790 444160 1 0 $X=232790 $Y=441460
X4695 VSS 985 SIGN_MEMFLCCMBLST2 $T=233790 444160 0 0 $X=232790 $Y=443160
X4696 VSS 985 SIGN_MEMFLCCMBLST2 $T=233790 447560 1 0 $X=232790 $Y=444860
X4697 VSS 986 SIGN_MEMFLCCMBLST2 $T=233790 447560 0 0 $X=232790 $Y=446560
X4698 VSS 986 SIGN_MEMFLCCMBLST2 $T=233790 450960 1 0 $X=232790 $Y=448260
X4699 VSS 987 SIGN_MEMFLCCMBLST2 $T=233790 450960 0 0 $X=232790 $Y=449960
X4700 VSS 987 SIGN_MEMFLCCMBLST2 $T=233790 454360 1 0 $X=232790 $Y=451660
X4701 VSS 988 SIGN_MEMFLCCMBLST2 $T=233790 454360 0 0 $X=232790 $Y=453360
X4702 VSS 988 SIGN_MEMFLCCMBLST2 $T=233790 457760 1 0 $X=232790 $Y=455060
X4703 VSS 989 SIGN_MEMFLCCMBLST2 $T=233790 457760 0 0 $X=232790 $Y=456760
X4704 VSS 989 SIGN_MEMFLCCMBLST2 $T=233790 461160 1 0 $X=232790 $Y=458460
X4705 VSS 990 SIGN_MEMFLCCMBLST2 $T=233790 461160 0 0 $X=232790 $Y=460160
X4706 VSS 990 SIGN_MEMFLCCMBLST2 $T=233790 464560 1 0 $X=232790 $Y=461860
X4707 VSS 991 SIGN_MEMFLCCMBLST2 $T=233790 464560 0 0 $X=232790 $Y=463560
X4708 VSS 991 SIGN_MEMFLCCMBLST2 $T=233790 467960 1 0 $X=232790 $Y=465260
X4709 VSS 992 SIGN_MEMFLCCMBLST2 $T=233790 467960 0 0 $X=232790 $Y=466960
X4710 VSS 992 SIGN_MEMFLCCMBLST2 $T=233790 471360 1 0 $X=232790 $Y=468660
X4711 VSS 993 SIGN_MEMFLCCMBLST2 $T=233790 471360 0 0 $X=232790 $Y=470360
X4712 VSS 993 SIGN_MEMFLCCMBLST2 $T=233790 474760 1 0 $X=232790 $Y=472060
X4713 VSS 994 SIGN_MEMFLCCMBLST2 $T=233790 474760 0 0 $X=232790 $Y=473760
X4714 VSS 994 SIGN_MEMFLCCMBLST2 $T=233790 478160 1 0 $X=232790 $Y=475460
X4715 VSS 995 SIGN_MEMFLCCMBLST2 $T=233790 478160 0 0 $X=232790 $Y=477160
X4716 VSS 995 SIGN_MEMFLCCMBLST2 $T=233790 481560 1 0 $X=232790 $Y=478860
X4717 VSS 996 SIGN_MEMFLCCMBLST2 $T=233790 481560 0 0 $X=232790 $Y=480560
X4718 VSS 996 SIGN_MEMFLCCMBLST2 $T=233790 484960 1 0 $X=232790 $Y=482260
X4719 VSS 997 SIGN_MEMFLCCMBLST2 $T=233790 484960 0 0 $X=232790 $Y=483960
X4720 VSS 997 SIGN_MEMFLCCMBLST2 $T=233790 488360 1 0 $X=232790 $Y=485660
X4721 VSS 998 SIGN_MEMFLCCMBLST2 $T=233790 488360 0 0 $X=232790 $Y=487360
X4722 VSS 998 SIGN_MEMFLCCMBLST2 $T=233790 491760 1 0 $X=232790 $Y=489060
X4723 VSS 999 SIGN_MEMFLCCMBLST2 $T=233790 491760 0 0 $X=232790 $Y=490760
X4724 VSS 999 SIGN_MEMFLCCMBLST2 $T=233790 495160 1 0 $X=232790 $Y=492460
X4725 VSS 1000 SIGN_MEMFLCCMBLST2 $T=233790 495160 0 0 $X=232790 $Y=494160
X4726 VSS 1000 SIGN_MEMFLCCMBLST2 $T=233790 498560 1 0 $X=232790 $Y=495860
X4727 VSS 1001 SIGN_MEMFLCCMBLST2 $T=233790 498560 0 0 $X=232790 $Y=497560
X4728 VSS 1001 SIGN_MEMFLCCMBLST2 $T=233790 501960 1 0 $X=232790 $Y=499260
X4729 VSS 1002 SIGN_MEMFLCCMBLST2 $T=233790 501960 0 0 $X=232790 $Y=500960
X4730 VSS 1002 SIGN_MEMFLCCMBLST2 $T=233790 505360 1 0 $X=232790 $Y=502660
X4731 VSS 1003 SIGN_MEMFLCCMBLST2 $T=233790 505360 0 0 $X=232790 $Y=504360
X4732 VSS 1003 SIGN_MEMFLCCMBLST2 $T=233790 508760 1 0 $X=232790 $Y=506060
X4733 VSS 63 1004 1005 VSS SIGN_MEMFLCCMBLST $T=236190 73560 0 0 $X=235190 $Y=72560
X4734 VSS 64 1004 1005 VSS SIGN_MEMFLCCMBLST $T=236190 76960 1 0 $X=235190 $Y=74260
X4735 VSS 65 1006 1007 VSS SIGN_MEMFLCCMBLST $T=236190 76960 0 0 $X=235190 $Y=75960
X4736 VSS 66 1006 1007 VSS SIGN_MEMFLCCMBLST $T=236190 80360 1 0 $X=235190 $Y=77660
X4737 VSS 67 1008 1009 VSS SIGN_MEMFLCCMBLST $T=236190 80360 0 0 $X=235190 $Y=79360
X4738 VSS 68 1008 1009 VSS SIGN_MEMFLCCMBLST $T=236190 83760 1 0 $X=235190 $Y=81060
X4739 VSS 69 1010 1011 VSS SIGN_MEMFLCCMBLST $T=236190 83760 0 0 $X=235190 $Y=82760
X4740 VSS 70 1010 1011 VSS SIGN_MEMFLCCMBLST $T=236190 87160 1 0 $X=235190 $Y=84460
X4741 VSS 71 1012 1013 VSS SIGN_MEMFLCCMBLST $T=236190 87160 0 0 $X=235190 $Y=86160
X4742 VSS 72 1012 1013 VSS SIGN_MEMFLCCMBLST $T=236190 90560 1 0 $X=235190 $Y=87860
X4743 VSS 73 1014 1015 VSS SIGN_MEMFLCCMBLST $T=236190 90560 0 0 $X=235190 $Y=89560
X4744 VSS 74 1014 1015 VSS SIGN_MEMFLCCMBLST $T=236190 93960 1 0 $X=235190 $Y=91260
X4745 VSS 75 1016 1017 VSS SIGN_MEMFLCCMBLST $T=236190 93960 0 0 $X=235190 $Y=92960
X4746 VSS 76 1016 1017 VSS SIGN_MEMFLCCMBLST $T=236190 97360 1 0 $X=235190 $Y=94660
X4747 VSS 77 1018 1019 VSS SIGN_MEMFLCCMBLST $T=236190 97360 0 0 $X=235190 $Y=96360
X4748 VSS 78 1018 1019 VSS SIGN_MEMFLCCMBLST $T=236190 100760 1 0 $X=235190 $Y=98060
X4749 VSS 79 1020 1021 VSS SIGN_MEMFLCCMBLST $T=236190 100760 0 0 $X=235190 $Y=99760
X4750 VSS 80 1020 1021 VSS SIGN_MEMFLCCMBLST $T=236190 104160 1 0 $X=235190 $Y=101460
X4751 VSS 81 1022 1023 VSS SIGN_MEMFLCCMBLST $T=236190 104160 0 0 $X=235190 $Y=103160
X4752 VSS 82 1022 1023 VSS SIGN_MEMFLCCMBLST $T=236190 107560 1 0 $X=235190 $Y=104860
X4753 VSS 83 1024 1025 VSS SIGN_MEMFLCCMBLST $T=236190 107560 0 0 $X=235190 $Y=106560
X4754 VSS 84 1024 1025 VSS SIGN_MEMFLCCMBLST $T=236190 110960 1 0 $X=235190 $Y=108260
X4755 VSS 85 1026 1027 VSS SIGN_MEMFLCCMBLST $T=236190 110960 0 0 $X=235190 $Y=109960
X4756 VSS 86 1026 1027 VSS SIGN_MEMFLCCMBLST $T=236190 114360 1 0 $X=235190 $Y=111660
X4757 VSS 87 1028 1029 VSS SIGN_MEMFLCCMBLST $T=236190 114360 0 0 $X=235190 $Y=113360
X4758 VSS 88 1028 1029 VSS SIGN_MEMFLCCMBLST $T=236190 117760 1 0 $X=235190 $Y=115060
X4759 VSS 89 1030 1031 VSS SIGN_MEMFLCCMBLST $T=236190 117760 0 0 $X=235190 $Y=116760
X4760 VSS 90 1030 1031 VSS SIGN_MEMFLCCMBLST $T=236190 121160 1 0 $X=235190 $Y=118460
X4761 VSS 91 1032 1033 VSS SIGN_MEMFLCCMBLST $T=236190 121160 0 0 $X=235190 $Y=120160
X4762 VSS 92 1032 1033 VSS SIGN_MEMFLCCMBLST $T=236190 124560 1 0 $X=235190 $Y=121860
X4763 VSS 93 1034 1035 VSS SIGN_MEMFLCCMBLST $T=236190 124560 0 0 $X=235190 $Y=123560
X4764 VSS 94 1034 1035 VSS SIGN_MEMFLCCMBLST $T=236190 127960 1 0 $X=235190 $Y=125260
X4765 VSS 95 1036 1037 VSS SIGN_MEMFLCCMBLST $T=236190 127960 0 0 $X=235190 $Y=126960
X4766 VSS 96 1036 1037 VSS SIGN_MEMFLCCMBLST $T=236190 131360 1 0 $X=235190 $Y=128660
X4767 VSS 97 1038 1039 VSS SIGN_MEMFLCCMBLST $T=236190 131360 0 0 $X=235190 $Y=130360
X4768 VSS 98 1038 1039 VSS SIGN_MEMFLCCMBLST $T=236190 134760 1 0 $X=235190 $Y=132060
X4769 VSS 99 1040 1041 VSS SIGN_MEMFLCCMBLST $T=236190 134760 0 0 $X=235190 $Y=133760
X4770 VSS 100 1040 1041 VSS SIGN_MEMFLCCMBLST $T=236190 138160 1 0 $X=235190 $Y=135460
X4771 VSS 101 1042 1043 VSS SIGN_MEMFLCCMBLST $T=236190 138160 0 0 $X=235190 $Y=137160
X4772 VSS 102 1042 1043 VSS SIGN_MEMFLCCMBLST $T=236190 141560 1 0 $X=235190 $Y=138860
X4773 VSS 103 1044 1045 VSS SIGN_MEMFLCCMBLST $T=236190 141560 0 0 $X=235190 $Y=140560
X4774 VSS 104 1044 1045 VSS SIGN_MEMFLCCMBLST $T=236190 144960 1 0 $X=235190 $Y=142260
X4775 VSS 105 1046 1047 VSS SIGN_MEMFLCCMBLST $T=236190 144960 0 0 $X=235190 $Y=143960
X4776 VSS 106 1046 1047 VSS SIGN_MEMFLCCMBLST $T=236190 148360 1 0 $X=235190 $Y=145660
X4777 VSS 107 1048 1049 VSS SIGN_MEMFLCCMBLST $T=236190 148360 0 0 $X=235190 $Y=147360
X4778 VSS 108 1048 1049 VSS SIGN_MEMFLCCMBLST $T=236190 151760 1 0 $X=235190 $Y=149060
X4779 VSS 109 1050 1051 VSS SIGN_MEMFLCCMBLST $T=236190 151760 0 0 $X=235190 $Y=150760
X4780 VSS 110 1050 1051 VSS SIGN_MEMFLCCMBLST $T=236190 155160 1 0 $X=235190 $Y=152460
X4781 VSS 111 1052 1053 VSS SIGN_MEMFLCCMBLST $T=236190 155160 0 0 $X=235190 $Y=154160
X4782 VSS 112 1052 1053 VSS SIGN_MEMFLCCMBLST $T=236190 158560 1 0 $X=235190 $Y=155860
X4783 VSS 113 1054 1055 VSS SIGN_MEMFLCCMBLST $T=236190 158560 0 0 $X=235190 $Y=157560
X4784 VSS 114 1054 1055 VSS SIGN_MEMFLCCMBLST $T=236190 161960 1 0 $X=235190 $Y=159260
X4785 VSS 115 1056 1057 VSS SIGN_MEMFLCCMBLST $T=236190 161960 0 0 $X=235190 $Y=160960
X4786 VSS 116 1056 1057 VSS SIGN_MEMFLCCMBLST $T=236190 165360 1 0 $X=235190 $Y=162660
X4787 VSS 117 1058 1059 VSS SIGN_MEMFLCCMBLST $T=236190 165360 0 0 $X=235190 $Y=164360
X4788 VSS 118 1058 1059 VSS SIGN_MEMFLCCMBLST $T=236190 168760 1 0 $X=235190 $Y=166060
X4789 VSS 119 1060 1061 VSS SIGN_MEMFLCCMBLST $T=236190 168760 0 0 $X=235190 $Y=167760
X4790 VSS 120 1060 1061 VSS SIGN_MEMFLCCMBLST $T=236190 172160 1 0 $X=235190 $Y=169460
X4791 VSS 121 1062 1063 VSS SIGN_MEMFLCCMBLST $T=236190 172160 0 0 $X=235190 $Y=171160
X4792 VSS 122 1062 1063 VSS SIGN_MEMFLCCMBLST $T=236190 175560 1 0 $X=235190 $Y=172860
X4793 VSS 123 1064 1065 VSS SIGN_MEMFLCCMBLST $T=236190 175560 0 0 $X=235190 $Y=174560
X4794 VSS 124 1064 1065 VSS SIGN_MEMFLCCMBLST $T=236190 178960 1 0 $X=235190 $Y=176260
X4795 VSS 125 1066 1067 VSS SIGN_MEMFLCCMBLST $T=236190 178960 0 0 $X=235190 $Y=177960
X4796 VSS 126 1066 1067 VSS SIGN_MEMFLCCMBLST $T=236190 182360 1 0 $X=235190 $Y=179660
X4797 VSS 127 1068 1069 VSS SIGN_MEMFLCCMBLST $T=236190 182360 0 0 $X=235190 $Y=181360
X4798 VSS 128 1068 1069 VSS SIGN_MEMFLCCMBLST $T=236190 185760 1 0 $X=235190 $Y=183060
X4799 VSS 129 1070 1071 VSS SIGN_MEMFLCCMBLST $T=236190 185760 0 0 $X=235190 $Y=184760
X4800 VSS 130 1070 1071 VSS SIGN_MEMFLCCMBLST $T=236190 189160 1 0 $X=235190 $Y=186460
X4801 VSS 131 1072 1073 VSS SIGN_MEMFLCCMBLST $T=236190 189160 0 0 $X=235190 $Y=188160
X4802 VSS 132 1072 1073 VSS SIGN_MEMFLCCMBLST $T=236190 192560 1 0 $X=235190 $Y=189860
X4803 VSS 133 1074 1075 VSS SIGN_MEMFLCCMBLST $T=236190 192560 0 0 $X=235190 $Y=191560
X4804 VSS 134 1074 1075 VSS SIGN_MEMFLCCMBLST $T=236190 195960 1 0 $X=235190 $Y=193260
X4805 VSS 135 1076 1077 VSS SIGN_MEMFLCCMBLST $T=236190 195960 0 0 $X=235190 $Y=194960
X4806 VSS 136 1076 1077 VSS SIGN_MEMFLCCMBLST $T=236190 199360 1 0 $X=235190 $Y=196660
X4807 VSS 137 1078 1079 VSS SIGN_MEMFLCCMBLST $T=236190 199360 0 0 $X=235190 $Y=198360
X4808 VSS 138 1078 1079 VSS SIGN_MEMFLCCMBLST $T=236190 202760 1 0 $X=235190 $Y=200060
X4809 VSS 139 1080 1081 VSS SIGN_MEMFLCCMBLST $T=236190 202760 0 0 $X=235190 $Y=201760
X4810 VSS 140 1080 1081 VSS SIGN_MEMFLCCMBLST $T=236190 206160 1 0 $X=235190 $Y=203460
X4811 VSS 141 1082 1083 VSS SIGN_MEMFLCCMBLST $T=236190 206160 0 0 $X=235190 $Y=205160
X4812 VSS 142 1082 1083 VSS SIGN_MEMFLCCMBLST $T=236190 209560 1 0 $X=235190 $Y=206860
X4813 VSS 143 1084 1085 VSS SIGN_MEMFLCCMBLST $T=236190 209560 0 0 $X=235190 $Y=208560
X4814 VSS 144 1084 1085 VSS SIGN_MEMFLCCMBLST $T=236190 212960 1 0 $X=235190 $Y=210260
X4815 VSS 145 1086 1087 VSS SIGN_MEMFLCCMBLST $T=236190 212960 0 0 $X=235190 $Y=211960
X4816 VSS 146 1086 1087 VSS SIGN_MEMFLCCMBLST $T=236190 216360 1 0 $X=235190 $Y=213660
X4817 VSS 147 1088 1089 VSS SIGN_MEMFLCCMBLST $T=236190 216360 0 0 $X=235190 $Y=215360
X4818 VSS 148 1088 1089 VSS SIGN_MEMFLCCMBLST $T=236190 219760 1 0 $X=235190 $Y=217060
X4819 VSS 149 1090 1091 VSS SIGN_MEMFLCCMBLST $T=236190 219760 0 0 $X=235190 $Y=218760
X4820 VSS 150 1090 1091 VSS SIGN_MEMFLCCMBLST $T=236190 223160 1 0 $X=235190 $Y=220460
X4821 VSS 151 1092 1093 VSS SIGN_MEMFLCCMBLST $T=236190 223160 0 0 $X=235190 $Y=222160
X4822 VSS 152 1092 1093 VSS SIGN_MEMFLCCMBLST $T=236190 226560 1 0 $X=235190 $Y=223860
X4823 VSS 153 1094 1095 VSS SIGN_MEMFLCCMBLST $T=236190 226560 0 0 $X=235190 $Y=225560
X4824 VSS 154 1094 1095 VSS SIGN_MEMFLCCMBLST $T=236190 229960 1 0 $X=235190 $Y=227260
X4825 VSS 155 1096 1097 VSS SIGN_MEMFLCCMBLST $T=236190 229960 0 0 $X=235190 $Y=228960
X4826 VSS 156 1096 1097 VSS SIGN_MEMFLCCMBLST $T=236190 233360 1 0 $X=235190 $Y=230660
X4827 VSS 157 1098 1099 VSS SIGN_MEMFLCCMBLST $T=236190 233360 0 0 $X=235190 $Y=232360
X4828 VSS 158 1098 1099 VSS SIGN_MEMFLCCMBLST $T=236190 236760 1 0 $X=235190 $Y=234060
X4829 VSS 159 1100 1101 VSS SIGN_MEMFLCCMBLST $T=236190 236760 0 0 $X=235190 $Y=235760
X4830 VSS 160 1100 1101 VSS SIGN_MEMFLCCMBLST $T=236190 240160 1 0 $X=235190 $Y=237460
X4831 VSS 161 1102 1103 VSS SIGN_MEMFLCCMBLST $T=236190 240160 0 0 $X=235190 $Y=239160
X4832 VSS 162 1102 1103 VSS SIGN_MEMFLCCMBLST $T=236190 243560 1 0 $X=235190 $Y=240860
X4833 VSS 163 1104 1105 VSS SIGN_MEMFLCCMBLST $T=236190 243560 0 0 $X=235190 $Y=242560
X4834 VSS 164 1104 1105 VSS SIGN_MEMFLCCMBLST $T=236190 246960 1 0 $X=235190 $Y=244260
X4835 VSS 165 1106 1107 VSS SIGN_MEMFLCCMBLST $T=236190 246960 0 0 $X=235190 $Y=245960
X4836 VSS 166 1106 1107 VSS SIGN_MEMFLCCMBLST $T=236190 250360 1 0 $X=235190 $Y=247660
X4837 VSS 167 1108 1109 VSS SIGN_MEMFLCCMBLST $T=236190 250360 0 0 $X=235190 $Y=249360
X4838 VSS 168 1108 1109 VSS SIGN_MEMFLCCMBLST $T=236190 253760 1 0 $X=235190 $Y=251060
X4839 VSS 169 1110 1111 VSS SIGN_MEMFLCCMBLST $T=236190 253760 0 0 $X=235190 $Y=252760
X4840 VSS 170 1110 1111 VSS SIGN_MEMFLCCMBLST $T=236190 257160 1 0 $X=235190 $Y=254460
X4841 VSS 171 1112 1113 VSS SIGN_MEMFLCCMBLST $T=236190 257160 0 0 $X=235190 $Y=256160
X4842 VSS 172 1112 1113 VSS SIGN_MEMFLCCMBLST $T=236190 260560 1 0 $X=235190 $Y=257860
X4843 VSS 173 1114 1115 VSS SIGN_MEMFLCCMBLST $T=236190 260560 0 0 $X=235190 $Y=259560
X4844 VSS 174 1114 1115 VSS SIGN_MEMFLCCMBLST $T=236190 263960 1 0 $X=235190 $Y=261260
X4845 VSS 175 1116 1117 VSS SIGN_MEMFLCCMBLST $T=236190 263960 0 0 $X=235190 $Y=262960
X4846 VSS 176 1116 1117 VSS SIGN_MEMFLCCMBLST $T=236190 267360 1 0 $X=235190 $Y=264660
X4847 VSS 177 1118 1119 VSS SIGN_MEMFLCCMBLST $T=236190 267360 0 0 $X=235190 $Y=266360
X4848 VSS 178 1118 1119 VSS SIGN_MEMFLCCMBLST $T=236190 270760 1 0 $X=235190 $Y=268060
X4849 VSS 179 1120 1121 VSS SIGN_MEMFLCCMBLST $T=236190 270760 0 0 $X=235190 $Y=269760
X4850 VSS 180 1120 1121 VSS SIGN_MEMFLCCMBLST $T=236190 274160 1 0 $X=235190 $Y=271460
X4851 VSS 181 1122 1123 VSS SIGN_MEMFLCCMBLST $T=236190 274160 0 0 $X=235190 $Y=273160
X4852 VSS 182 1122 1123 VSS SIGN_MEMFLCCMBLST $T=236190 277560 1 0 $X=235190 $Y=274860
X4853 VSS 183 1124 1125 VSS SIGN_MEMFLCCMBLST $T=236190 277560 0 0 $X=235190 $Y=276560
X4854 VSS 184 1124 1125 VSS SIGN_MEMFLCCMBLST $T=236190 280960 1 0 $X=235190 $Y=278260
X4855 VSS 185 1126 1127 VSS SIGN_MEMFLCCMBLST $T=236190 280960 0 0 $X=235190 $Y=279960
X4856 VSS 186 1126 1127 VSS SIGN_MEMFLCCMBLST $T=236190 284360 1 0 $X=235190 $Y=281660
X4857 VSS 187 1128 1129 VSS SIGN_MEMFLCCMBLST $T=236190 284360 0 0 $X=235190 $Y=283360
X4858 VSS 188 1128 1129 VSS SIGN_MEMFLCCMBLST $T=236190 287760 1 0 $X=235190 $Y=285060
X4859 VSS 189 1130 1131 VSS SIGN_MEMFLCCMBLST $T=236190 287760 0 0 $X=235190 $Y=286760
X4860 VSS 190 1130 1131 VSS SIGN_MEMFLCCMBLST $T=236190 291160 1 0 $X=235190 $Y=288460
X4861 VSS 191 1132 1133 VSS SIGN_MEMFLCCMBLST $T=236190 291160 0 0 $X=235190 $Y=290160
X4862 VSS 192 1132 1133 VSS SIGN_MEMFLCCMBLST $T=236190 294560 1 0 $X=235190 $Y=291860
X4863 VSS 193 1134 1135 VSS SIGN_MEMFLCCMBLST $T=236190 294560 0 0 $X=235190 $Y=293560
X4864 VSS 194 1134 1135 VSS SIGN_MEMFLCCMBLST $T=236190 297960 1 0 $X=235190 $Y=295260
X4865 VSS 195 1136 1137 VSS SIGN_MEMFLCCMBLST $T=236190 297960 0 0 $X=235190 $Y=296960
X4866 VSS 196 1136 1137 VSS SIGN_MEMFLCCMBLST $T=236190 301360 1 0 $X=235190 $Y=298660
X4867 VSS 197 1138 1139 VSS SIGN_MEMFLCCMBLST $T=236190 301360 0 0 $X=235190 $Y=300360
X4868 VSS 198 1138 1139 VSS SIGN_MEMFLCCMBLST $T=236190 304760 1 0 $X=235190 $Y=302060
X4869 VSS 199 1140 1141 VSS SIGN_MEMFLCCMBLST $T=236190 304760 0 0 $X=235190 $Y=303760
X4870 VSS 200 1140 1141 VSS SIGN_MEMFLCCMBLST $T=236190 308160 1 0 $X=235190 $Y=305460
X4871 VSS 201 1142 1143 VSS SIGN_MEMFLCCMBLST $T=236190 308160 0 0 $X=235190 $Y=307160
X4872 VSS 202 1142 1143 VSS SIGN_MEMFLCCMBLST $T=236190 311560 1 0 $X=235190 $Y=308860
X4873 VSS 203 1144 1145 VSS SIGN_MEMFLCCMBLST $T=236190 311560 0 0 $X=235190 $Y=310560
X4874 VSS 204 1144 1145 VSS SIGN_MEMFLCCMBLST $T=236190 314960 1 0 $X=235190 $Y=312260
X4875 VSS 205 1146 1147 VSS SIGN_MEMFLCCMBLST $T=236190 314960 0 0 $X=235190 $Y=313960
X4876 VSS 206 1146 1147 VSS SIGN_MEMFLCCMBLST $T=236190 318360 1 0 $X=235190 $Y=315660
X4877 VSS 207 1148 1149 VSS SIGN_MEMFLCCMBLST $T=236190 318360 0 0 $X=235190 $Y=317360
X4878 VSS 208 1148 1149 VSS SIGN_MEMFLCCMBLST $T=236190 321760 1 0 $X=235190 $Y=319060
X4879 VSS 209 1150 1151 VSS SIGN_MEMFLCCMBLST $T=236190 321760 0 0 $X=235190 $Y=320760
X4880 VSS 210 1150 1151 VSS SIGN_MEMFLCCMBLST $T=236190 325160 1 0 $X=235190 $Y=322460
X4881 VSS 211 1152 1153 VSS SIGN_MEMFLCCMBLST $T=236190 325160 0 0 $X=235190 $Y=324160
X4882 VSS 212 1152 1153 VSS SIGN_MEMFLCCMBLST $T=236190 328560 1 0 $X=235190 $Y=325860
X4883 VSS 213 1154 1155 VSS SIGN_MEMFLCCMBLST $T=236190 328560 0 0 $X=235190 $Y=327560
X4884 VSS 214 1154 1155 VSS SIGN_MEMFLCCMBLST $T=236190 331960 1 0 $X=235190 $Y=329260
X4885 VSS 215 1156 1157 VSS SIGN_MEMFLCCMBLST $T=236190 331960 0 0 $X=235190 $Y=330960
X4886 VSS 216 1156 1157 VSS SIGN_MEMFLCCMBLST $T=236190 335360 1 0 $X=235190 $Y=332660
X4887 VSS 217 1158 1159 VSS SIGN_MEMFLCCMBLST $T=236190 335360 0 0 $X=235190 $Y=334360
X4888 VSS 218 1158 1159 VSS SIGN_MEMFLCCMBLST $T=236190 338760 1 0 $X=235190 $Y=336060
X4889 VSS 219 1160 1161 VSS SIGN_MEMFLCCMBLST $T=236190 338760 0 0 $X=235190 $Y=337760
X4890 VSS 220 1160 1161 VSS SIGN_MEMFLCCMBLST $T=236190 342160 1 0 $X=235190 $Y=339460
X4891 VSS 221 1162 1163 VSS SIGN_MEMFLCCMBLST $T=236190 342160 0 0 $X=235190 $Y=341160
X4892 VSS 222 1162 1163 VSS SIGN_MEMFLCCMBLST $T=236190 345560 1 0 $X=235190 $Y=342860
X4893 VSS 223 1164 1165 VSS SIGN_MEMFLCCMBLST $T=236190 345560 0 0 $X=235190 $Y=344560
X4894 VSS 224 1164 1165 VSS SIGN_MEMFLCCMBLST $T=236190 348960 1 0 $X=235190 $Y=346260
X4895 VSS 225 1166 1167 VSS SIGN_MEMFLCCMBLST $T=236190 348960 0 0 $X=235190 $Y=347960
X4896 VSS 226 1166 1167 VSS SIGN_MEMFLCCMBLST $T=236190 352360 1 0 $X=235190 $Y=349660
X4897 VSS 227 1168 1169 VSS SIGN_MEMFLCCMBLST $T=236190 352360 0 0 $X=235190 $Y=351360
X4898 VSS 228 1168 1169 VSS SIGN_MEMFLCCMBLST $T=236190 355760 1 0 $X=235190 $Y=353060
X4899 VSS 229 1170 1171 VSS SIGN_MEMFLCCMBLST $T=236190 355760 0 0 $X=235190 $Y=354760
X4900 VSS 230 1170 1171 VSS SIGN_MEMFLCCMBLST $T=236190 359160 1 0 $X=235190 $Y=356460
X4901 VSS 231 1172 1173 VSS SIGN_MEMFLCCMBLST $T=236190 359160 0 0 $X=235190 $Y=358160
X4902 VSS 232 1172 1173 VSS SIGN_MEMFLCCMBLST $T=236190 362560 1 0 $X=235190 $Y=359860
X4903 VSS 233 1174 1175 VSS SIGN_MEMFLCCMBLST $T=236190 362560 0 0 $X=235190 $Y=361560
X4904 VSS 234 1174 1175 VSS SIGN_MEMFLCCMBLST $T=236190 365960 1 0 $X=235190 $Y=363260
X4905 VSS 235 1176 1177 VSS SIGN_MEMFLCCMBLST $T=236190 365960 0 0 $X=235190 $Y=364960
X4906 VSS 236 1176 1177 VSS SIGN_MEMFLCCMBLST $T=236190 369360 1 0 $X=235190 $Y=366660
X4907 VSS 237 1178 1179 VSS SIGN_MEMFLCCMBLST $T=236190 369360 0 0 $X=235190 $Y=368360
X4908 VSS 238 1178 1179 VSS SIGN_MEMFLCCMBLST $T=236190 372760 1 0 $X=235190 $Y=370060
X4909 VSS 239 1180 1181 VSS SIGN_MEMFLCCMBLST $T=236190 372760 0 0 $X=235190 $Y=371760
X4910 VSS 240 1180 1181 VSS SIGN_MEMFLCCMBLST $T=236190 376160 1 0 $X=235190 $Y=373460
X4911 VSS 241 1182 1183 VSS SIGN_MEMFLCCMBLST $T=236190 376160 0 0 $X=235190 $Y=375160
X4912 VSS 242 1182 1183 VSS SIGN_MEMFLCCMBLST $T=236190 379560 1 0 $X=235190 $Y=376860
X4913 VSS 243 1184 1185 VSS SIGN_MEMFLCCMBLST $T=236190 379560 0 0 $X=235190 $Y=378560
X4914 VSS 244 1184 1185 VSS SIGN_MEMFLCCMBLST $T=236190 382960 1 0 $X=235190 $Y=380260
X4915 VSS 245 1186 1187 VSS SIGN_MEMFLCCMBLST $T=236190 382960 0 0 $X=235190 $Y=381960
X4916 VSS 246 1186 1187 VSS SIGN_MEMFLCCMBLST $T=236190 386360 1 0 $X=235190 $Y=383660
X4917 VSS 247 1188 1189 VSS SIGN_MEMFLCCMBLST $T=236190 386360 0 0 $X=235190 $Y=385360
X4918 VSS 248 1188 1189 VSS SIGN_MEMFLCCMBLST $T=236190 389760 1 0 $X=235190 $Y=387060
X4919 VSS 249 1190 1191 VSS SIGN_MEMFLCCMBLST $T=236190 389760 0 0 $X=235190 $Y=388760
X4920 VSS 250 1190 1191 VSS SIGN_MEMFLCCMBLST $T=236190 393160 1 0 $X=235190 $Y=390460
X4921 VSS 251 1192 1193 VSS SIGN_MEMFLCCMBLST $T=236190 393160 0 0 $X=235190 $Y=392160
X4922 VSS 252 1192 1193 VSS SIGN_MEMFLCCMBLST $T=236190 396560 1 0 $X=235190 $Y=393860
X4923 VSS 253 1194 1195 VSS SIGN_MEMFLCCMBLST $T=236190 396560 0 0 $X=235190 $Y=395560
X4924 VSS 254 1194 1195 VSS SIGN_MEMFLCCMBLST $T=236190 399960 1 0 $X=235190 $Y=397260
X4925 VSS 255 1196 1197 VSS SIGN_MEMFLCCMBLST $T=236190 399960 0 0 $X=235190 $Y=398960
X4926 VSS 256 1196 1197 VSS SIGN_MEMFLCCMBLST $T=236190 403360 1 0 $X=235190 $Y=400660
X4927 VSS 257 1198 1199 VSS SIGN_MEMFLCCMBLST $T=236190 403360 0 0 $X=235190 $Y=402360
X4928 VSS 258 1198 1199 VSS SIGN_MEMFLCCMBLST $T=236190 406760 1 0 $X=235190 $Y=404060
X4929 VSS 259 1200 1201 VSS SIGN_MEMFLCCMBLST $T=236190 406760 0 0 $X=235190 $Y=405760
X4930 VSS 260 1200 1201 VSS SIGN_MEMFLCCMBLST $T=236190 410160 1 0 $X=235190 $Y=407460
X4931 VSS 261 1202 1203 VSS SIGN_MEMFLCCMBLST $T=236190 410160 0 0 $X=235190 $Y=409160
X4932 VSS 262 1202 1203 VSS SIGN_MEMFLCCMBLST $T=236190 413560 1 0 $X=235190 $Y=410860
X4933 VSS 263 1204 1205 VSS SIGN_MEMFLCCMBLST $T=236190 413560 0 0 $X=235190 $Y=412560
X4934 VSS 264 1204 1205 VSS SIGN_MEMFLCCMBLST $T=236190 416960 1 0 $X=235190 $Y=414260
X4935 VSS 265 1206 1207 VSS SIGN_MEMFLCCMBLST $T=236190 416960 0 0 $X=235190 $Y=415960
X4936 VSS 266 1206 1207 VSS SIGN_MEMFLCCMBLST $T=236190 420360 1 0 $X=235190 $Y=417660
X4937 VSS 267 1208 1209 VSS SIGN_MEMFLCCMBLST $T=236190 420360 0 0 $X=235190 $Y=419360
X4938 VSS 268 1208 1209 VSS SIGN_MEMFLCCMBLST $T=236190 423760 1 0 $X=235190 $Y=421060
X4939 VSS 269 1210 1211 VSS SIGN_MEMFLCCMBLST $T=236190 423760 0 0 $X=235190 $Y=422760
X4940 VSS 270 1210 1211 VSS SIGN_MEMFLCCMBLST $T=236190 427160 1 0 $X=235190 $Y=424460
X4941 VSS 271 1212 1213 VSS SIGN_MEMFLCCMBLST $T=236190 427160 0 0 $X=235190 $Y=426160
X4942 VSS 272 1212 1213 VSS SIGN_MEMFLCCMBLST $T=236190 430560 1 0 $X=235190 $Y=427860
X4943 VSS 273 1214 1215 VSS SIGN_MEMFLCCMBLST $T=236190 430560 0 0 $X=235190 $Y=429560
X4944 VSS 274 1214 1215 VSS SIGN_MEMFLCCMBLST $T=236190 433960 1 0 $X=235190 $Y=431260
X4945 VSS 275 1216 1217 VSS SIGN_MEMFLCCMBLST $T=236190 433960 0 0 $X=235190 $Y=432960
X4946 VSS 276 1216 1217 VSS SIGN_MEMFLCCMBLST $T=236190 437360 1 0 $X=235190 $Y=434660
X4947 VSS 277 1218 1219 VSS SIGN_MEMFLCCMBLST $T=236190 437360 0 0 $X=235190 $Y=436360
X4948 VSS 278 1218 1219 VSS SIGN_MEMFLCCMBLST $T=236190 440760 1 0 $X=235190 $Y=438060
X4949 VSS 279 1220 1221 VSS SIGN_MEMFLCCMBLST $T=236190 440760 0 0 $X=235190 $Y=439760
X4950 VSS 280 1220 1221 VSS SIGN_MEMFLCCMBLST $T=236190 444160 1 0 $X=235190 $Y=441460
X4951 VSS 281 1222 1223 VSS SIGN_MEMFLCCMBLST $T=236190 444160 0 0 $X=235190 $Y=443160
X4952 VSS 282 1222 1223 VSS SIGN_MEMFLCCMBLST $T=236190 447560 1 0 $X=235190 $Y=444860
X4953 VSS 283 1224 1225 VSS SIGN_MEMFLCCMBLST $T=236190 447560 0 0 $X=235190 $Y=446560
X4954 VSS 284 1224 1225 VSS SIGN_MEMFLCCMBLST $T=236190 450960 1 0 $X=235190 $Y=448260
X4955 VSS 285 1226 1227 VSS SIGN_MEMFLCCMBLST $T=236190 450960 0 0 $X=235190 $Y=449960
X4956 VSS 286 1226 1227 VSS SIGN_MEMFLCCMBLST $T=236190 454360 1 0 $X=235190 $Y=451660
X4957 VSS 287 1228 1229 VSS SIGN_MEMFLCCMBLST $T=236190 454360 0 0 $X=235190 $Y=453360
X4958 VSS 288 1228 1229 VSS SIGN_MEMFLCCMBLST $T=236190 457760 1 0 $X=235190 $Y=455060
X4959 VSS 289 1230 1231 VSS SIGN_MEMFLCCMBLST $T=236190 457760 0 0 $X=235190 $Y=456760
X4960 VSS 290 1230 1231 VSS SIGN_MEMFLCCMBLST $T=236190 461160 1 0 $X=235190 $Y=458460
X4961 VSS 291 1232 1233 VSS SIGN_MEMFLCCMBLST $T=236190 461160 0 0 $X=235190 $Y=460160
X4962 VSS 292 1232 1233 VSS SIGN_MEMFLCCMBLST $T=236190 464560 1 0 $X=235190 $Y=461860
X4963 VSS 293 1234 1235 VSS SIGN_MEMFLCCMBLST $T=236190 464560 0 0 $X=235190 $Y=463560
X4964 VSS 294 1234 1235 VSS SIGN_MEMFLCCMBLST $T=236190 467960 1 0 $X=235190 $Y=465260
X4965 VSS 295 1236 1237 VSS SIGN_MEMFLCCMBLST $T=236190 467960 0 0 $X=235190 $Y=466960
X4966 VSS 296 1236 1237 VSS SIGN_MEMFLCCMBLST $T=236190 471360 1 0 $X=235190 $Y=468660
X4967 VSS 297 1238 1239 VSS SIGN_MEMFLCCMBLST $T=236190 471360 0 0 $X=235190 $Y=470360
X4968 VSS 298 1238 1239 VSS SIGN_MEMFLCCMBLST $T=236190 474760 1 0 $X=235190 $Y=472060
X4969 VSS 299 1240 1241 VSS SIGN_MEMFLCCMBLST $T=236190 474760 0 0 $X=235190 $Y=473760
X4970 VSS 300 1240 1241 VSS SIGN_MEMFLCCMBLST $T=236190 478160 1 0 $X=235190 $Y=475460
X4971 VSS 301 1242 1243 VSS SIGN_MEMFLCCMBLST $T=236190 478160 0 0 $X=235190 $Y=477160
X4972 VSS 302 1242 1243 VSS SIGN_MEMFLCCMBLST $T=236190 481560 1 0 $X=235190 $Y=478860
X4973 VSS 303 1244 1245 VSS SIGN_MEMFLCCMBLST $T=236190 481560 0 0 $X=235190 $Y=480560
X4974 VSS 304 1244 1245 VSS SIGN_MEMFLCCMBLST $T=236190 484960 1 0 $X=235190 $Y=482260
X4975 VSS 305 1246 1247 VSS SIGN_MEMFLCCMBLST $T=236190 484960 0 0 $X=235190 $Y=483960
X4976 VSS 306 1246 1247 VSS SIGN_MEMFLCCMBLST $T=236190 488360 1 0 $X=235190 $Y=485660
X4977 VSS 307 1248 1249 VSS SIGN_MEMFLCCMBLST $T=236190 488360 0 0 $X=235190 $Y=487360
X4978 VSS 308 1248 1249 VSS SIGN_MEMFLCCMBLST $T=236190 491760 1 0 $X=235190 $Y=489060
X4979 VSS 309 1250 1251 VSS SIGN_MEMFLCCMBLST $T=236190 491760 0 0 $X=235190 $Y=490760
X4980 VSS 310 1250 1251 VSS SIGN_MEMFLCCMBLST $T=236190 495160 1 0 $X=235190 $Y=492460
X4981 VSS 311 1252 1253 VSS SIGN_MEMFLCCMBLST $T=236190 495160 0 0 $X=235190 $Y=494160
X4982 VSS 312 1252 1253 VSS SIGN_MEMFLCCMBLST $T=236190 498560 1 0 $X=235190 $Y=495860
X4983 VSS 313 1254 1255 VSS SIGN_MEMFLCCMBLST $T=236190 498560 0 0 $X=235190 $Y=497560
X4984 VSS 314 1254 1255 VSS SIGN_MEMFLCCMBLST $T=236190 501960 1 0 $X=235190 $Y=499260
X4985 VSS 315 1256 1257 VSS SIGN_MEMFLCCMBLST $T=236190 501960 0 0 $X=235190 $Y=500960
X4986 VSS 316 1256 1257 VSS SIGN_MEMFLCCMBLST $T=236190 505360 1 0 $X=235190 $Y=502660
X4987 VSS 317 1258 1259 VSS SIGN_MEMFLCCMBLST $T=236190 505360 0 0 $X=235190 $Y=504360
X4988 VSS 318 1258 1259 VSS SIGN_MEMFLCCMBLST $T=236190 508760 1 0 $X=235190 $Y=506060
X4989 VSS 50 1260 SIGN_MEMFLCCMBLSTU $T=236190 509800 0 0 $X=235190 $Y=508800
X4990 VSS 50 1260 SIGN_MEMFLCCMBLSTU $T=236190 513200 1 0 $X=235190 $Y=510500
X4991 VSS VDD D<8> Q<8> D<9> Q<9> D<10> Q<10> D<11> Q<11> D<12> Q<12> D<13> Q<13> D<14> Q<14> D<15> Q<15> 63 64
+ 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84
+ 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264
+ 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284
+ 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304
+ 305 306 307 308 309 310 311 312 313 314 315 316 317 318 324 325 326 327 328 329
+ 330 331 332 333 51 323 51 VSS 51 5375 5376 5377 5378 5379 5380 5381 5382 5383 5384 5385
+ 5386 5387 5388 5389 5390 5391 5392 5393 5394 5395 5396 5397 5398 5399 5400 5401 5402 5403 5404 5405
+ 5406 5407 5408 5409 5410 5411 5412 5413 5414 5415 5416 5417 5418 5419 5420 5421 5422 5423 5424 5425
+ 5426 5427 5428 5429 5430 5431 5432 5433 5434 5435 5436 5437 5438 5439 5440 5441 5442 5443 5444 5445
+ 5446 5447 5448 5449 5450 5451 5452 5453 5454 5455 5456 5457 5458 5459 5460 5461 5462 5463 5464 5465
+ 5466 5467 5468 5469 5470 5471 5472 5473 5474 5475 5476 5477 5478 5479 5480 5481 5482 5483 5484 5485
+ 5486 5487 5488 5489 5490 5491 5492 5493 5494 5495 5496 5497 5498 5499 5500 5501 5502 5503 5504 5505
+ 5506 5507 5508 5509 5510 5511 5512 5513 5514 5515 5516 5517 5518 5519 5520 5521 5522 5523 5524 5525
+ 5526 5527 5528 5529 5530 5531 5532 5533 5534 5535 5536 5537 5538 5539 5540 5541 5542 5543 5544 5545
+ 5546 5547 5548 5549 5550 5551 5552 5553 5554 5555 5556 5557 5558 5559 5560 5561 5562 5563 5564 5565
+ 5566 5567 5568 5569 5570 5571 5572 5573 5574 5575 5576 5577 5578 5579 5580 5581 5582 5583 5584 5585
+ 5586 5587 5588 5589 5590 5591 5592 5593 5594 5595 5596 5597 5598 5599 5600 5601 5602 5603 5604 5605
+ 5606 5607 5608 5609 5610 5611 5612 5613 5614 5615 5616 5617 5618 5619 5620 5621 5622 5623 5624 5625
+ 5626 5627 5628 5629 5630 5631 5632 5633 5634 5635 5636 5637 5638 5639 5640 5641 5642 5643 5644 5645
+ 5646 5647 5648 5649 5650 5651 5652 5653 5654 5655 5656 5657 5658 5659 5660 5661 5662 5663 5664 5665
+ 5666 5667 5668 5669 5670 5671 5672 5673 5674 5675 5676 5677 5678 5679 5680 5681 5682 5683 5684 5685
+ 5686 5687 5688 5689 5690 5691 5692 5693 5694 5695 5696 5697 5698 5699 5700 5701 5702 5703 5704 5705
+ 5706 5707 5708 5709 5710 5711 5712 5713 5714 5715 5716 5717 5718 5719 5720 5721 5722 5723 5724 5725
+ 5726 5727 5728 5729 5730 5731 5732 5733 5734 5735 5736 5737 5738 5739 5740 5741 5742 5743 5744 5745
+ 5746 5747 5748 5749 5750 5751 5752 5753 5754 5755 5756 5757 5758 5759 5760 5761 5762 5763 5764 5765
+ 5766 5767 5768 5769 5770 5771 5772 5773 5774 5775 5776 5777 5778 5779 5780 5781 5782 5783 5784 5785
+ 5786 5787 5788 5789 5790 5791 5792 5793 5794 5795 5796 5797 5798 5799 5800 5801 5802 5803 5804 5805
+ 5806 5807 5808 5809 5810 5811 5812 5813 5814 5815 5816 5817 5818 5819 5820 5821 5822 5823 5824 5825
+ 5826 5827 5828 5829 5830 5831 5832 5833 5834 5835 5836 5837 5838 5839 5840 5841 5842 5843 5844 5845
+ 5846 5847 5848 5849 5850 5851 5852 5853 5854 5855 5856 5857 5858 5859 5860 5861 5862 5863 5864 5865
+ 5866 5867 5868 5869 5870 5871 5872 5873 5874 5875 5876 5877 5878 5879 5880 5881 5882 5883 5884 5885
+ 5886 5887 5888
+ SIGN_MEMWING_8_RIGHT $T=237390 10240 0 0 $X=236390 $Y=9240
X4992 VDD VSS 5889 5890 base_flme_nvpv $T=316590 509800 0 0 $X=315590 $Y=508800
X4993 VDD VSS 5891 5892 base_flme_nvpv $T=317790 513200 0 180 $X=315590 $Y=510500
.ENDS
***************************************
.SUBCKT ICV_143 1 2 327 831 832 833 849 852 854 881 882 885 887 915 916 917 919 939 941 942
+ 943 954 955 960 962 965 972 974 976 979 982 985 988 996 1019 1020 1022 1024 1048 1050
+ 1052 1054 1082 1085 1088 1111 1113 1115 1117
** N=37952 EP=49 IP=49 FDC=420541
X0 1 2 943 942 941 939 919 917 916 915 887 885 882 881 854 852 831 849 954 955
+ 960 962 965 972 974 976 979 982 985 988 832 996 327 1019 1020 1022 1024 1048 1050 1052
+ 1054 1082 1085 833 1088 1111 1113 1115 1117
+ SIGN_MEM $T=0 0 0 0 $X=-2 $Y=-2
.ENDS
***************************************
.SUBCKT ICV_147 1 2 3 4
** N=4 EP=4 IP=4 FDC=0
X0 1 2 3 4 PDVSS $T=0 0 0 0 $X=-140 $Y=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_175
** N=5 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_174 1 2 3 4
** N=1584 EP=4 IP=60 FDC=220
X13 2 3 4 1 PVDD $T=2000000 255000 0 90 $X=1753000 $Y=254860
X14 2 3 4 1 PVSS $T=2000000 330000 0 90 $X=1753000 $Y=329860
.ENDS
***************************************
.SUBCKT ICV_157 1 2 3 4 21 22 23 24 25 26
** N=1643 EP=10 IP=69 FDC=807
X4 3 2 4 1 1 22 21 PICS $T=2000000 405000 0 90 $X=1752998 $Y=404750
X5 3 2 4 1 1 24 23 PICS $T=2000000 480000 0 90 $X=1752998 $Y=479750
X6 3 2 4 1 1 26 25 PICS $T=2000000 555000 0 90 $X=1752998 $Y=554750
.ENDS
***************************************
.SUBCKT ICV_156 1 2 5 6 46 53 56 57 58 59 60 61 62 63 64 65 66 67
** N=2104 EP=18 IP=133 FDC=1883
X7 5 1 6 2 2 53 57 PICS $T=705000 -2000000 0 0 $X=704750 $Y=-2000000
X8 5 1 6 2 2 46 58 PICS $T=780000 -2000000 0 0 $X=779750 $Y=-2000000
X9 5 1 6 2 2 60 59 PICS $T=855000 -2000000 0 0 $X=854750 $Y=-2000000
X10 5 1 6 2 2 62 61 PICS $T=930000 -2000000 0 0 $X=929750 $Y=-2000000
X11 5 1 6 2 2 64 63 PICS $T=1005000 -2000000 0 0 $X=1004750 $Y=-2000000
X12 5 1 6 2 2 66 65 PICS $T=1080000 -2000000 0 0 $X=1079750 $Y=-2000000
X13 5 1 6 2 2 56 67 PICS $T=1155000 -2000000 0 0 $X=1154750 $Y=-2000000
.ENDS
***************************************
.SUBCKT ICV_155 1 2 5 6 27 28 29 30
** N=844 EP=8 IP=74 FDC=538
X15 5 2 6 1 1 28 27 PICS $T=2000000 1230000 0 90 $X=1752998 $Y=1229750
X16 5 2 6 1 1 30 29 PICS $T=2000000 1305000 0 90 $X=1752998 $Y=1304750
.ENDS
***************************************
.SUBCKT ICV_154 1 2 5 6 45 46 47 48
** N=1169 EP=8 IP=66 FDC=758
X4 2 5 6 1 PDVDD $T=2000000 1605000 0 90 $X=1753000 $Y=1604860
X5 5 2 6 1 1 46 45 PICS $T=2000000 1455000 0 90 $X=1752998 $Y=1454750
X6 5 2 6 1 1 48 47 PICS $T=2000000 1530000 0 90 $X=1752998 $Y=1529750
.ENDS
***************************************
.SUBCKT ICV_149
** N=125 EP=0 IP=40 FDC=0
.ENDS
***************************************
.SUBCKT ICV_146
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_144 1 2 3 4 5 6
** N=6 EP=6 IP=7 FDC=269
X0 2 1 3 4 4 6 5 PICS $T=0 0 0 0 $X=-250 $Y=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6
** N=6 EP=6 IP=7 FDC=269
X0 2 1 3 4 4 6 5 PICS $T=0 0 0 0 $X=-250 $Y=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4
** N=4 EP=4 IP=4 FDC=0
X0 1 2 3 4 PDVSS $T=0 0 0 0 $X=-140 $Y=0
.ENDS
***************************************
.SUBCKT mult_chip VSS DVSS DVDD VDD i_clk i_reset o_smem_rdata<0> o_smem_rdata<1> o_smem_rdata<2> o_smem_rdata<3> o_smem_rdata<4> o_smem_rdata<5> o_smem_rdata<6> o_smem_rdata<7> o_smem_rdata<8> o_smem_rdata<9> o_smem_rdata<10> o_smem_rdata<11> o_smem_rdata<12> o_smem_rdata<13>
+ o_smem_rdata<14> o_smem_rdata<15> i_smem_ext i_smem_cen i_smem_wen i_smem_addr<0> i_smem_addr<1> i_smem_addr<2> i_smem_addr<3> i_smem_addr<4> i_smem_addr<5> i_smem_addr<6> i_smem_addr<7> i_smem_addr<8> i_smem_addr<9> i_smem_addr<10> i_smem_addr<11> i_smem_wdata<0> i_smem_wdata<1> i_smem_wdata<2>
+ i_smem_wdata<4> i_smem_wdata<5> i_smem_wdata<6> i_smem_wdata<7> i_smem_wdata<8> i_smem_wdata<9> i_smem_wdata<10> i_smem_wdata<11> i_smem_wdata<12> i_smem_wdata<14> i_smem_wdata<15> i_smem_wdata<3> i_smem_wdata<13>
** N=8050 EP=53 IP=16320 FDC=445052
X4 VSS DVSS DVDD VDD i_clk 4985 i_reset 932 ICV_260 $T=0 0 0 90 $X=0 $Y=687400
X11 VSS DVSS DVDD VDD o_smem_rdata<0> o_smem_rdata<1> o_smem_rdata<2> o_smem_rdata<3> o_smem_rdata<4> o_smem_rdata<5> o_smem_rdata<6> o_smem_rdata<7> o_smem_rdata<8> o_smem_rdata<9> o_smem_rdata<10> o_smem_rdata<11> o_smem_rdata<12> o_smem_rdata<13> o_smem_rdata<14> o_smem_rdata<15>
+ 5410 5411 5412 5413 5414 5415 5416 5417 5418 5419 5420 5421 5422 5423 5424 5425
+ ICV_256 $T=0 0 0 0 $X=246860 $Y=-2
X12 VSS VDD DVSS DVDD i_smem_ext 5469 i_smem_cen 5495 i_smem_wen 5480 i_smem_addr<0> 5506 i_smem_addr<1> 5515 i_smem_addr<2> 5520 i_smem_addr<3> 4047 i_smem_addr<4> 5539
+ i_smem_addr<5> 5559 i_smem_addr<6> 5594 i_smem_addr<7> 5616 i_smem_addr<8> 5701 i_smem_addr<9> 5682 i_smem_addr<10> 5700 i_smem_addr<11> 5735
+ ICV_179 $T=0 0 0 0 $X=246860 $Y=1735700
X14 VSS VDD 6521 6518 ICV_239 $T=0 0 0 0 $X=247000 $Y=399400
X15 VSS VDD 5224 4047 6981 1757 4264 6972 6961 6959 6872 3970 5227 5217 5230 5223 6886 5229 5216 6848
+ 6873 6885 6887 6888 2196 6897 6898 6900 6852 6906 6915 6909 6914 6916 6984 6917 6918 6919 6983 6931
+ 6930 6945 6948 5235 6975 7058 4985 6706 5233 6858 5215 5225 5219 5220 3971 5506 6859 6518 6874 6845
+ 6905 6913 6910 5234 6982 6922 6933 6844 6990 6993 7078 5713 7076 7077 7085 7030 4980 5469 6707 6754
+ 6755 5228 5221 5226 5218 6763 5515 5520 5222 5414 5415 6839 6840 6847 6849 6850 6857 6871 5417 6899
+ 6911 6932 6946 6960 6973 5424 5704 6989 6987 6974 6985 6988 6986 6991 5425 5708 5735 5243 6629 5410
+ 5411 5412 5413 5416 5418 5419 5420 5421 6947 5422 5423 6992 5398 5323 5766
+ ICV_235 $T=0 0 0 0 $X=247000 $Y=687400
X16 VSS VDD 3971 3970 6763 6850 6849 6987 6988 6993 4264 6839 6840 6848 5594 7739 5700 5701 6986 6985
+ 5682 5753 5539 6852 5559 6982 6983 6984 5752 6521 7030 7740 5334 1984 5335 5243 6845
+ ICV_210 $T=0 0 0 0 $X=247000 $Y=1220200
X17 VSS VDD 932 5616 4983 5093 1986 4982 5480 6989 5708 6991 6992 5753 7058 5704 7076 7077 7739 7078
+ 7085 5752 5323 5723 4981 5397 1985 5090 6629 6754 5495 6755 6847 5092 6990 1983 5713 5091 5094 5095
+ 5766 7740 5096
+ ICV_202 $T=0 0 0 0 $X=247000 $Y=1436200
X18 VDD VSS 6706 5215 5220 5221 5223 5224 5225 5229 5216 6707 5218 5222 5217 5219 5226 5227 5228 5230 ICV_1 $T=500000 925000 0 0 $X=500000 $Y=924900
X19 VDD VSS 1757 5233 5234 5235 6857 6858 6859 6871 6872 6873 6874 6885 6886 6887 6888 6897 6898 6899
+ 6900 6905 6906 6909 6910 6911 6913 6914 6915 6916 6917 6918 6919 6922 6930 6931 6932 6933 6945 6946
+ 6947 6948 6959 6960 6961 6972 6973 6974 6975
+ ICV_143 $T=1000000 750000 0 0 $X=999998 $Y=749998
X20 VSS DVSS DVDD VDD ICV_147 $T=1680000 0 0 0 $X=1679860 $Y=0
X23 VDD VSS DVSS DVDD ICV_174 $T=0 0 0 0 $X=1737400 $Y=246860
X24 VDD VSS DVSS DVDD i_smem_wdata<0> 5398 i_smem_wdata<1> 1984 i_smem_wdata<2> 4980 ICV_157 $T=0 0 0 0 $X=1737400 $Y=399860
X25 VSS VDD DVSS DVDD 4982 5335 5094 i_smem_wdata<4> i_smem_wdata<5> i_smem_wdata<6> 5397 i_smem_wdata<7> 5095 i_smem_wdata<8> 5096 i_smem_wdata<9> 5093 i_smem_wdata<10> ICV_156 $T=0 0 0 90 $X=1737400 $Y=687400
X26 VDD VSS DVSS DVDD i_smem_wdata<11> 5091 i_smem_wdata<12> 4983 ICV_155 $T=0 0 0 0 $X=1737400 $Y=1220200
X27 VDD VSS DVSS DVDD i_smem_wdata<14> 1986 i_smem_wdata<15> 5092 ICV_154 $T=0 0 0 0 $X=1737400 $Y=1437000
X31 VSS DVSS DVDD VDD i_smem_wdata<3> 4981 ICV_144 $T=2000000 630000 0 90 $X=1752998 $Y=629750
X32 VSS DVSS DVDD VDD i_smem_wdata<13> 1983 ICV_41 $T=2000000 1380000 0 90 $X=1752998 $Y=1379750
X33 VSS DVSS DVDD VDD ICV_27 $T=2000000 1680000 0 90 $X=1753000 $Y=1679860
.ENDS
***************************************
