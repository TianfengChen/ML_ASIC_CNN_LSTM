SITE IBM13SITE
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.400 BY 3.600 ;
END IBM13SITE

MACRO XOR3XLTR
    CLASS CORE ;
    FOREIGN XOR3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.030 7.520 3.160 ;
        RECT  7.280 2.040 7.290 3.160 ;
        END
        ANTENNADIFFAREA 1.202 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.480 2.350 6.720 2.830 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.300 1.640 4.460 2.360 ;
        RECT  4.200 1.640 4.300 1.960 ;
        RECT  4.040 1.180 4.200 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.440 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.070 -0.280 7.600 0.280 ;
        RECT  6.780 -0.280 7.070 0.340 ;
        RECT  1.840 -0.280 6.780 0.280 ;
        RECT  1.560 -0.280 1.840 0.610 ;
        RECT  0.360 -0.280 1.560 0.280 ;
        RECT  0.090 -0.280 0.360 0.770 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.040 3.320 7.600 3.880 ;
        RECT  6.880 1.970 7.040 3.880 ;
        RECT  6.710 1.970 6.880 2.130 ;
        RECT  2.300 3.320 6.880 3.880 ;
        RECT  2.020 2.930 2.300 3.880 ;
        RECT  0.380 3.320 2.020 3.880 ;
        RECT  0.120 3.190 0.380 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.970 0.540 7.130 1.750 ;
        RECT  5.430 0.540 6.970 0.700 ;
        RECT  6.330 0.910 6.490 2.190 ;
        RECT  6.290 0.910 6.330 1.620 ;
        RECT  6.060 1.460 6.290 1.620 ;
        RECT  5.900 0.890 6.120 1.050 ;
        RECT  6.110 2.450 6.120 3.090 ;
        RECT  5.950 1.800 6.110 3.090 ;
        RECT  5.900 1.800 5.950 1.960 ;
        RECT  2.620 2.930 5.950 3.090 ;
        RECT  5.740 0.890 5.900 1.960 ;
        RECT  5.430 2.550 5.700 2.710 ;
        RECT  5.270 0.540 5.430 2.710 ;
        RECT  4.940 0.830 5.100 2.770 ;
        RECT  4.890 0.830 4.940 1.110 ;
        RECT  4.710 0.450 4.890 1.110 ;
        RECT  4.620 1.320 4.780 2.710 ;
        RECT  3.880 0.450 4.710 0.610 ;
        RECT  4.530 1.320 4.620 1.480 ;
        RECT  3.240 2.550 4.620 2.710 ;
        RECT  4.370 0.840 4.530 1.480 ;
        RECT  4.090 0.840 4.370 1.000 ;
        RECT  3.880 2.120 4.040 2.360 ;
        RECT  3.720 0.450 3.880 2.360 ;
        RECT  3.400 0.450 3.560 2.360 ;
        RECT  2.160 0.450 3.400 0.610 ;
        RECT  3.080 0.770 3.240 2.710 ;
        RECT  2.480 0.770 3.080 0.930 ;
        RECT  2.640 1.090 2.920 2.450 ;
        RECT  1.400 2.290 2.640 2.450 ;
        RECT  2.460 2.610 2.620 3.090 ;
        RECT  2.320 0.770 2.480 2.130 ;
        RECT  1.080 2.610 2.460 2.770 ;
        RECT  1.720 1.970 2.320 2.130 ;
        RECT  2.000 0.450 2.160 1.790 ;
        RECT  0.850 0.770 2.000 0.930 ;
        RECT  1.900 1.510 2.000 1.790 ;
        RECT  1.720 1.090 1.840 1.310 ;
        RECT  1.560 1.090 1.720 2.130 ;
        RECT  1.240 1.960 1.400 2.450 ;
        RECT  1.080 1.090 1.320 1.250 ;
        RECT  0.920 1.090 1.080 2.770 ;
        RECT  0.760 0.510 0.850 0.930 ;
        RECT  0.600 0.510 0.760 2.830 ;
    END
END XOR3XLTR

MACRO XOR3X4TR
    CLASS CORE ;
    FOREIGN XOR3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.320 1.280 10.420 2.280 ;
        RECT  10.220 0.440 10.320 2.280 ;
        RECT  10.180 0.440 10.220 3.160 ;
        RECT  9.910 0.440 10.180 1.440 ;
        RECT  9.940 2.040 10.180 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.460 1.240 9.560 1.560 ;
        RECT  9.240 1.240 9.460 1.680 ;
        RECT  9.180 1.400 9.240 1.680 ;
        END
        ANTENNAGATEAREA 0.5832 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.800 1.390 6.020 2.340 ;
        RECT  5.740 1.390 5.800 1.960 ;
        RECT  5.640 1.270 5.740 1.960 ;
        RECT  5.520 1.270 5.640 1.550 ;
        END
        ANTENNAGATEAREA 0.8904 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.600 0.570 1.860 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 -0.280 10.800 0.280 ;
        RECT  10.480 -0.280 10.710 1.120 ;
        RECT  9.670 -0.280 10.480 0.280 ;
        RECT  9.390 -0.280 9.670 0.800 ;
        RECT  4.240 -0.280 9.390 0.280 ;
        RECT  3.960 -0.280 4.240 0.350 ;
        RECT  3.140 -0.280 3.960 0.280 ;
        RECT  2.980 -0.280 3.140 0.350 ;
        RECT  0.370 -0.280 2.980 0.280 ;
        RECT  0.090 -0.280 0.370 1.010 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.320 10.800 3.880 ;
        RECT  10.420 2.590 10.700 3.880 ;
        RECT  9.700 3.320 10.420 3.880 ;
        RECT  9.420 2.730 9.700 3.880 ;
        RECT  4.060 3.260 9.420 3.880 ;
        RECT  3.760 3.020 4.060 3.880 ;
        RECT  3.000 3.320 3.760 3.880 ;
        RECT  2.720 2.680 3.000 3.880 ;
        RECT  0.370 3.320 2.720 3.880 ;
        RECT  0.090 2.590 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.780 1.600 10.020 1.880 ;
        RECT  9.740 1.600 9.780 2.570 ;
        RECT  9.620 1.720 9.740 2.570 ;
        RECT  9.020 2.410 9.620 2.570 ;
        RECT  9.020 1.970 9.180 2.250 ;
        RECT  9.020 0.960 9.080 1.240 ;
        RECT  8.860 0.960 9.020 2.250 ;
        RECT  8.860 2.410 9.020 3.100 ;
        RECT  8.800 0.960 8.860 1.850 ;
        RECT  8.260 2.940 8.860 3.100 ;
        RECT  8.740 1.570 8.800 1.850 ;
        RECT  8.580 0.440 8.740 0.780 ;
        RECT  8.580 2.010 8.700 2.780 ;
        RECT  8.420 0.440 8.580 2.780 ;
        RECT  6.820 0.440 8.420 0.600 ;
        RECT  8.100 0.760 8.260 3.100 ;
        RECT  7.980 0.760 8.100 1.100 ;
        RECT  7.940 2.240 8.100 2.800 ;
        RECT  7.300 0.760 7.980 0.920 ;
        RECT  7.620 1.080 7.780 1.310 ;
        RECT  7.620 2.240 7.740 3.100 ;
        RECT  7.460 1.080 7.620 3.100 ;
        RECT  4.400 2.940 7.460 3.100 ;
        RECT  7.140 0.760 7.300 1.100 ;
        RECT  7.140 2.240 7.260 2.780 ;
        RECT  6.980 0.760 7.140 2.780 ;
        RECT  6.660 0.440 6.820 2.780 ;
        RECT  6.540 0.440 6.660 1.260 ;
        RECT  6.500 1.960 6.660 2.780 ;
        RECT  5.780 0.440 6.540 0.660 ;
        RECT  6.180 0.940 6.340 2.780 ;
        RECT  6.060 0.940 6.180 1.220 ;
        RECT  6.020 2.500 6.180 2.780 ;
        RECT  4.720 2.620 6.020 2.780 ;
        RECT  5.460 0.440 5.780 1.090 ;
        RECT  5.480 2.120 5.640 2.400 ;
        RECT  5.360 1.710 5.480 2.400 ;
        RECT  5.360 0.930 5.460 1.090 ;
        RECT  5.320 0.930 5.360 2.400 ;
        RECT  5.200 0.930 5.320 1.870 ;
        RECT  5.040 0.510 5.240 0.720 ;
        RECT  5.040 2.030 5.160 2.310 ;
        RECT  4.880 0.510 5.040 2.310 ;
        RECT  4.040 0.510 4.880 0.720 ;
        RECT  4.640 1.610 4.720 1.890 ;
        RECT  4.560 2.380 4.720 2.780 ;
        RECT  4.570 0.940 4.700 1.220 ;
        RECT  4.570 1.610 4.640 2.220 ;
        RECT  4.410 0.940 4.570 2.220 ;
        RECT  3.990 2.380 4.560 2.540 ;
        RECT  4.360 1.650 4.410 2.220 ;
        RECT  4.240 2.700 4.400 3.100 ;
        RECT  2.090 1.650 4.360 1.810 ;
        RECT  3.670 2.700 4.240 2.860 ;
        RECT  3.880 0.510 4.040 1.490 ;
        RECT  3.830 2.040 3.990 2.540 ;
        RECT  2.820 0.510 3.880 0.670 ;
        RECT  3.170 1.270 3.880 1.490 ;
        RECT  1.810 2.040 3.830 2.200 ;
        RECT  3.440 0.830 3.720 1.110 ;
        RECT  3.510 2.360 3.670 2.860 ;
        RECT  2.290 2.360 3.510 2.520 ;
        RECT  2.940 0.950 3.440 1.110 ;
        RECT  2.750 0.950 2.940 1.370 ;
        RECT  2.660 0.440 2.820 0.670 ;
        RECT  2.010 1.210 2.750 1.370 ;
        RECT  0.890 0.440 2.660 0.600 ;
        RECT  2.240 0.760 2.470 1.040 ;
        RECT  2.170 2.360 2.290 2.630 ;
        RECT  1.330 0.760 2.240 0.920 ;
        RECT  2.010 2.360 2.170 3.160 ;
        RECT  1.810 1.650 2.090 1.880 ;
        RECT  1.650 1.080 2.010 1.370 ;
        RECT  1.330 3.000 2.010 3.160 ;
        RECT  1.650 2.040 1.810 2.840 ;
        RECT  1.490 1.080 1.650 2.840 ;
        RECT  1.210 0.760 1.330 1.080 ;
        RECT  1.210 2.020 1.330 3.160 ;
        RECT  1.170 0.760 1.210 3.160 ;
        RECT  1.050 0.760 1.170 2.890 ;
        RECT  0.730 0.440 0.890 3.160 ;
        RECT  0.570 0.440 0.730 1.310 ;
        RECT  0.570 2.020 0.730 3.160 ;
    END
END XOR3X4TR

MACRO XOR3X2TR
    CLASS CORE ;
    FOREIGN XOR3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.360 0.440 7.520 3.160 ;
        RECT  7.230 0.440 7.360 1.310 ;
        RECT  7.280 1.920 7.360 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 2.360 6.750 2.760 ;
        END
        ANTENNAGATEAREA 0.2856 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 2.040 4.350 2.520 ;
        RECT  4.080 1.250 4.240 2.520 ;
        END
        ANTENNAGATEAREA 0.6408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.990 -0.280 7.600 0.280 ;
        RECT  6.710 -0.280 6.990 0.400 ;
        RECT  2.450 -0.280 6.710 0.340 ;
        RECT  2.290 -0.280 2.450 1.320 ;
        RECT  0.370 -0.280 2.290 0.280 ;
        RECT  0.090 -0.280 0.370 1.070 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 3.320 7.600 3.880 ;
        RECT  6.670 3.020 6.950 3.880 ;
        RECT  2.480 3.320 6.670 3.880 ;
        RECT  2.200 2.990 2.480 3.880 ;
        RECT  0.370 3.320 2.200 3.880 ;
        RECT  0.090 2.530 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.070 1.470 7.200 1.750 ;
        RECT  6.910 0.560 7.070 1.750 ;
        RECT  5.590 0.560 6.910 0.720 ;
        RECT  6.350 1.030 6.630 2.200 ;
        RECT  6.340 1.470 6.350 2.200 ;
        RECT  6.230 1.470 6.340 1.750 ;
        RECT  6.070 2.770 6.170 3.160 ;
        RECT  5.890 0.880 6.070 3.160 ;
        RECT  5.790 0.880 5.890 1.160 ;
        RECT  2.800 3.000 5.890 3.160 ;
        RECT  5.590 2.140 5.690 2.840 ;
        RECT  5.430 0.560 5.590 2.840 ;
        RECT  5.410 0.830 5.430 2.840 ;
        RECT  5.310 0.830 5.410 1.140 ;
        RECT  5.110 2.140 5.210 2.840 ;
        RECT  4.930 0.500 5.110 2.840 ;
        RECT  4.830 0.500 4.930 1.320 ;
        RECT  4.100 0.500 4.830 0.660 ;
        RECT  4.570 1.480 4.730 2.840 ;
        RECT  4.410 0.820 4.570 1.640 ;
        RECT  4.510 2.560 4.570 2.840 ;
        RECT  3.120 2.680 4.510 2.840 ;
        RECT  3.910 0.500 4.100 1.090 ;
        RECT  3.910 1.900 3.920 2.450 ;
        RECT  3.750 0.500 3.910 2.450 ;
        RECT  3.700 1.920 3.750 2.450 ;
        RECT  3.520 0.500 3.550 1.210 ;
        RECT  3.360 0.500 3.520 2.290 ;
        RECT  2.770 0.500 3.360 0.660 ;
        RECT  3.280 2.010 3.360 2.290 ;
        RECT  2.960 2.350 3.120 2.840 ;
        RECT  2.930 0.930 3.090 2.190 ;
        RECT  1.430 2.350 2.960 2.510 ;
        RECT  1.750 2.030 2.930 2.190 ;
        RECT  2.640 2.670 2.800 3.160 ;
        RECT  2.610 0.500 2.770 1.640 ;
        RECT  1.110 2.670 2.640 2.830 ;
        RECT  2.250 1.480 2.610 1.640 ;
        RECT  2.130 1.480 2.250 1.760 ;
        RECT  1.970 0.440 2.130 1.760 ;
        RECT  0.790 0.440 1.970 0.600 ;
        RECT  1.530 0.790 1.810 1.360 ;
        RECT  1.590 1.520 1.750 2.190 ;
        RECT  1.430 1.200 1.530 1.360 ;
        RECT  1.270 1.200 1.430 2.510 ;
        RECT  1.110 0.760 1.330 1.040 ;
        RECT  0.950 0.760 1.110 2.830 ;
        RECT  0.570 0.440 0.790 3.160 ;
    END
END XOR3X2TR

MACRO XOR3X1TR
    CLASS CORE ;
    FOREIGN XOR3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 0.920 7.520 2.550 ;
        RECT  7.200 0.920 7.280 1.200 ;
        RECT  7.250 1.910 7.280 2.550 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.400 2.380 6.720 2.760 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.640 4.420 2.180 ;
        RECT  4.200 1.640 4.260 1.960 ;
        RECT  4.040 1.180 4.200 1.960 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.380 1.960 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.940 -0.280 7.600 0.280 ;
        RECT  6.660 -0.280 6.940 0.340 ;
        RECT  1.840 -0.280 6.660 0.280 ;
        RECT  1.560 -0.280 1.840 0.580 ;
        RECT  0.400 -0.280 1.560 0.280 ;
        RECT  0.090 -0.280 0.400 0.560 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 3.320 7.600 3.880 ;
        RECT  6.670 2.920 6.950 3.880 ;
        RECT  2.340 3.320 6.670 3.880 ;
        RECT  2.060 2.930 2.340 3.880 ;
        RECT  0.410 3.320 2.060 3.880 ;
        RECT  0.100 3.260 0.410 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.840 1.360 7.120 1.640 ;
        RECT  6.680 0.590 6.840 1.640 ;
        RECT  5.380 0.590 6.680 0.750 ;
        RECT  6.160 1.030 6.320 2.190 ;
        RECT  5.860 1.500 6.160 1.660 ;
        RECT  5.860 2.370 6.020 2.650 ;
        RECT  5.700 0.910 5.920 1.070 ;
        RECT  5.700 1.820 5.860 3.000 ;
        RECT  5.540 0.910 5.700 1.980 ;
        RECT  2.660 2.840 5.700 3.000 ;
        RECT  5.380 2.140 5.540 2.650 ;
        RECT  5.220 0.590 5.380 2.300 ;
        RECT  4.900 0.830 5.060 2.650 ;
        RECT  4.840 0.830 4.900 0.990 ;
        RECT  4.680 0.540 4.840 0.990 ;
        RECT  4.580 1.150 4.740 2.680 ;
        RECT  3.880 0.540 4.680 0.700 ;
        RECT  4.520 1.150 4.580 1.310 ;
        RECT  3.240 2.520 4.580 2.680 ;
        RECT  4.360 0.860 4.520 1.310 ;
        RECT  4.200 0.860 4.360 1.020 ;
        RECT  3.880 2.200 4.100 2.360 ;
        RECT  3.720 0.540 3.880 2.360 ;
        RECT  3.400 0.450 3.560 2.190 ;
        RECT  2.160 0.450 3.400 0.610 ;
        RECT  3.080 0.770 3.240 2.680 ;
        RECT  2.480 0.770 3.080 0.930 ;
        RECT  2.760 1.090 2.920 2.450 ;
        RECT  2.640 1.090 2.760 1.250 ;
        RECT  2.640 2.170 2.760 2.450 ;
        RECT  2.500 2.610 2.660 3.000 ;
        RECT  1.400 2.290 2.640 2.450 ;
        RECT  1.080 2.610 2.500 2.770 ;
        RECT  2.320 0.770 2.480 2.130 ;
        RECT  1.720 1.970 2.320 2.130 ;
        RECT  2.000 0.450 2.160 1.580 ;
        RECT  0.760 0.770 2.000 0.930 ;
        RECT  1.880 1.420 2.000 1.580 ;
        RECT  1.720 1.090 1.840 1.250 ;
        RECT  1.560 1.090 1.720 2.130 ;
        RECT  1.240 1.700 1.400 2.450 ;
        RECT  1.080 1.090 1.320 1.250 ;
        RECT  0.920 1.090 1.080 2.770 ;
        RECT  0.600 0.770 0.760 2.950 ;
    END
END XOR3X1TR

MACRO XOR2XLTR
    CLASS CORE ;
    FOREIGN XOR2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.950 2.320 2.560 ;
        RECT  1.980 0.950 2.040 1.230 ;
        RECT  1.980 2.280 2.040 2.560 ;
        END
        ANTENNADIFFAREA 1.893 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.100 1.180 1.380 ;
        RECT  0.900 1.100 1.120 1.560 ;
        RECT  0.840 1.220 0.900 1.560 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 2.720 0.720 3.160 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 -0.280 3.200 0.280 ;
        RECT  1.040 -0.280 2.760 0.340 ;
        RECT  0.760 -0.280 1.040 0.940 ;
        RECT  0.000 -0.280 0.760 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 3.320 3.200 3.880 ;
        RECT  2.480 3.200 2.760 3.880 ;
        RECT  1.160 3.260 2.480 3.880 ;
        RECT  0.880 2.330 1.160 3.880 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 0.630 3.080 1.550 ;
        RECT  1.820 0.630 2.920 0.790 ;
        RECT  2.480 0.950 2.760 3.000 ;
        RECT  1.660 0.630 1.820 2.370 ;
        RECT  1.340 0.770 1.660 1.050 ;
        RECT  1.640 2.210 1.660 2.370 ;
        RECT  1.360 2.210 1.640 2.490 ;
        RECT  1.280 1.540 1.500 1.880 ;
        RECT  0.480 1.720 1.280 1.880 ;
        RECT  0.320 0.850 0.480 2.490 ;
        RECT  0.200 0.850 0.320 1.130 ;
        RECT  0.200 2.210 0.320 2.490 ;
    END
END XOR2XLTR

MACRO XOR2X4TR
    CLASS CORE ;
    FOREIGN XOR2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.580 0.910 5.860 1.190 ;
        RECT  5.520 1.970 5.700 2.330 ;
        RECT  5.520 0.950 5.580 1.190 ;
        RECT  5.420 0.950 5.520 2.330 ;
        RECT  5.280 0.950 5.420 2.210 ;
        RECT  4.900 0.950 5.280 1.190 ;
        RECT  4.740 1.960 5.280 2.210 ;
        RECT  4.620 0.470 4.900 1.190 ;
        RECT  4.460 1.960 4.740 2.330 ;
        RECT  3.940 0.950 4.620 1.190 ;
        RECT  3.780 1.960 4.460 2.210 ;
        RECT  3.660 0.910 3.940 1.190 ;
        RECT  3.500 1.960 3.780 2.330 ;
        END
        ANTENNADIFFAREA 9.504 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.610 1.180 1.960 ;
        END
        ANTENNAGATEAREA 0.6384 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.470 2.700 1.750 ;
        RECT  2.320 1.590 2.480 1.750 ;
        RECT  2.040 1.240 2.320 1.750 ;
        END
        ANTENNAGATEAREA 0.8856 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.780 -0.280 8.000 0.280 ;
        RECT  7.500 -0.280 7.780 1.190 ;
        RECT  6.820 -0.280 7.500 0.280 ;
        RECT  6.540 -0.280 6.820 0.750 ;
        RECT  2.460 -0.280 6.540 0.280 ;
        RECT  2.180 -0.280 2.460 0.400 ;
        RECT  1.460 -0.280 2.180 0.340 ;
        RECT  1.180 -0.280 1.460 1.040 ;
        RECT  0.460 -0.280 1.180 0.340 ;
        RECT  0.180 -0.280 0.460 1.260 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.880 3.320 8.000 3.880 ;
        RECT  7.600 3.200 7.880 3.880 ;
        RECT  7.000 3.260 7.600 3.880 ;
        RECT  6.720 2.110 7.000 3.880 ;
        RECT  2.440 3.260 6.720 3.880 ;
        RECT  2.160 3.100 2.440 3.880 ;
        RECT  1.460 3.260 2.160 3.880 ;
        RECT  1.180 2.440 1.460 3.880 ;
        RECT  0.460 3.260 1.180 3.880 ;
        RECT  0.180 2.220 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.340 1.790 7.480 2.890 ;
        RECT  7.200 0.470 7.340 2.890 ;
        RECT  7.180 0.470 7.200 1.950 ;
        RECT  7.020 0.470 7.180 1.190 ;
        RECT  6.520 1.790 7.180 1.950 ;
        RECT  6.340 1.030 7.020 1.190 ;
        RECT  6.340 1.350 7.020 1.630 ;
        RECT  6.360 1.790 6.520 3.090 ;
        RECT  6.240 1.910 6.360 2.190 ;
        RECT  3.020 2.810 6.360 3.090 ;
        RECT  6.060 0.470 6.340 1.190 ;
        RECT  6.060 1.470 6.340 1.630 ;
        RECT  6.060 2.370 6.180 2.650 ;
        RECT  5.380 0.470 6.060 0.630 ;
        RECT  5.900 1.470 6.060 2.650 ;
        RECT  5.220 2.490 5.900 2.650 ;
        RECT  5.100 0.470 5.380 0.750 ;
        RECT  4.940 2.370 5.220 2.650 ;
        RECT  4.740 1.350 5.120 1.630 ;
        RECT  1.940 2.490 4.940 2.650 ;
        RECT  3.020 1.350 4.740 1.510 ;
        RECT  4.140 0.460 4.420 0.750 ;
        RECT  3.460 0.460 4.140 0.630 ;
        RECT  3.180 0.460 3.460 1.190 ;
        RECT  1.940 0.710 3.180 0.870 ;
        RECT  2.860 1.030 3.020 2.190 ;
        RECT  2.700 1.030 2.860 1.310 ;
        RECT  2.680 1.910 2.860 2.190 ;
        RECT  1.780 0.710 1.940 1.040 ;
        RECT  1.780 2.120 1.940 2.650 ;
        RECT  1.660 0.760 1.780 2.650 ;
        RECT  1.620 0.760 1.660 2.280 ;
        RECT  0.980 1.200 1.620 1.360 ;
        RECT  0.980 2.120 1.620 2.280 ;
        RECT  0.820 1.030 0.980 1.360 ;
        RECT  0.700 2.120 0.980 2.720 ;
        RECT  0.700 1.030 0.820 1.310 ;
    END
END XOR2X4TR

MACRO XOR2X2TR
    CLASS CORE ;
    FOREIGN XOR2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.990 0.840 5.120 2.950 ;
        RECT  4.830 0.590 4.990 2.950 ;
        RECT  4.150 0.590 4.830 0.750 ;
        RECT  3.990 0.590 4.150 2.780 ;
        RECT  3.870 0.590 3.990 1.020 ;
        RECT  3.870 2.170 3.990 2.780 ;
        RECT  3.230 0.590 3.870 0.750 ;
        RECT  3.070 0.590 3.230 2.450 ;
        RECT  2.910 0.920 3.070 1.200 ;
        RECT  2.910 2.170 3.070 2.450 ;
        END
        ANTENNADIFFAREA 6.602 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.360 0.970 1.640 ;
        RECT  0.440 1.240 0.760 1.640 ;
        RECT  0.330 1.360 0.440 1.640 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.640 2.430 1.960 ;
        RECT  2.040 1.630 2.260 1.960 ;
        END
        ANTENNAGATEAREA 0.444 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.280 5.200 0.280 ;
        RECT  0.930 -0.280 1.210 0.400 ;
        RECT  0.410 -0.280 0.930 0.280 ;
        RECT  0.130 -0.280 0.410 0.400 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 3.320 5.200 3.880 ;
        RECT  0.410 3.260 2.480 3.880 ;
        RECT  0.130 3.200 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.510 0.910 4.630 1.190 ;
        RECT  4.510 2.170 4.630 2.950 ;
        RECT  4.350 0.910 4.510 3.100 ;
        RECT  1.290 2.940 4.350 3.100 ;
        RECT  3.510 1.010 3.670 2.780 ;
        RECT  3.390 1.010 3.510 1.290 ;
        RECT  3.390 2.170 3.510 2.780 ;
        RECT  1.790 2.620 3.390 2.780 ;
        RECT  2.750 1.360 2.910 1.640 ;
        RECT  2.590 0.960 2.750 2.400 ;
        RECT  2.430 0.960 2.590 1.240 ;
        RECT  2.430 2.120 2.590 2.400 ;
        RECT  1.730 1.030 1.790 1.310 ;
        RECT  1.730 2.030 1.790 2.780 ;
        RECT  1.570 1.030 1.730 2.780 ;
        RECT  1.510 1.030 1.570 1.310 ;
        RECT  1.290 1.360 1.350 1.640 ;
        RECT  1.130 0.920 1.290 3.100 ;
        RECT  0.810 0.920 1.130 1.080 ;
        RECT  0.810 2.030 1.130 2.190 ;
        RECT  0.530 0.800 0.810 1.080 ;
        RECT  0.530 2.030 0.810 2.810 ;
    END
END XOR2X2TR

MACRO XOR2X1TR
    CLASS CORE ;
    FOREIGN XOR2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.910 2.150 2.760 ;
        RECT  1.650 0.910 1.990 1.190 ;
        RECT  1.640 2.440 1.990 2.760 ;
        END
        ANTENNADIFFAREA 2.603 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.240 1.160 1.560 ;
        RECT  0.820 1.240 1.130 1.630 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 2.440 0.720 2.760 ;
        END
        ANTENNAGATEAREA 0.2184 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.280 3.200 0.280 ;
        RECT  2.830 -0.280 3.110 0.400 ;
        RECT  0.970 -0.280 2.830 0.340 ;
        RECT  0.690 -0.280 0.970 1.020 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 3.320 3.200 3.880 ;
        RECT  2.790 2.240 3.070 3.880 ;
        RECT  0.930 3.260 2.790 3.880 ;
        RECT  0.650 2.920 0.930 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.910 1.540 3.030 1.820 ;
        RECT  2.750 0.590 2.910 1.820 ;
        RECT  1.490 0.590 2.750 0.750 ;
        RECT  2.310 0.980 2.590 2.950 ;
        RECT  1.670 1.350 1.830 2.270 ;
        RECT  1.490 1.350 1.670 1.510 ;
        RECT  1.450 2.110 1.670 2.270 ;
        RECT  1.290 1.670 1.510 1.950 ;
        RECT  1.330 0.590 1.490 1.510 ;
        RECT  1.170 2.110 1.450 2.590 ;
        RECT  1.170 0.740 1.330 1.020 ;
        RECT  0.450 1.790 1.290 1.950 ;
        RECT  0.410 1.790 0.450 2.280 ;
        RECT  0.250 0.980 0.410 2.280 ;
        RECT  0.090 0.980 0.250 1.260 ;
        RECT  0.130 2.000 0.250 2.280 ;
    END
END XOR2X1TR

MACRO XNOR3XLTR
    CLASS CORE ;
    FOREIGN XNOR3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.030 7.520 3.160 ;
        RECT  7.280 2.040 7.290 3.160 ;
        END
        ANTENNADIFFAREA 1.202 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.480 2.350 6.720 2.830 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.300 1.640 4.460 2.360 ;
        RECT  4.200 1.640 4.300 1.960 ;
        RECT  4.040 1.180 4.200 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.440 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.070 -0.280 7.600 0.280 ;
        RECT  6.780 -0.280 7.070 0.340 ;
        RECT  1.840 -0.280 6.780 0.280 ;
        RECT  1.560 -0.280 1.840 0.610 ;
        RECT  0.360 -0.280 1.560 0.280 ;
        RECT  0.090 -0.280 0.360 0.770 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.040 3.320 7.600 3.880 ;
        RECT  6.880 1.970 7.040 3.880 ;
        RECT  6.710 1.970 6.880 2.130 ;
        RECT  2.300 3.320 6.880 3.880 ;
        RECT  2.020 2.930 2.300 3.880 ;
        RECT  0.380 3.320 2.020 3.880 ;
        RECT  0.120 3.190 0.380 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.970 0.540 7.130 1.750 ;
        RECT  5.430 0.540 6.970 0.700 ;
        RECT  6.330 0.910 6.490 2.190 ;
        RECT  6.290 0.910 6.330 1.620 ;
        RECT  6.060 1.460 6.290 1.620 ;
        RECT  5.900 0.890 6.120 1.050 ;
        RECT  6.110 2.450 6.120 2.740 ;
        RECT  5.950 1.800 6.110 3.070 ;
        RECT  5.900 1.800 5.950 1.960 ;
        RECT  2.620 2.910 5.950 3.070 ;
        RECT  5.740 0.890 5.900 1.960 ;
        RECT  5.480 2.130 5.640 2.740 ;
        RECT  5.430 2.130 5.480 2.290 ;
        RECT  5.270 0.540 5.430 2.290 ;
        RECT  4.940 0.830 5.100 2.740 ;
        RECT  4.890 0.830 4.940 1.110 ;
        RECT  4.710 0.450 4.890 1.110 ;
        RECT  4.620 1.320 4.780 2.680 ;
        RECT  3.880 0.450 4.710 0.610 ;
        RECT  4.530 1.320 4.620 1.480 ;
        RECT  3.240 2.520 4.620 2.680 ;
        RECT  4.370 0.840 4.530 1.480 ;
        RECT  4.090 0.840 4.370 1.000 ;
        RECT  3.880 2.120 4.040 2.360 ;
        RECT  3.720 0.450 3.880 2.330 ;
        RECT  3.400 0.450 3.560 2.360 ;
        RECT  2.160 0.450 3.400 0.610 ;
        RECT  3.080 0.770 3.240 2.680 ;
        RECT  2.480 0.770 3.080 0.930 ;
        RECT  2.640 1.090 2.920 2.450 ;
        RECT  1.400 2.290 2.640 2.450 ;
        RECT  2.460 2.610 2.620 3.070 ;
        RECT  2.320 0.770 2.480 2.130 ;
        RECT  1.080 2.610 2.460 2.770 ;
        RECT  1.720 1.970 2.320 2.130 ;
        RECT  2.000 0.450 2.160 1.790 ;
        RECT  0.850 0.770 2.000 0.930 ;
        RECT  1.900 1.510 2.000 1.790 ;
        RECT  1.720 1.090 1.840 1.310 ;
        RECT  1.560 1.090 1.720 2.130 ;
        RECT  1.240 1.960 1.400 2.450 ;
        RECT  1.080 1.090 1.320 1.250 ;
        RECT  0.920 1.090 1.080 2.770 ;
        RECT  0.760 0.510 0.850 0.930 ;
        RECT  0.600 0.510 0.760 2.830 ;
    END
END XNOR3XLTR

MACRO XNOR3X4TR
    CLASS CORE ;
    FOREIGN XNOR3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.320 1.280 10.420 2.280 ;
        RECT  10.220 0.440 10.320 2.280 ;
        RECT  10.180 0.440 10.220 3.160 ;
        RECT  9.910 0.440 10.180 1.440 ;
        RECT  9.940 2.040 10.180 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.460 1.240 9.560 1.560 ;
        RECT  9.280 1.240 9.460 1.680 ;
        RECT  9.180 1.400 9.280 1.680 ;
        END
        ANTENNAGATEAREA 0.5544 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.800 1.390 6.020 2.340 ;
        RECT  5.740 1.390 5.800 1.960 ;
        RECT  5.640 1.270 5.740 1.960 ;
        RECT  5.520 1.270 5.640 1.550 ;
        END
        ANTENNAGATEAREA 0.8904 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.600 0.570 1.860 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 -0.280 10.800 0.280 ;
        RECT  10.480 -0.280 10.710 1.120 ;
        RECT  9.670 -0.280 10.480 0.280 ;
        RECT  9.390 -0.280 9.670 0.800 ;
        RECT  4.240 -0.280 9.390 0.280 ;
        RECT  3.960 -0.280 4.240 0.350 ;
        RECT  3.140 -0.280 3.960 0.280 ;
        RECT  2.980 -0.280 3.140 0.350 ;
        RECT  0.370 -0.280 2.980 0.280 ;
        RECT  0.090 -0.280 0.370 1.010 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.320 10.800 3.880 ;
        RECT  10.420 2.590 10.700 3.880 ;
        RECT  9.700 3.320 10.420 3.880 ;
        RECT  9.420 2.730 9.700 3.880 ;
        RECT  4.060 3.260 9.420 3.880 ;
        RECT  3.760 3.020 4.060 3.880 ;
        RECT  3.000 3.320 3.760 3.880 ;
        RECT  2.710 2.680 3.000 3.880 ;
        RECT  0.370 3.320 2.710 3.880 ;
        RECT  0.090 2.590 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.780 1.600 10.020 1.880 ;
        RECT  9.740 1.600 9.780 2.570 ;
        RECT  9.620 1.720 9.740 2.570 ;
        RECT  9.020 2.410 9.620 2.570 ;
        RECT  9.020 1.970 9.180 2.250 ;
        RECT  9.020 0.960 9.090 1.240 ;
        RECT  8.860 0.960 9.020 2.250 ;
        RECT  8.860 2.410 9.020 3.100 ;
        RECT  8.800 0.960 8.860 1.850 ;
        RECT  8.260 2.940 8.860 3.100 ;
        RECT  8.740 1.570 8.800 1.850 ;
        RECT  8.580 0.440 8.740 0.780 ;
        RECT  8.580 2.310 8.700 2.690 ;
        RECT  8.420 0.440 8.580 2.690 ;
        RECT  6.820 0.440 8.420 0.600 ;
        RECT  8.100 0.760 8.260 3.100 ;
        RECT  7.980 0.760 8.100 1.100 ;
        RECT  7.940 2.240 8.100 2.800 ;
        RECT  7.300 0.760 7.980 0.920 ;
        RECT  7.620 1.080 7.780 1.310 ;
        RECT  7.620 1.960 7.680 3.100 ;
        RECT  7.460 1.080 7.620 3.100 ;
        RECT  4.400 2.940 7.460 3.100 ;
        RECT  7.140 0.760 7.300 1.100 ;
        RECT  7.140 2.240 7.260 2.780 ;
        RECT  6.980 0.760 7.140 2.780 ;
        RECT  6.660 0.440 6.820 2.780 ;
        RECT  6.540 0.440 6.660 1.260 ;
        RECT  6.500 2.460 6.660 2.780 ;
        RECT  5.780 0.440 6.540 0.660 ;
        RECT  6.180 0.940 6.340 2.780 ;
        RECT  6.060 0.940 6.180 1.220 ;
        RECT  6.020 2.500 6.180 2.780 ;
        RECT  4.720 2.620 6.020 2.780 ;
        RECT  5.460 0.440 5.780 1.090 ;
        RECT  5.480 2.120 5.640 2.400 ;
        RECT  5.360 1.710 5.480 2.400 ;
        RECT  5.360 0.930 5.460 1.090 ;
        RECT  5.320 0.930 5.360 2.400 ;
        RECT  5.200 0.930 5.320 1.870 ;
        RECT  5.040 0.510 5.240 0.720 ;
        RECT  5.040 2.030 5.160 2.310 ;
        RECT  4.880 0.510 5.040 2.310 ;
        RECT  4.040 0.510 4.880 0.720 ;
        RECT  4.640 1.610 4.720 1.890 ;
        RECT  4.560 2.380 4.720 2.780 ;
        RECT  4.570 0.940 4.700 1.220 ;
        RECT  4.570 1.610 4.640 2.220 ;
        RECT  4.410 0.940 4.570 2.220 ;
        RECT  3.990 2.380 4.560 2.540 ;
        RECT  4.360 1.650 4.410 2.220 ;
        RECT  4.240 2.700 4.400 3.100 ;
        RECT  2.090 1.650 4.360 1.810 ;
        RECT  3.670 2.700 4.240 2.860 ;
        RECT  3.880 0.510 4.040 1.490 ;
        RECT  3.830 2.040 3.990 2.540 ;
        RECT  2.820 0.510 3.880 0.670 ;
        RECT  3.170 1.270 3.880 1.490 ;
        RECT  1.810 2.040 3.830 2.200 ;
        RECT  3.440 0.830 3.720 1.110 ;
        RECT  3.510 2.360 3.670 2.860 ;
        RECT  2.290 2.360 3.510 2.520 ;
        RECT  2.940 0.950 3.440 1.110 ;
        RECT  2.750 0.950 2.940 1.370 ;
        RECT  2.660 0.440 2.820 0.670 ;
        RECT  2.010 1.210 2.750 1.370 ;
        RECT  0.890 0.440 2.660 0.600 ;
        RECT  2.240 0.760 2.470 1.040 ;
        RECT  2.170 2.360 2.290 2.630 ;
        RECT  1.330 0.760 2.240 0.920 ;
        RECT  2.010 2.360 2.170 3.160 ;
        RECT  1.810 1.650 2.090 1.880 ;
        RECT  1.650 1.080 2.010 1.370 ;
        RECT  1.330 3.000 2.010 3.160 ;
        RECT  1.650 2.040 1.810 2.840 ;
        RECT  1.490 1.080 1.650 2.840 ;
        RECT  1.210 0.760 1.330 1.080 ;
        RECT  1.210 2.020 1.330 3.160 ;
        RECT  1.170 0.760 1.210 3.160 ;
        RECT  1.050 0.760 1.170 2.890 ;
        RECT  0.730 0.440 0.890 3.160 ;
        RECT  0.570 0.440 0.730 1.310 ;
        RECT  0.570 2.020 0.730 3.160 ;
    END
END XNOR3X4TR

MACRO XNOR3X2TR
    CLASS CORE ;
    FOREIGN XNOR3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.360 0.440 7.520 3.160 ;
        RECT  7.230 0.440 7.360 1.310 ;
        RECT  7.280 1.920 7.360 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 2.360 6.750 2.760 ;
        END
        ANTENNAGATEAREA 0.2976 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 2.040 4.350 2.380 ;
        RECT  4.080 1.210 4.250 2.380 ;
        END
        ANTENNAGATEAREA 0.6408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.990 -0.280 7.600 0.280 ;
        RECT  6.710 -0.280 6.990 0.400 ;
        RECT  2.450 -0.280 6.710 0.340 ;
        RECT  2.290 -0.280 2.450 1.320 ;
        RECT  0.370 -0.280 2.290 0.280 ;
        RECT  0.090 -0.280 0.370 1.070 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 3.320 7.600 3.880 ;
        RECT  6.670 3.020 6.950 3.880 ;
        RECT  2.480 3.320 6.670 3.880 ;
        RECT  2.200 2.990 2.480 3.880 ;
        RECT  0.370 3.320 2.200 3.880 ;
        RECT  0.090 2.530 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.070 1.470 7.200 1.750 ;
        RECT  6.910 0.560 7.070 1.750 ;
        RECT  5.590 0.560 6.910 0.720 ;
        RECT  6.350 0.940 6.630 2.200 ;
        RECT  6.340 1.470 6.350 2.200 ;
        RECT  6.230 1.470 6.340 1.750 ;
        RECT  6.070 2.020 6.170 2.890 ;
        RECT  6.050 0.880 6.070 2.890 ;
        RECT  5.890 0.880 6.050 3.160 ;
        RECT  5.790 0.880 5.890 1.160 ;
        RECT  2.800 3.000 5.890 3.160 ;
        RECT  5.590 2.140 5.690 2.840 ;
        RECT  5.430 0.560 5.590 2.840 ;
        RECT  5.410 0.650 5.430 2.840 ;
        RECT  5.310 0.650 5.410 0.930 ;
        RECT  5.110 2.140 5.210 2.840 ;
        RECT  4.930 0.500 5.110 2.840 ;
        RECT  4.830 0.500 4.930 1.320 ;
        RECT  4.100 0.500 4.830 0.660 ;
        RECT  4.570 1.480 4.730 2.840 ;
        RECT  4.410 0.820 4.570 1.640 ;
        RECT  4.510 2.560 4.570 2.840 ;
        RECT  3.120 2.680 4.510 2.840 ;
        RECT  3.910 0.500 4.100 1.000 ;
        RECT  3.910 2.140 3.920 2.450 ;
        RECT  3.750 0.500 3.910 2.450 ;
        RECT  3.700 2.150 3.750 2.450 ;
        RECT  3.520 0.500 3.550 1.210 ;
        RECT  3.360 0.500 3.520 2.290 ;
        RECT  2.770 0.500 3.360 0.660 ;
        RECT  3.280 2.010 3.360 2.290 ;
        RECT  2.960 2.350 3.120 2.840 ;
        RECT  2.930 0.930 3.090 2.190 ;
        RECT  1.430 2.350 2.960 2.510 ;
        RECT  1.750 2.030 2.930 2.190 ;
        RECT  2.640 2.670 2.800 3.160 ;
        RECT  2.610 0.500 2.770 1.640 ;
        RECT  1.110 2.670 2.640 2.830 ;
        RECT  2.250 1.480 2.610 1.640 ;
        RECT  2.130 1.480 2.250 1.760 ;
        RECT  1.970 0.440 2.130 1.760 ;
        RECT  0.790 0.440 1.970 0.600 ;
        RECT  1.530 0.790 1.810 1.360 ;
        RECT  1.590 1.520 1.750 2.190 ;
        RECT  1.430 1.200 1.530 1.360 ;
        RECT  1.270 1.200 1.430 2.510 ;
        RECT  1.110 0.760 1.330 1.040 ;
        RECT  0.950 0.760 1.110 2.830 ;
        RECT  0.570 0.440 0.790 3.160 ;
    END
END XNOR3X2TR

MACRO XNOR3X1TR
    CLASS CORE ;
    FOREIGN XNOR3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.380 2.020 7.520 3.160 ;
        RECT  7.210 0.920 7.380 3.160 ;
        END
        ANTENNADIFFAREA 1.879 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 2.380 6.720 2.920 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.640 4.370 2.180 ;
        RECT  4.040 1.180 4.200 1.960 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.380 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.000 -0.280 7.600 0.280 ;
        RECT  6.710 -0.280 7.000 0.340 ;
        RECT  1.840 -0.280 6.710 0.280 ;
        RECT  1.560 -0.280 1.840 0.580 ;
        RECT  0.370 -0.280 1.560 0.280 ;
        RECT  0.090 -0.280 0.370 0.450 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.040 3.320 7.600 3.880 ;
        RECT  6.880 1.970 7.040 3.880 ;
        RECT  6.620 1.970 6.880 2.130 ;
        RECT  2.340 3.320 6.880 3.880 ;
        RECT  2.060 2.930 2.340 3.880 ;
        RECT  0.340 3.320 2.060 3.880 ;
        RECT  0.090 3.180 0.340 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.890 0.590 7.050 1.640 ;
        RECT  5.430 0.590 6.890 0.750 ;
        RECT  6.210 0.920 6.430 2.190 ;
        RECT  6.150 0.920 6.210 1.790 ;
        RECT  5.970 1.500 6.150 1.790 ;
        RECT  5.810 0.910 5.970 1.070 ;
        RECT  5.810 2.370 5.970 2.650 ;
        RECT  5.650 0.910 5.810 3.160 ;
        RECT  2.660 3.000 5.650 3.160 ;
        RECT  5.430 2.370 5.490 2.650 ;
        RECT  5.270 0.590 5.430 2.650 ;
        RECT  4.850 0.540 5.010 2.650 ;
        RECT  4.730 0.540 4.850 0.990 ;
        RECT  3.880 0.540 4.730 0.700 ;
        RECT  4.530 1.150 4.690 2.810 ;
        RECT  4.370 0.860 4.530 1.310 ;
        RECT  3.240 2.650 4.530 2.810 ;
        RECT  4.250 0.860 4.370 1.020 ;
        RECT  3.880 2.330 4.100 2.490 ;
        RECT  3.720 0.540 3.880 2.490 ;
        RECT  3.400 0.450 3.560 2.190 ;
        RECT  2.160 0.450 3.400 0.610 ;
        RECT  3.080 0.770 3.240 2.810 ;
        RECT  2.480 0.770 3.080 0.930 ;
        RECT  2.640 1.090 2.920 2.450 ;
        RECT  2.500 2.610 2.660 3.160 ;
        RECT  1.400 2.290 2.640 2.450 ;
        RECT  1.080 2.610 2.500 2.770 ;
        RECT  2.320 0.770 2.480 2.130 ;
        RECT  1.720 1.970 2.320 2.130 ;
        RECT  2.000 0.450 2.160 1.690 ;
        RECT  0.760 0.770 2.000 0.930 ;
        RECT  1.900 1.410 2.000 1.690 ;
        RECT  1.720 1.090 1.840 1.250 ;
        RECT  1.560 1.090 1.720 2.130 ;
        RECT  1.240 1.700 1.400 2.450 ;
        RECT  1.080 1.090 1.320 1.250 ;
        RECT  0.920 1.090 1.080 2.770 ;
        RECT  0.600 0.770 0.760 2.950 ;
    END
END XNOR3X1TR

MACRO XNOR2XLTR
    CLASS CORE ;
    FOREIGN XNOR2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.180 1.210 2.320 1.570 ;
        RECT  1.890 0.970 2.180 2.490 ;
        END
        ANTENNADIFFAREA 1.768 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.840 1.120 1.380 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 2.820 0.720 3.160 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.800 -0.280 3.200 0.280 ;
        RECT  0.930 -0.280 2.800 0.340 ;
        RECT  0.650 -0.280 0.930 0.680 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.730 3.320 3.200 3.880 ;
        RECT  2.450 3.200 2.730 3.880 ;
        RECT  1.050 3.260 2.450 3.880 ;
        RECT  0.880 2.330 1.050 3.880 ;
        RECT  0.770 2.330 0.880 2.620 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.960 0.630 3.120 1.710 ;
        RECT  1.730 0.630 2.960 0.790 ;
        RECT  2.840 1.430 2.960 1.710 ;
        RECT  2.680 0.950 2.800 1.230 ;
        RECT  2.680 2.210 2.800 3.000 ;
        RECT  2.520 0.950 2.680 3.000 ;
        RECT  1.570 0.630 1.730 2.370 ;
        RECT  1.310 0.770 1.570 1.050 ;
        RECT  1.530 2.210 1.570 2.370 ;
        RECT  1.250 2.210 1.530 2.490 ;
        RECT  1.130 1.540 1.410 1.820 ;
        RECT  0.370 1.660 1.130 1.820 ;
        RECT  0.210 0.850 0.370 2.490 ;
        RECT  0.090 0.850 0.210 1.130 ;
        RECT  0.090 2.210 0.210 2.490 ;
    END
END XNOR2XLTR

MACRO XNOR2X4TR
    CLASS CORE ;
    FOREIGN XNOR2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.260 0.800 5.480 1.030 ;
        RECT  4.880 0.800 5.260 2.460 ;
        RECT  4.520 0.800 4.880 1.040 ;
        RECT  3.060 2.180 4.880 2.460 ;
        RECT  4.240 0.440 4.520 1.040 ;
        RECT  3.560 0.800 4.240 1.040 ;
        RECT  3.280 0.760 3.560 1.040 ;
        END
        ANTENNADIFFAREA 9.396 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.520 1.050 1.720 ;
        RECT  0.370 1.520 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.6336 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.640 4.020 1.960 ;
        END
        ANTENNAGATEAREA 0.8784 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.460 -0.280 7.600 0.280 ;
        RECT  7.180 -0.280 7.460 1.090 ;
        RECT  6.490 -0.280 7.180 0.280 ;
        RECT  6.220 -0.280 6.490 0.670 ;
        RECT  1.850 -0.280 6.220 0.280 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  0.850 -0.280 1.570 0.340 ;
        RECT  0.570 -0.280 0.850 0.930 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.460 3.320 7.600 3.880 ;
        RECT  7.180 1.910 7.460 3.880 ;
        RECT  6.460 3.320 7.180 3.880 ;
        RECT  6.220 2.010 6.460 3.880 ;
        RECT  1.810 3.320 6.220 3.880 ;
        RECT  1.530 2.670 1.810 3.880 ;
        RECT  0.850 3.260 1.530 3.880 ;
        RECT  0.570 2.670 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.860 0.600 7.020 2.950 ;
        RECT  6.700 0.600 6.860 1.090 ;
        RECT  6.700 1.690 6.860 2.950 ;
        RECT  5.960 0.930 6.700 1.090 ;
        RECT  6.020 1.690 6.700 1.850 ;
        RECT  6.000 1.250 6.640 1.530 ;
        RECT  5.740 1.690 6.020 3.160 ;
        RECT  5.580 1.370 6.000 1.530 ;
        RECT  5.680 0.480 5.960 1.090 ;
        RECT  4.500 2.940 5.740 3.160 ;
        RECT  4.720 0.480 5.680 0.640 ;
        RECT  5.420 1.370 5.580 2.780 ;
        RECT  3.830 2.620 5.420 2.780 ;
        RECT  4.280 1.260 4.590 2.020 ;
        RECT  2.370 1.260 4.280 1.420 ;
        RECT  3.740 0.440 4.040 0.640 ;
        RECT  3.550 2.620 3.830 2.890 ;
        RECT  3.060 0.440 3.740 0.600 ;
        RECT  2.850 2.620 3.550 2.780 ;
        RECT  2.770 0.440 3.060 1.040 ;
        RECT  2.560 2.350 2.850 3.160 ;
        RECT  1.370 0.710 2.770 0.870 ;
        RECT  1.370 2.350 2.560 2.510 ;
        RECT  2.310 1.030 2.370 1.420 ;
        RECT  2.090 1.030 2.310 2.190 ;
        RECT  2.010 1.910 2.090 2.190 ;
        RECT  1.330 0.710 1.370 2.510 ;
        RECT  1.210 0.710 1.330 2.950 ;
        RECT  1.050 0.970 1.210 1.250 ;
        RECT  1.050 2.120 1.210 2.950 ;
        RECT  0.370 1.090 1.050 1.250 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 0.970 0.370 1.250 ;
        RECT  0.090 2.120 0.370 2.950 ;
    END
END XNOR2X4TR

MACRO XNOR2X2TR
    CLASS CORE ;
    FOREIGN XNOR2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.990 0.840 5.120 2.890 ;
        RECT  4.830 0.550 4.990 2.890 ;
        RECT  4.150 0.550 4.830 0.710 ;
        RECT  3.990 0.550 4.150 2.780 ;
        RECT  3.870 0.550 3.990 0.930 ;
        RECT  3.870 2.130 3.990 2.780 ;
        RECT  3.230 0.550 3.870 0.710 ;
        RECT  3.070 0.550 3.230 2.410 ;
        RECT  2.910 0.870 3.070 1.150 ;
        RECT  2.910 2.130 3.070 2.410 ;
        END
        ANTENNADIFFAREA 6.66 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.360 1.030 1.640 ;
        RECT  0.480 1.240 0.760 1.640 ;
        RECT  0.450 1.410 0.480 1.640 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.240 2.430 1.640 ;
        END
        ANTENNAGATEAREA 0.4464 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 -0.280 5.200 0.280 ;
        RECT  2.030 -0.280 2.310 0.400 ;
        RECT  1.270 -0.280 2.030 0.340 ;
        RECT  0.990 -0.280 1.270 0.400 ;
        RECT  0.410 -0.280 0.990 0.280 ;
        RECT  0.090 -0.280 0.410 1.050 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 3.320 5.200 3.880 ;
        RECT  0.990 3.260 2.410 3.880 ;
        RECT  0.410 3.320 0.990 3.880 ;
        RECT  0.090 1.990 0.410 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.510 0.870 4.630 1.150 ;
        RECT  4.510 2.130 4.630 2.890 ;
        RECT  4.350 0.870 4.510 3.100 ;
        RECT  1.350 2.940 4.350 3.100 ;
        RECT  3.510 0.870 3.670 2.780 ;
        RECT  3.390 0.870 3.510 1.150 ;
        RECT  3.390 2.130 3.510 2.780 ;
        RECT  1.830 2.620 3.390 2.780 ;
        RECT  2.750 1.540 2.910 1.820 ;
        RECT  2.590 0.800 2.750 2.220 ;
        RECT  2.430 0.800 2.590 1.080 ;
        RECT  2.430 1.940 2.590 2.220 ;
        RECT  1.670 0.920 1.830 2.780 ;
        RECT  1.510 0.920 1.670 1.200 ;
        RECT  1.510 1.910 1.670 2.780 ;
        RECT  1.350 1.360 1.510 1.640 ;
        RECT  1.190 0.920 1.350 3.100 ;
        RECT  0.870 0.920 1.190 1.080 ;
        RECT  0.870 2.940 1.190 3.100 ;
        RECT  0.590 0.800 0.870 1.080 ;
        RECT  0.670 1.910 0.870 3.100 ;
        RECT  0.590 1.910 0.670 2.690 ;
    END
END XNOR2X2TR

MACRO XNOR2X1TR
    CLASS CORE ;
    FOREIGN XNOR2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.940 2.090 2.850 ;
        RECT  1.890 0.940 1.930 1.100 ;
        RECT  1.680 2.600 1.930 3.160 ;
        RECT  1.610 0.820 1.890 1.100 ;
        RECT  1.590 2.600 1.680 2.880 ;
        END
        ANTENNADIFFAREA 2.602 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.900 1.070 2.120 ;
        RECT  0.480 1.640 0.760 2.120 ;
        END
        ANTENNAGATEAREA 0.1536 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.840 1.160 3.160 ;
        RECT  0.500 3.000 0.880 3.160 ;
        END
        ANTENNAGATEAREA 0.2232 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.050 -0.280 3.200 0.280 ;
        RECT  2.770 -0.280 3.050 0.400 ;
        RECT  0.930 -0.280 2.770 0.340 ;
        RECT  0.650 -0.280 0.930 1.030 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.010 3.320 3.200 3.880 ;
        RECT  2.730 2.100 3.010 3.880 ;
        RECT  0.340 3.320 2.730 3.880 ;
        RECT  0.710 2.510 0.950 2.680 ;
        RECT  0.520 2.510 0.710 2.770 ;
        RECT  0.340 2.610 0.520 2.770 ;
        RECT  0.160 2.610 0.340 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 1.360 2.970 1.640 ;
        RECT  2.690 0.560 2.850 1.640 ;
        RECT  2.210 0.560 2.690 0.720 ;
        RECT  2.250 1.030 2.530 2.880 ;
        RECT  2.050 0.500 2.210 0.720 ;
        RECT  1.450 0.500 2.050 0.660 ;
        RECT  1.610 1.260 1.770 2.440 ;
        RECT  1.450 1.260 1.610 1.420 ;
        RECT  1.390 2.280 1.610 2.440 ;
        RECT  1.290 0.500 1.450 1.420 ;
        RECT  1.230 1.580 1.450 1.900 ;
        RECT  1.170 2.280 1.390 2.590 ;
        RECT  1.130 0.750 1.290 1.030 ;
        RECT  1.080 1.580 1.230 1.740 ;
        RECT  0.920 1.320 1.080 1.740 ;
        RECT  0.370 1.320 0.920 1.480 ;
        RECT  0.320 1.030 0.370 1.480 ;
        RECT  0.160 1.030 0.320 2.450 ;
        RECT  0.090 1.030 0.160 1.310 ;
        RECT  0.100 2.170 0.160 2.450 ;
    END
END XNOR2X1TR

MACRO TLATSRXLTR
    CLASS CORE ;
    FOREIGN TLATSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.350 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.540 2.380 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.590 0.840 6.720 1.960 ;
        RECT  6.430 0.840 6.590 2.280 ;
        RECT  6.150 2.120 6.430 2.280 ;
        RECT  5.870 2.120 6.150 2.400 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.990 2.580 6.110 2.860 ;
        RECT  5.830 2.560 5.990 2.860 ;
        RECT  5.830 1.640 5.960 1.960 ;
        RECT  5.710 0.970 5.830 1.960 ;
        RECT  5.710 2.560 5.830 2.720 ;
        RECT  5.550 0.970 5.710 2.720 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.970 1.470 4.250 1.750 ;
        RECT  3.960 1.470 3.970 1.630 ;
        RECT  3.680 1.240 3.960 1.630 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.720 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.470 -0.280 6.800 0.280 ;
        RECT  6.190 -0.280 6.470 0.400 ;
        RECT  5.170 -0.280 6.190 0.280 ;
        RECT  4.890 -0.280 5.170 0.400 ;
        RECT  4.050 -0.280 4.890 0.280 ;
        RECT  3.770 -0.280 4.050 0.400 ;
        RECT  1.850 -0.280 3.770 0.280 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  0.370 -0.280 1.570 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.700 3.320 6.800 3.880 ;
        RECT  6.420 2.440 6.700 3.880 ;
        RECT  5.590 3.320 6.420 3.880 ;
        RECT  5.310 2.880 5.590 3.880 ;
        RECT  4.370 3.260 5.310 3.880 ;
        RECT  4.090 3.200 4.370 3.880 ;
        RECT  2.290 3.320 4.090 3.880 ;
        RECT  2.010 3.200 2.290 3.880 ;
        RECT  0.370 3.320 2.010 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 1.170 6.270 1.450 ;
        RECT  5.990 0.630 6.150 1.450 ;
        RECT  5.830 0.630 5.990 0.790 ;
        RECT  5.550 0.490 5.830 0.790 ;
        RECT  5.390 0.630 5.550 0.790 ;
        RECT  5.230 0.630 5.390 2.510 ;
        RECT  5.150 2.350 5.230 2.510 ;
        RECT  4.990 2.350 5.150 3.040 ;
        RECT  4.850 0.710 5.010 2.190 ;
        RECT  3.930 2.820 4.990 3.040 ;
        RECT  4.610 0.710 4.850 0.870 ;
        RECT  4.550 2.350 4.830 2.660 ;
        RECT  4.610 1.510 4.690 1.790 ;
        RECT  4.330 0.570 4.610 0.870 ;
        RECT  4.570 1.030 4.610 1.790 ;
        RECT  4.410 1.030 4.570 2.190 ;
        RECT  1.130 2.440 4.550 2.660 ;
        RECT  4.330 1.030 4.410 1.310 ;
        RECT  4.380 1.910 4.410 2.190 ;
        RECT  4.220 1.910 4.380 2.280 ;
        RECT  3.520 0.710 4.330 0.870 ;
        RECT  2.850 2.120 4.220 2.280 ;
        RECT  3.650 2.820 3.930 3.100 ;
        RECT  3.360 0.710 3.520 1.960 ;
        RECT  3.010 1.680 3.360 1.960 ;
        RECT  3.040 0.480 3.200 1.520 ;
        RECT  2.900 0.480 3.040 0.760 ;
        RECT  2.850 1.360 3.040 1.520 ;
        RECT  2.660 0.920 2.880 1.200 ;
        RECT  2.690 1.360 2.850 2.280 ;
        RECT  2.530 2.880 2.810 3.160 ;
        RECT  1.510 2.120 2.690 2.280 ;
        RECT  1.270 0.920 2.660 1.080 ;
        RECT  0.750 2.880 2.530 3.040 ;
        RECT  1.290 1.700 1.510 2.280 ;
        RECT  1.130 0.480 1.410 0.760 ;
        RECT  1.130 0.920 1.270 1.230 ;
        RECT  0.810 0.600 1.130 0.760 ;
        RECT  0.990 0.920 1.130 2.660 ;
        RECT  0.970 1.070 0.990 2.660 ;
        RECT  0.910 2.380 0.970 2.660 ;
        RECT  0.690 0.600 0.810 1.310 ;
        RECT  0.750 1.910 0.810 2.190 ;
        RECT  0.690 1.910 0.750 3.040 ;
        RECT  0.530 0.600 0.690 3.040 ;
    END
END TLATSRXLTR

MACRO TLATSRX4TR
    CLASS CORE ;
    FOREIGN TLATSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.610 0.530 1.890 ;
        RECT  0.320 1.610 0.360 2.360 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.190 6.320 1.630 ;
        END
        ANTENNAGATEAREA 0.432 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.310 0.440 10.630 2.190 ;
        RECT  10.080 1.440 10.310 2.190 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.390 0.440 9.670 2.190 ;
        RECT  9.280 1.310 9.390 2.190 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.360 7.210 1.640 ;
        RECT  6.480 0.840 6.760 1.640 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 1.500 4.380 1.720 ;
        RECT  3.200 1.500 3.360 1.840 ;
        RECT  2.360 1.680 3.200 1.840 ;
        RECT  2.040 1.240 2.360 1.840 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 -0.280 11.200 0.280 ;
        RECT  10.830 -0.280 11.110 1.310 ;
        RECT  10.150 -0.280 10.830 0.280 ;
        RECT  9.870 -0.280 10.150 1.280 ;
        RECT  9.190 -0.280 9.870 0.280 ;
        RECT  8.910 -0.280 9.190 0.760 ;
        RECT  8.330 -0.280 8.910 0.340 ;
        RECT  8.050 -0.280 8.330 0.360 ;
        RECT  6.970 -0.280 8.050 0.280 ;
        RECT  6.690 -0.280 6.970 0.360 ;
        RECT  4.400 -0.280 6.690 0.280 ;
        RECT  4.120 -0.280 4.400 0.640 ;
        RECT  2.080 -0.280 4.120 0.280 ;
        RECT  1.800 -0.280 2.080 0.400 ;
        RECT  0.850 -0.280 1.800 0.280 ;
        RECT  0.570 -0.280 0.850 0.710 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 3.320 11.200 3.880 ;
        RECT  10.830 2.910 11.110 3.880 ;
        RECT  10.150 3.320 10.830 3.880 ;
        RECT  9.870 2.910 10.150 3.880 ;
        RECT  9.150 3.320 9.870 3.880 ;
        RECT  8.870 3.200 9.150 3.880 ;
        RECT  8.330 3.320 8.870 3.880 ;
        RECT  8.050 3.200 8.330 3.880 ;
        RECT  6.970 3.260 8.050 3.880 ;
        RECT  6.810 3.200 6.970 3.880 ;
        RECT  4.900 3.320 6.810 3.880 ;
        RECT  4.620 2.900 4.900 3.880 ;
        RECT  2.610 3.320 4.620 3.880 ;
        RECT  2.330 3.020 2.610 3.880 ;
        RECT  0.890 3.320 2.330 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.790 1.580 11.070 2.750 ;
        RECT  8.980 2.590 10.790 2.750 ;
        RECT  8.820 1.030 8.980 2.750 ;
        RECT  8.570 1.030 8.820 1.310 ;
        RECT  8.730 1.910 8.820 2.750 ;
        RECT  8.570 1.910 8.730 3.040 ;
        RECT  8.410 1.470 8.650 1.750 ;
        RECT  6.650 2.880 8.570 3.040 ;
        RECT  8.370 1.470 8.410 2.720 ;
        RECT  8.250 1.590 8.370 2.720 ;
        RECT  5.700 2.560 8.250 2.720 ;
        RECT  7.930 0.520 8.090 2.280 ;
        RECT  7.870 0.520 7.930 0.680 ;
        RECT  7.650 2.120 7.930 2.400 ;
        RECT  7.590 0.460 7.870 0.680 ;
        RECT  7.490 0.920 7.770 1.960 ;
        RECT  5.920 0.520 7.590 0.680 ;
        RECT  7.210 0.920 7.490 1.200 ;
        RECT  7.470 1.800 7.490 1.960 ;
        RECT  7.190 1.800 7.470 2.190 ;
        RECT  5.920 1.800 7.190 2.100 ;
        RECT  6.370 2.880 6.650 3.120 ;
        RECT  5.220 2.940 6.200 3.160 ;
        RECT  5.760 0.520 5.920 1.070 ;
        RECT  5.640 1.250 5.920 2.100 ;
        RECT  5.360 0.910 5.760 1.070 ;
        RECT  5.580 2.500 5.700 2.780 ;
        RECT  3.680 1.880 5.640 2.100 ;
        RECT  4.720 0.470 5.600 0.750 ;
        RECT  5.420 2.260 5.580 2.780 ;
        RECT  4.100 2.260 5.420 2.420 ;
        RECT  5.200 0.910 5.360 1.520 ;
        RECT  5.060 2.580 5.220 3.160 ;
        RECT  5.080 1.180 5.200 1.520 ;
        RECT  3.040 1.180 5.080 1.340 ;
        RECT  4.420 2.580 5.060 2.740 ;
        RECT  4.560 0.470 4.720 1.020 ;
        RECT  1.410 0.800 4.560 1.020 ;
        RECT  4.260 2.580 4.420 2.860 ;
        RECT  1.240 2.700 4.260 2.860 ;
        RECT  3.940 2.260 4.100 2.540 ;
        RECT  1.450 2.320 3.940 2.540 ;
        RECT  3.520 1.880 3.680 2.160 ;
        RECT  1.770 2.000 3.520 2.160 ;
        RECT  2.760 1.180 3.040 1.520 ;
        RECT  1.610 1.240 1.770 2.160 ;
        RECT  1.450 1.240 1.610 1.520 ;
        RECT  1.290 1.910 1.450 2.540 ;
        RECT  1.290 0.440 1.410 1.080 ;
        RECT  1.130 0.440 1.290 2.540 ;
        RECT  0.970 2.700 1.240 3.040 ;
        RECT  0.810 0.920 0.970 3.040 ;
        RECT  0.690 0.920 0.810 2.680 ;
        RECT  0.370 0.920 0.690 1.080 ;
        RECT  0.370 2.520 0.690 2.680 ;
        RECT  0.090 0.440 0.370 1.080 ;
        RECT  0.090 2.520 0.370 3.160 ;
    END
END TLATSRX4TR

MACRO TLATSRX2TR
    CLASS CORE ;
    FOREIGN TLATSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.400 2.760 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.640 2.760 1.960 ;
        RECT  2.440 1.640 2.640 2.020 ;
        RECT  2.360 1.740 2.440 2.020 ;
        END
        ANTENNAGATEAREA 0.2208 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 0.440 7.520 3.160 ;
        RECT  7.230 1.910 7.280 3.160 ;
        END
        ANTENNADIFFAREA 3.47 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.640 6.720 1.960 ;
        RECT  6.490 1.640 6.530 2.190 ;
        RECT  6.270 1.020 6.490 2.190 ;
        RECT  6.190 1.020 6.270 1.300 ;
        END
        ANTENNADIFFAREA 2.516 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.040 1.580 4.560 1.960 ;
        END
        ANTENNAGATEAREA 0.084 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.620 2.160 1.960 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.990 -0.280 7.600 0.280 ;
        RECT  6.710 -0.280 6.990 0.400 ;
        RECT  5.610 -0.280 6.710 0.280 ;
        RECT  5.330 -0.280 5.610 0.400 ;
        RECT  4.360 -0.280 5.330 0.280 ;
        RECT  4.080 -0.280 4.360 0.400 ;
        RECT  2.080 -0.280 4.080 0.280 ;
        RECT  1.800 -0.280 2.080 0.800 ;
        RECT  0.400 -0.280 1.800 0.340 ;
        RECT  0.090 -0.280 0.400 0.970 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.030 3.320 7.600 3.880 ;
        RECT  6.750 2.910 7.030 3.880 ;
        RECT  2.400 3.320 6.750 3.880 ;
        RECT  2.120 3.200 2.400 3.880 ;
        RECT  0.370 3.320 2.120 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.040 1.460 7.120 1.740 ;
        RECT  6.880 0.570 7.040 2.700 ;
        RECT  6.130 0.570 6.880 0.730 ;
        RECT  6.210 2.540 6.880 2.700 ;
        RECT  6.110 2.370 6.210 2.700 ;
        RECT  5.850 0.450 6.130 0.730 ;
        RECT  5.930 2.370 6.110 3.160 ;
        RECT  5.770 1.530 6.010 1.810 ;
        RECT  4.240 3.000 5.930 3.160 ;
        RECT  5.610 1.530 5.770 2.840 ;
        RECT  4.560 2.680 5.610 2.840 ;
        RECT  5.290 0.580 5.450 2.060 ;
        RECT  4.920 0.580 5.290 0.740 ;
        RECT  5.040 1.780 5.290 2.060 ;
        RECT  4.880 1.300 5.130 1.580 ;
        RECT  4.880 2.240 5.000 2.520 ;
        RECT  4.640 0.440 4.920 0.740 ;
        RECT  4.720 0.900 4.880 2.520 ;
        RECT  4.600 0.900 4.720 1.180 ;
        RECT  3.080 2.180 4.720 2.340 ;
        RECT  3.880 0.580 4.640 0.740 ;
        RECT  4.400 2.500 4.560 2.840 ;
        RECT  1.240 2.500 4.400 2.720 ;
        RECT  3.960 2.880 4.240 3.160 ;
        RECT  3.720 0.580 3.880 2.020 ;
        RECT  3.240 1.740 3.720 2.020 ;
        RECT  3.400 0.540 3.560 1.580 ;
        RECT  3.150 2.880 3.450 3.160 ;
        RECT  3.200 0.540 3.400 0.820 ;
        RECT  3.080 1.420 3.400 1.580 ;
        RECT  2.960 0.980 3.240 1.260 ;
        RECT  1.620 2.880 3.150 3.040 ;
        RECT  2.920 1.420 3.080 2.340 ;
        RECT  1.560 0.980 2.960 1.230 ;
        RECT  1.480 2.180 2.920 2.340 ;
        RECT  0.850 0.560 1.640 0.780 ;
        RECT  1.430 2.880 1.620 3.150 ;
        RECT  1.280 0.950 1.560 1.230 ;
        RECT  1.320 1.390 1.480 2.340 ;
        RECT  0.720 2.990 1.430 3.150 ;
        RECT  1.220 1.390 1.320 1.670 ;
        RECT  1.060 1.070 1.280 1.230 ;
        RECT  1.160 2.500 1.240 2.830 ;
        RECT  1.060 1.830 1.160 2.830 ;
        RECT  1.000 1.070 1.060 2.830 ;
        RECT  0.900 1.070 1.000 1.990 ;
        RECT  0.960 2.550 1.000 2.830 ;
        RECT  0.720 0.560 0.850 0.910 ;
        RECT  0.720 2.150 0.840 2.370 ;
        RECT  0.560 0.560 0.720 3.150 ;
    END
END TLATSRX2TR

MACRO TLATSRX1TR
    CLASS CORE ;
    FOREIGN TLATSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.370 1.670 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.630 2.470 1.960 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.640 0.640 6.760 1.200 ;
        RECT  6.480 0.640 6.640 2.280 ;
        RECT  6.380 2.120 6.480 2.280 ;
        RECT  6.100 2.120 6.380 2.400 ;
        END
        ANTENNADIFFAREA 1.724 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 2.630 6.320 3.010 ;
        RECT  5.940 2.630 6.040 2.790 ;
        RECT  5.880 1.640 5.940 2.790 ;
        RECT  5.780 0.980 5.880 2.790 ;
        RECT  5.600 0.980 5.780 1.970 ;
        END
        ANTENNADIFFAREA 1.568 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.070 1.240 4.360 1.680 ;
        RECT  4.040 1.240 4.070 1.560 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.750 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.590 -0.280 7.200 0.280 ;
        RECT  6.310 -0.280 6.590 0.400 ;
        RECT  5.360 -0.280 6.310 0.280 ;
        RECT  5.080 -0.280 5.360 0.400 ;
        RECT  4.110 -0.280 5.080 0.280 ;
        RECT  3.830 -0.280 4.110 0.400 ;
        RECT  1.950 -0.280 3.830 0.280 ;
        RECT  1.670 -0.280 1.950 0.400 ;
        RECT  0.370 -0.280 1.670 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.900 3.320 7.200 3.880 ;
        RECT  6.620 2.600 6.900 3.880 ;
        RECT  5.620 3.320 6.620 3.880 ;
        RECT  5.340 2.930 5.620 3.880 ;
        RECT  4.430 3.260 5.340 3.880 ;
        RECT  4.150 3.200 4.430 3.880 ;
        RECT  2.350 3.320 4.150 3.880 ;
        RECT  2.070 3.200 2.350 3.880 ;
        RECT  0.370 3.320 2.070 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.200 0.970 6.320 1.250 ;
        RECT  6.040 0.660 6.200 1.250 ;
        RECT  5.920 0.660 6.040 0.820 ;
        RECT  5.640 0.440 5.920 0.820 ;
        RECT  5.440 0.660 5.640 0.820 ;
        RECT  5.280 0.660 5.440 2.600 ;
        RECT  5.180 2.440 5.280 2.600 ;
        RECT  5.020 2.440 5.180 3.040 ;
        RECT  4.960 0.590 5.120 2.280 ;
        RECT  4.810 2.820 5.020 3.040 ;
        RECT  4.800 0.590 4.960 0.750 ;
        RECT  4.840 2.000 4.960 2.280 ;
        RECT  3.070 2.440 4.860 2.660 ;
        RECT  3.990 2.880 4.810 3.040 ;
        RECT  4.520 0.450 4.800 0.750 ;
        RECT  4.680 0.910 4.800 1.840 ;
        RECT  4.520 0.910 4.680 2.280 ;
        RECT  3.630 0.590 4.520 0.750 ;
        RECT  4.350 1.990 4.520 2.280 ;
        RECT  2.830 2.120 4.350 2.280 ;
        RECT  3.710 2.880 3.990 3.160 ;
        RECT  3.470 0.590 3.630 1.820 ;
        RECT  3.270 1.660 3.470 1.820 ;
        RECT  3.150 0.440 3.310 1.500 ;
        RECT  2.990 1.660 3.270 1.940 ;
        RECT  2.950 0.440 3.150 0.720 ;
        RECT  2.830 1.340 3.150 1.500 ;
        RECT  1.190 2.440 3.070 2.720 ;
        RECT  2.710 0.900 2.990 1.180 ;
        RECT  2.590 2.880 2.870 3.160 ;
        RECT  2.670 1.340 2.830 2.280 ;
        RECT  1.270 0.900 2.710 1.060 ;
        RECT  1.510 2.120 2.670 2.280 ;
        RECT  1.550 2.880 2.590 3.040 ;
        RECT  1.350 2.880 1.550 3.160 ;
        RECT  1.230 0.460 1.510 0.740 ;
        RECT  1.290 1.580 1.510 2.280 ;
        RECT  0.750 3.000 1.350 3.160 ;
        RECT  1.130 0.900 1.270 1.190 ;
        RECT  0.810 0.580 1.230 0.740 ;
        RECT  1.130 2.440 1.190 2.840 ;
        RECT  0.990 0.900 1.130 2.840 ;
        RECT  0.970 1.030 0.990 2.840 ;
        RECT  0.910 2.560 0.970 2.840 ;
        RECT  0.690 0.580 0.810 1.250 ;
        RECT  0.750 1.870 0.810 2.220 ;
        RECT  0.690 1.870 0.750 3.160 ;
        RECT  0.530 0.580 0.690 3.160 ;
    END
END TLATSRX1TR

MACRO TLATNTSCAX8TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.540 3.040 1.960 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.420 0.440 16.700 3.160 ;
        RECT  16.240 0.440 16.420 2.960 ;
        RECT  11.300 0.440 16.240 0.840 ;
        RECT  15.880 2.080 16.240 2.960 ;
        RECT  15.020 2.080 15.880 2.560 ;
        RECT  14.740 2.080 15.020 3.160 ;
        RECT  13.420 2.080 14.740 2.560 ;
        RECT  13.140 2.080 13.420 3.160 ;
        RECT  11.820 2.080 13.140 2.560 ;
        RECT  11.540 2.080 11.820 3.160 ;
        END
        ANTENNADIFFAREA 12.596 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.240 3.560 1.710 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.520 1.500 1.800 ;
        RECT  0.480 1.520 0.760 1.960 ;
        RECT  0.420 1.520 0.480 1.800 ;
        END
        ANTENNAGATEAREA 0.7992 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.980 -0.280 16.800 0.280 ;
        RECT  10.700 -0.280 10.980 0.400 ;
        RECT  8.540 -0.280 10.700 0.340 ;
        RECT  8.260 -0.280 8.540 0.790 ;
        RECT  6.480 -0.280 8.260 0.280 ;
        RECT  6.200 -0.280 6.480 0.930 ;
        RECT  4.840 -0.280 6.200 0.280 ;
        RECT  4.560 -0.280 4.840 0.380 ;
        RECT  3.800 -0.280 4.560 0.280 ;
        RECT  3.520 -0.280 3.800 0.380 ;
        RECT  2.800 -0.280 3.520 0.280 ;
        RECT  2.520 -0.280 2.800 0.380 ;
        RECT  1.820 -0.280 2.520 0.280 ;
        RECT  1.540 -0.280 1.820 0.860 ;
        RECT  0.860 -0.280 1.540 0.280 ;
        RECT  0.580 -0.280 0.860 1.360 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.860 3.320 16.800 3.880 ;
        RECT  15.580 3.180 15.860 3.880 ;
        RECT  14.220 3.320 15.580 3.880 ;
        RECT  13.940 2.930 14.220 3.880 ;
        RECT  12.620 3.320 13.940 3.880 ;
        RECT  12.340 2.930 12.620 3.880 ;
        RECT  10.980 3.320 12.340 3.880 ;
        RECT  10.280 3.180 10.980 3.880 ;
        RECT  8.520 3.320 10.280 3.880 ;
        RECT  8.240 3.260 8.520 3.880 ;
        RECT  6.840 3.320 8.240 3.880 ;
        RECT  6.560 3.260 6.840 3.880 ;
        RECT  5.080 3.320 6.560 3.880 ;
        RECT  4.800 3.260 5.080 3.880 ;
        RECT  4.040 3.320 4.800 3.880 ;
        RECT  3.760 3.260 4.040 3.880 ;
        RECT  2.800 3.320 3.760 3.880 ;
        RECT  2.520 3.260 2.800 3.880 ;
        RECT  1.860 3.320 2.520 3.880 ;
        RECT  1.580 3.260 1.860 3.880 ;
        RECT  0.860 3.320 1.580 3.880 ;
        RECT  0.580 2.930 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.860 1.240 16.080 1.520 ;
        RECT  15.700 1.000 15.860 1.860 ;
        RECT  11.140 1.000 15.700 1.160 ;
        RECT  11.580 1.640 15.700 1.860 ;
        RECT  11.140 1.320 15.540 1.480 ;
        RECT  10.980 0.650 11.140 1.160 ;
        RECT  10.980 1.320 11.140 2.680 ;
        RECT  9.800 0.650 10.980 0.810 ;
        RECT  10.120 2.520 10.980 2.680 ;
        RECT  10.660 1.090 10.820 2.120 ;
        RECT  10.420 1.090 10.660 1.250 ;
        RECT  10.580 1.960 10.660 2.120 ;
        RECT  10.300 1.960 10.580 2.240 ;
        RECT  9.800 1.410 10.500 1.690 ;
        RECT  10.140 0.970 10.420 1.250 ;
        RECT  10.180 2.080 10.300 2.240 ;
        RECT  9.960 2.080 10.180 2.360 ;
        RECT  9.960 2.520 10.120 3.100 ;
        RECT  9.680 2.940 9.960 3.100 ;
        RECT  9.640 0.650 9.800 2.770 ;
        RECT  9.400 2.940 9.680 3.160 ;
        RECT  9.100 0.950 9.640 1.170 ;
        RECT  5.720 2.550 9.640 2.770 ;
        RECT  9.320 1.480 9.480 2.390 ;
        RECT  5.560 2.940 9.400 3.100 ;
        RECT  9.180 1.480 9.320 1.640 ;
        RECT  5.560 2.230 9.320 2.390 ;
        RECT  8.900 1.360 9.180 1.640 ;
        RECT  7.480 1.820 9.160 2.010 ;
        RECT  7.700 0.950 9.100 1.110 ;
        RECT  7.490 1.410 8.900 1.570 ;
        RECT  7.000 0.710 7.700 1.110 ;
        RECT  7.210 1.280 7.490 1.570 ;
        RECT  7.200 1.740 7.480 2.010 ;
        RECT  5.720 1.410 7.210 1.570 ;
        RECT  6.200 1.850 7.200 2.010 ;
        RECT  6.800 0.950 7.000 1.110 ;
        RECT  6.640 0.950 6.800 1.250 ;
        RECT  6.040 1.090 6.640 1.250 ;
        RECT  5.920 1.760 6.200 2.010 ;
        RECT  5.880 1.070 6.040 1.250 ;
        RECT  5.240 1.850 5.920 2.010 ;
        RECT  5.680 1.070 5.880 1.230 ;
        RECT  5.440 1.390 5.720 1.580 ;
        RECT  5.400 0.950 5.680 1.230 ;
        RECT  5.400 2.230 5.560 3.100 ;
        RECT  1.340 2.940 5.400 3.100 ;
        RECT  5.080 0.540 5.240 2.780 ;
        RECT  2.380 0.540 5.080 0.700 ;
        RECT  2.280 2.620 5.080 2.780 ;
        RECT  4.800 1.410 4.920 1.690 ;
        RECT  4.640 1.150 4.800 2.450 ;
        RECT  4.320 1.150 4.640 1.310 ;
        RECT  4.280 2.170 4.640 2.450 ;
        RECT  3.880 1.730 4.480 2.010 ;
        RECT  4.040 1.030 4.320 1.310 ;
        RECT  3.720 0.860 3.880 2.240 ;
        RECT  3.040 0.860 3.720 1.080 ;
        RECT  3.360 1.960 3.720 2.240 ;
        RECT  2.280 0.540 2.380 1.360 ;
        RECT  2.100 0.540 2.280 2.780 ;
        RECT  2.000 1.960 2.100 2.780 ;
        RECT  1.820 1.410 1.940 1.690 ;
        RECT  1.660 1.200 1.820 2.120 ;
        RECT  1.340 1.200 1.660 1.360 ;
        RECT  1.340 1.960 1.660 2.120 ;
        RECT  1.060 0.440 1.340 1.360 ;
        RECT  1.060 1.960 1.340 3.100 ;
        RECT  0.380 2.120 1.060 2.280 ;
        RECT  0.260 0.500 0.380 1.360 ;
        RECT  0.320 2.120 0.380 3.160 ;
        RECT  0.260 1.960 0.320 3.160 ;
        RECT  0.100 0.500 0.260 3.160 ;
    END
END TLATNTSCAX8TR

MACRO TLATNTSCAX6TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 1.320 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.390 0.500 10.650 2.280 ;
        RECT  10.290 0.500 10.390 3.160 ;
        RECT  8.270 0.500 10.290 0.790 ;
        RECT  10.110 1.910 10.290 3.160 ;
        RECT  8.920 1.910 10.110 2.270 ;
        RECT  8.280 1.910 8.920 3.130 ;
        END
        ANTENNADIFFAREA 6.4005 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.640 2.870 1.970 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.520 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.110 -0.280 10.800 0.280 ;
        RECT  9.830 -0.280 10.110 0.340 ;
        RECT  9.070 -0.280 9.830 0.280 ;
        RECT  8.790 -0.280 9.070 0.340 ;
        RECT  8.020 -0.280 8.790 0.280 ;
        RECT  7.170 -0.280 8.020 0.340 ;
        RECT  5.610 -0.280 7.170 0.280 ;
        RECT  5.330 -0.280 5.610 0.340 ;
        RECT  3.040 -0.280 5.330 0.280 ;
        RECT  2.760 -0.280 3.040 0.330 ;
        RECT  1.410 -0.280 2.760 0.280 ;
        RECT  1.130 -0.280 1.410 0.340 ;
        RECT  0.410 -0.280 1.130 0.280 ;
        RECT  0.140 -0.280 0.410 1.200 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.620 3.320 10.800 3.880 ;
        RECT  9.270 2.510 9.620 3.880 ;
        RECT  7.950 3.320 9.270 3.880 ;
        RECT  7.670 2.820 7.950 3.880 ;
        RECT  5.730 3.320 7.670 3.880 ;
        RECT  5.450 3.260 5.730 3.880 ;
        RECT  4.050 3.320 5.450 3.880 ;
        RECT  3.770 2.710 4.050 3.880 ;
        RECT  1.770 3.320 3.770 3.880 ;
        RECT  1.080 2.930 1.770 3.880 ;
        RECT  0.410 3.320 1.080 3.880 ;
        RECT  0.140 2.120 0.410 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.110 1.470 10.130 1.750 ;
        RECT  9.950 0.950 10.110 1.750 ;
        RECT  8.110 0.950 9.950 1.110 ;
        RECT  8.550 1.590 9.950 1.750 ;
        RECT  8.190 1.270 9.790 1.430 ;
        RECT  8.120 1.270 8.190 1.560 ;
        RECT  7.960 1.270 8.120 2.450 ;
        RECT  7.950 0.650 8.110 1.110 ;
        RECT  7.330 2.290 7.960 2.450 ;
        RECT  6.830 0.650 7.950 0.810 ;
        RECT  7.630 0.970 7.790 2.130 ;
        RECT  6.990 0.970 7.630 1.290 ;
        RECT  7.170 1.970 7.630 2.130 ;
        RECT  7.010 1.450 7.470 1.730 ;
        RECT  7.170 2.290 7.330 3.100 ;
        RECT  4.490 2.940 7.170 3.100 ;
        RECT  6.850 1.450 7.010 2.660 ;
        RECT  6.830 1.450 6.850 1.610 ;
        RECT  4.830 2.500 6.850 2.660 ;
        RECT  6.670 0.650 6.830 1.610 ;
        RECT  6.510 1.770 6.690 2.010 ;
        RECT  6.170 0.650 6.670 0.930 ;
        RECT  6.350 1.090 6.510 2.010 ;
        RECT  4.330 1.090 6.350 1.250 ;
        RECT  5.150 1.850 6.350 2.010 ;
        RECT  6.030 1.410 6.190 1.690 ;
        RECT  4.490 0.770 6.170 0.930 ;
        RECT  4.490 1.440 6.030 1.600 ;
        RECT  4.990 1.760 5.150 2.010 ;
        RECT  4.810 1.760 4.990 1.920 ;
        RECT  4.670 2.270 4.830 2.660 ;
        RECT  4.330 1.440 4.490 3.100 ;
        RECT  4.170 0.500 4.330 1.250 ;
        RECT  3.510 2.390 4.330 2.550 ;
        RECT  1.900 0.500 4.170 0.660 ;
        RECT  4.010 1.420 4.170 1.580 ;
        RECT  3.850 1.000 4.010 1.900 ;
        RECT  3.470 1.000 3.850 1.160 ;
        RECT  3.510 1.740 3.850 1.900 ;
        RECT  3.190 1.320 3.690 1.580 ;
        RECT  3.350 1.740 3.510 2.190 ;
        RECT  3.350 2.390 3.510 2.680 ;
        RECT  3.310 0.880 3.470 1.160 ;
        RECT  1.150 2.520 3.350 2.680 ;
        RECT  3.030 1.320 3.190 2.290 ;
        RECT  2.640 1.320 3.030 1.480 ;
        RECT  2.550 2.130 3.030 2.290 ;
        RECT  2.480 0.820 2.640 1.480 ;
        RECT  2.180 0.820 2.480 0.980 ;
        RECT  1.780 0.500 1.900 1.130 ;
        RECT  1.740 0.500 1.780 2.130 ;
        RECT  1.620 0.970 1.740 2.130 ;
        RECT  1.310 1.970 1.620 2.130 ;
        RECT  1.150 1.460 1.460 1.740 ;
        RECT  0.990 1.040 1.150 2.680 ;
        RECT  0.890 1.040 0.990 1.200 ;
        RECT  0.880 2.380 0.990 2.680 ;
        RECT  0.600 0.510 0.890 1.200 ;
        RECT  0.620 2.380 0.880 3.160 ;
    END
END TLATNTSCAX6TR

MACRO TLATNTSCAX4TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.320 1.960 1.960 ;
        RECT  1.640 1.640 1.670 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 1.840 7.520 2.670 ;
        RECT  6.970 1.050 7.210 2.670 ;
        RECT  6.890 1.050 6.970 1.330 ;
        END
        ANTENNADIFFAREA 4.228 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 2.430 2.360 2.760 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.430 2.760 ;
        END
        ANTENNAGATEAREA 0.2736 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.850 -0.280 8.400 0.280 ;
        RECT  7.690 -0.280 7.850 1.260 ;
        RECT  6.650 -0.280 7.690 0.280 ;
        RECT  4.650 -0.280 6.650 0.340 ;
        RECT  3.250 -0.280 4.650 0.280 ;
        RECT  2.470 -0.280 3.250 0.400 ;
        RECT  0.850 -0.280 2.470 0.280 ;
        RECT  0.570 -0.280 0.850 0.800 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.310 3.320 8.400 3.880 ;
        RECT  8.030 2.190 8.310 3.880 ;
        RECT  6.670 3.320 8.030 3.880 ;
        RECT  4.650 3.260 6.670 3.880 ;
        RECT  3.250 3.320 4.650 3.880 ;
        RECT  1.140 3.260 3.250 3.880 ;
        RECT  0.370 3.320 1.140 3.880 ;
        RECT  0.090 2.920 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.890 1.600 8.050 2.030 ;
        RECT  7.870 1.870 7.890 2.030 ;
        RECT  7.710 1.870 7.870 3.100 ;
        RECT  6.810 2.940 7.710 3.100 ;
        RECT  7.530 1.520 7.670 1.680 ;
        RECT  7.370 0.500 7.530 1.680 ;
        RECT  5.750 0.500 7.370 0.660 ;
        RECT  6.650 1.600 6.810 3.100 ;
        RECT  3.710 2.820 6.650 3.100 ;
        RECT  6.330 1.110 6.490 2.090 ;
        RECT  5.910 1.110 6.330 1.270 ;
        RECT  6.210 1.930 6.330 2.090 ;
        RECT  5.930 1.930 6.210 2.210 ;
        RECT  5.750 1.460 6.170 1.740 ;
        RECT  5.810 1.930 5.930 2.120 ;
        RECT  5.530 1.900 5.810 2.120 ;
        RECT  5.590 0.500 5.750 1.740 ;
        RECT  5.270 0.500 5.590 0.660 ;
        RECT  5.270 1.580 5.590 1.740 ;
        RECT  4.290 1.090 5.430 1.370 ;
        RECT  4.990 0.500 5.270 0.930 ;
        RECT  5.110 1.580 5.270 2.660 ;
        RECT  4.990 2.140 5.110 2.660 ;
        RECT  3.810 0.500 4.990 0.780 ;
        RECT  4.090 2.140 4.990 2.300 ;
        RECT  4.130 0.940 4.290 1.900 ;
        RECT  3.650 0.940 4.130 1.100 ;
        RECT  4.070 1.620 4.130 1.900 ;
        RECT  3.870 2.140 4.090 2.420 ;
        RECT  3.710 1.260 3.890 1.540 ;
        RECT  3.550 1.260 3.710 3.100 ;
        RECT  3.490 0.560 3.650 1.100 ;
        RECT  0.870 2.940 3.550 3.100 ;
        RECT  1.510 0.560 3.490 0.720 ;
        RECT  3.330 1.380 3.390 1.660 ;
        RECT  3.170 1.170 3.330 2.300 ;
        RECT  2.850 1.170 3.170 1.330 ;
        RECT  2.850 2.140 3.170 2.300 ;
        RECT  2.470 1.700 3.010 1.980 ;
        RECT  2.570 1.050 2.850 1.330 ;
        RECT  2.630 2.140 2.850 2.730 ;
        RECT  2.350 1.700 2.470 2.270 ;
        RECT  2.190 0.880 2.350 2.270 ;
        RECT  1.910 0.880 2.190 1.160 ;
        RECT  1.390 0.560 1.510 1.290 ;
        RECT  1.350 0.560 1.390 2.150 ;
        RECT  1.230 1.000 1.350 2.150 ;
        RECT  1.190 1.990 1.230 2.150 ;
        RECT  0.910 1.990 1.190 2.270 ;
        RECT  0.750 1.360 1.070 1.640 ;
        RECT  0.750 2.880 0.870 3.160 ;
        RECT  0.590 1.150 0.750 3.160 ;
        RECT  0.370 1.150 0.590 1.310 ;
        RECT  0.090 0.500 0.370 1.310 ;
    END
END TLATNTSCAX4TR

MACRO TLATNTSCAX3TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.260 1.980 1.540 ;
        RECT  1.700 1.260 1.960 1.960 ;
        RECT  1.640 1.640 1.700 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.030 1.960 6.360 2.780 ;
        RECT  5.870 1.030 6.030 2.120 ;
        RECT  5.750 1.030 5.870 1.310 ;
        END
        ANTENNADIFFAREA 3.128 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.440 2.320 2.780 ;
        RECT  2.140 2.370 2.300 2.780 ;
        RECT  2.020 2.370 2.140 2.760 ;
        RECT  2.010 2.370 2.020 2.530 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.850 -0.280 7.200 0.280 ;
        RECT  6.570 -0.280 6.850 1.310 ;
        RECT  5.470 -0.280 6.570 0.340 ;
        RECT  4.760 -0.280 5.470 0.400 ;
        RECT  3.180 -0.280 4.760 0.280 ;
        RECT  2.500 -0.280 3.180 0.340 ;
        RECT  1.500 -0.280 2.500 0.280 ;
        RECT  0.980 -0.280 1.500 0.340 ;
        RECT  0.700 -0.280 0.980 0.860 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.320 7.200 3.880 ;
        RECT  6.890 2.020 7.110 3.880 ;
        RECT  0.450 3.320 6.890 3.880 ;
        RECT  0.160 2.920 0.450 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.730 1.580 6.910 1.860 ;
        RECT  6.570 1.580 6.730 3.140 ;
        RECT  5.710 2.940 6.570 3.140 ;
        RECT  6.190 0.630 6.410 1.800 ;
        RECT  4.580 0.630 6.190 0.790 ;
        RECT  5.490 1.580 5.710 3.140 ;
        RECT  3.500 2.940 5.490 3.140 ;
        RECT  5.170 1.150 5.330 2.070 ;
        RECT  5.030 1.150 5.170 1.310 ;
        RECT  5.040 1.910 5.170 2.070 ;
        RECT  4.960 1.910 5.040 2.190 ;
        RECT  4.750 1.030 5.030 1.310 ;
        RECT  4.580 1.470 5.010 1.750 ;
        RECT  4.740 1.910 4.960 2.590 ;
        RECT  4.420 0.630 4.580 2.540 ;
        RECT  4.060 0.630 4.420 0.790 ;
        RECT  3.940 2.380 4.420 2.540 ;
        RECT  4.040 0.950 4.260 1.870 ;
        RECT  3.780 0.440 4.060 0.790 ;
        RECT  3.620 0.950 4.040 1.110 ;
        RECT  3.660 2.380 3.940 2.660 ;
        RECT  3.740 1.280 3.860 1.560 ;
        RECT  3.580 1.280 3.740 2.220 ;
        RECT  3.460 0.500 3.620 1.110 ;
        RECT  3.500 2.060 3.580 2.220 ;
        RECT  3.340 2.060 3.500 3.140 ;
        RECT  1.540 0.500 3.460 0.660 ;
        RECT  3.300 1.280 3.420 1.560 ;
        RECT  0.860 2.940 3.340 3.140 ;
        RECT  3.140 0.980 3.300 1.900 ;
        RECT  2.540 0.980 3.140 1.140 ;
        RECT  2.820 1.740 3.140 1.900 ;
        RECT  2.500 1.300 2.980 1.580 ;
        RECT  2.660 1.740 2.820 2.780 ;
        RECT  2.480 2.500 2.660 2.780 ;
        RECT  2.340 1.300 2.500 2.210 ;
        RECT  2.300 1.300 2.340 1.460 ;
        RECT  2.220 1.930 2.340 2.210 ;
        RECT  2.140 0.820 2.300 1.460 ;
        RECT  1.940 0.820 2.140 1.100 ;
        RECT  1.420 0.500 1.540 1.300 ;
        RECT  1.380 0.500 1.420 1.950 ;
        RECT  1.260 0.940 1.380 1.950 ;
        RECT  1.240 1.790 1.260 1.950 ;
        RECT  1.020 1.790 1.240 2.210 ;
        RECT  0.860 1.350 1.100 1.630 ;
        RECT  0.700 1.140 0.860 3.140 ;
        RECT  0.500 1.140 0.700 1.300 ;
        RECT  0.160 0.580 0.500 1.300 ;
    END
END TLATNTSCAX3TR

MACRO TLATNTSCAX2TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 1.140 1.920 1.750 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 1.910 6.210 3.160 ;
        RECT  5.840 1.910 5.930 2.360 ;
        RECT  5.680 1.090 5.840 2.360 ;
        RECT  5.510 1.090 5.680 1.250 ;
        END
        ANTENNADIFFAREA 2.764 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.360 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.380 2.760 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.310 -0.280 6.400 0.280 ;
        RECT  6.030 -0.280 6.310 0.340 ;
        RECT  5.270 -0.280 6.030 0.280 ;
        RECT  4.580 -0.280 5.270 0.460 ;
        RECT  3.040 -0.280 4.580 0.280 ;
        RECT  2.480 -0.280 3.040 0.340 ;
        RECT  0.890 -0.280 2.480 0.280 ;
        RECT  0.830 -0.280 0.890 0.340 ;
        RECT  0.670 -0.280 0.830 0.800 ;
        RECT  0.610 -0.280 0.670 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.370 3.320 6.400 3.880 ;
        RECT  5.090 3.260 5.370 3.880 ;
        RECT  3.160 3.320 5.090 3.880 ;
        RECT  2.880 3.250 3.160 3.880 ;
        RECT  1.400 3.320 2.880 3.880 ;
        RECT  1.120 2.800 1.400 3.880 ;
        RECT  0.310 3.320 1.120 3.880 ;
        RECT  0.150 2.930 0.310 3.880 ;
        RECT  0.000 3.320 0.150 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.000 0.710 6.160 1.640 ;
        RECT  4.350 0.710 6.000 0.870 ;
        RECT  5.360 1.580 5.520 3.090 ;
        RECT  4.240 2.930 5.360 3.090 ;
        RECT  5.040 1.150 5.200 2.130 ;
        RECT  4.770 1.150 5.040 1.310 ;
        RECT  4.670 1.970 5.040 2.130 ;
        RECT  4.350 1.470 4.880 1.750 ;
        RECT  4.610 1.030 4.770 1.310 ;
        RECT  4.510 1.970 4.670 2.590 ;
        RECT  4.190 0.710 4.350 2.060 ;
        RECT  3.960 2.930 4.240 3.130 ;
        RECT  3.820 0.710 4.190 0.870 ;
        RECT  3.940 1.900 4.190 2.060 ;
        RECT  3.870 1.030 4.030 1.730 ;
        RECT  3.560 2.930 3.960 3.090 ;
        RECT  3.780 1.900 3.940 2.660 ;
        RECT  3.500 1.030 3.870 1.190 ;
        RECT  3.660 0.590 3.820 0.870 ;
        RECT  3.560 1.360 3.680 1.520 ;
        RECT  3.400 1.360 3.560 3.090 ;
        RECT  3.340 0.500 3.500 1.190 ;
        RECT  1.780 2.930 3.400 3.090 ;
        RECT  1.450 0.500 3.340 0.660 ;
        RECT  3.180 1.620 3.220 1.900 ;
        RECT  3.020 1.000 3.180 2.770 ;
        RECT  2.400 1.000 3.020 1.160 ;
        RECT  2.120 2.610 3.020 2.770 ;
        RECT  2.680 1.320 2.860 1.590 ;
        RECT  2.520 1.320 2.680 2.310 ;
        RECT  2.240 1.320 2.520 1.480 ;
        RECT  2.080 2.150 2.520 2.310 ;
        RECT  2.080 0.820 2.240 1.480 ;
        RECT  1.800 0.820 2.080 0.980 ;
        RECT  1.620 2.480 1.780 3.090 ;
        RECT  0.790 2.480 1.620 2.640 ;
        RECT  1.290 0.500 1.450 1.950 ;
        RECT  1.020 1.790 1.290 1.950 ;
        RECT  0.700 1.320 1.070 1.630 ;
        RECT  0.860 1.790 1.020 2.190 ;
        RECT  0.700 2.480 0.790 3.130 ;
        RECT  0.630 1.320 0.700 3.130 ;
        RECT  0.540 1.320 0.630 2.640 ;
        RECT  0.310 1.320 0.540 1.480 ;
        RECT  0.150 1.020 0.310 1.480 ;
    END
END TLATNTSCAX2TR

MACRO TLATNTSCAX20TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.160 2.000 1.560 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.230 1.010 19.510 3.160 ;
        RECT  18.550 1.010 19.230 2.360 ;
        RECT  18.280 1.010 18.550 3.160 ;
        RECT  18.270 0.510 18.280 3.160 ;
        RECT  18.080 0.510 18.270 2.740 ;
        RECT  11.870 0.510 18.080 1.230 ;
        RECT  17.590 1.860 18.080 2.740 ;
        RECT  17.310 1.860 17.590 3.160 ;
        RECT  16.630 1.860 17.310 2.740 ;
        RECT  16.350 1.860 16.630 3.160 ;
        RECT  15.670 1.860 16.350 2.740 ;
        RECT  15.390 1.860 15.670 3.160 ;
        RECT  14.710 1.860 15.390 2.740 ;
        RECT  14.430 1.860 14.710 3.160 ;
        RECT  13.750 1.860 14.430 2.740 ;
        RECT  13.470 1.860 13.750 3.160 ;
        RECT  12.790 1.860 13.470 2.740 ;
        RECT  12.510 1.860 12.790 3.160 ;
        RECT  11.830 1.860 12.510 2.740 ;
        RECT  11.550 1.860 11.830 3.160 ;
        END
        ANTENNADIFFAREA 30.796 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.020 2.350 2.340 2.760 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.480 2.360 ;
        END
        ANTENNAGATEAREA 0.2736 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.990 -0.280 19.600 0.280 ;
        RECT  11.470 -0.280 18.990 0.340 ;
        RECT  10.510 -0.280 11.470 0.280 ;
        RECT  10.230 -0.280 10.510 0.800 ;
        RECT  9.470 -0.280 10.230 0.340 ;
        RECT  9.190 -0.280 9.470 0.800 ;
        RECT  8.430 -0.280 9.190 0.340 ;
        RECT  8.130 -0.280 8.430 1.010 ;
        RECT  6.740 -0.280 8.130 0.280 ;
        RECT  4.720 -0.280 6.740 0.340 ;
        RECT  3.320 -0.280 4.720 0.280 ;
        RECT  2.620 -0.280 3.320 0.300 ;
        RECT  0.950 -0.280 2.620 0.280 ;
        RECT  0.650 -0.280 0.950 0.720 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.030 3.320 19.600 3.880 ;
        RECT  18.750 2.720 19.030 3.880 ;
        RECT  18.070 3.320 18.750 3.880 ;
        RECT  17.790 2.930 18.070 3.880 ;
        RECT  17.110 3.320 17.790 3.880 ;
        RECT  16.830 2.930 17.110 3.880 ;
        RECT  16.150 3.320 16.830 3.880 ;
        RECT  15.870 2.930 16.150 3.880 ;
        RECT  15.190 3.320 15.870 3.880 ;
        RECT  14.910 2.930 15.190 3.880 ;
        RECT  14.230 3.320 14.910 3.880 ;
        RECT  13.950 2.930 14.230 3.880 ;
        RECT  13.270 3.320 13.950 3.880 ;
        RECT  12.990 2.930 13.270 3.880 ;
        RECT  12.310 3.320 12.990 3.880 ;
        RECT  12.030 2.930 12.310 3.880 ;
        RECT  11.350 3.320 12.030 3.880 ;
        RECT  11.070 2.040 11.350 3.880 ;
        RECT  10.390 3.320 11.070 3.880 ;
        RECT  10.110 2.040 10.390 3.880 ;
        RECT  9.430 3.320 10.110 3.880 ;
        RECT  9.150 2.040 9.430 3.880 ;
        RECT  8.470 3.320 9.150 3.880 ;
        RECT  8.190 1.980 8.470 3.880 ;
        RECT  6.770 3.320 8.190 3.880 ;
        RECT  6.090 3.240 6.770 3.880 ;
        RECT  3.320 3.320 6.090 3.880 ;
        RECT  1.160 3.260 3.320 3.880 ;
        RECT  0.390 3.320 1.160 3.880 ;
        RECT  0.110 2.520 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.670 1.390 17.890 1.670 ;
        RECT  11.390 1.390 11.670 1.550 ;
        RECT  11.230 0.960 11.390 1.880 ;
        RECT  11.030 0.960 11.230 1.120 ;
        RECT  10.870 1.720 11.230 1.880 ;
        RECT  8.470 1.280 11.070 1.560 ;
        RECT  10.750 0.840 11.030 1.120 ;
        RECT  10.590 1.720 10.870 3.160 ;
        RECT  9.990 0.960 10.750 1.120 ;
        RECT  9.910 1.720 10.590 1.880 ;
        RECT  9.710 0.840 9.990 1.120 ;
        RECT  9.630 1.720 9.910 3.160 ;
        RECT  8.950 0.960 9.710 1.120 ;
        RECT  8.950 1.720 9.630 1.880 ;
        RECT  8.670 0.840 8.950 1.120 ;
        RECT  8.670 1.720 8.950 3.160 ;
        RECT  7.670 1.280 8.470 1.440 ;
        RECT  7.990 1.600 8.270 1.820 ;
        RECT  7.830 1.600 7.990 3.120 ;
        RECT  7.660 0.500 7.950 1.120 ;
        RECT  7.070 2.960 7.830 3.120 ;
        RECT  7.390 1.280 7.670 2.800 ;
        RECT  5.710 0.500 7.660 0.660 ;
        RECT  7.230 0.950 7.390 1.460 ;
        RECT  6.980 0.950 7.230 1.230 ;
        RECT  6.910 1.540 7.070 3.120 ;
        RECT  6.790 1.540 6.910 1.820 ;
        RECT  5.920 2.790 6.910 2.950 ;
        RECT  6.470 1.070 6.630 2.030 ;
        RECT  6.230 1.070 6.470 1.230 ;
        RECT  6.230 1.870 6.470 2.030 ;
        RECT  5.710 1.390 6.310 1.670 ;
        RECT  5.950 0.950 6.230 1.230 ;
        RECT  5.870 1.870 6.230 2.490 ;
        RECT  5.750 2.790 5.920 3.150 ;
        RECT  3.720 2.990 5.750 3.150 ;
        RECT  5.550 0.500 5.710 2.300 ;
        RECT  5.340 0.500 5.550 0.660 ;
        RECT  5.350 2.140 5.550 2.300 ;
        RECT  5.110 0.960 5.390 1.240 ;
        RECT  5.070 2.140 5.350 2.820 ;
        RECT  5.060 0.500 5.340 0.800 ;
        RECT  4.360 1.080 5.110 1.240 ;
        RECT  4.150 2.140 5.070 2.300 ;
        RECT  3.880 0.500 5.060 0.780 ;
        RECT  4.280 1.080 4.360 1.980 ;
        RECT  4.120 0.940 4.280 1.980 ;
        RECT  3.880 2.140 4.150 2.420 ;
        RECT  3.600 0.940 4.120 1.100 ;
        RECT  4.080 1.700 4.120 1.980 ;
        RECT  3.720 1.260 3.960 1.540 ;
        RECT  3.560 1.260 3.720 3.150 ;
        RECT  3.440 0.460 3.600 1.100 ;
        RECT  0.870 2.920 3.560 3.080 ;
        RECT  1.490 0.460 3.440 0.620 ;
        RECT  3.280 1.320 3.400 1.600 ;
        RECT  3.120 0.950 3.280 2.530 ;
        RECT  2.520 0.950 3.120 1.230 ;
        RECT  2.800 2.370 3.120 2.530 ;
        RECT  2.680 1.390 2.960 2.190 ;
        RECT  2.520 2.370 2.800 2.730 ;
        RECT  2.320 1.390 2.680 1.550 ;
        RECT  2.390 1.910 2.680 2.190 ;
        RECT  2.160 0.780 2.320 1.550 ;
        RECT  1.960 0.780 2.160 1.000 ;
        RECT  1.330 0.460 1.490 2.190 ;
        RECT  1.100 1.910 1.330 2.190 ;
        RECT  0.800 1.360 1.110 1.640 ;
        RECT  0.800 2.880 0.870 3.160 ;
        RECT  0.640 0.910 0.800 3.160 ;
        RECT  0.390 0.910 0.640 1.070 ;
        RECT  0.110 0.440 0.390 1.070 ;
    END
END TLATNTSCAX20TR

MACRO TLATNTSCAX16TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.640 1.920 1.960 ;
        RECT  1.680 1.250 1.860 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.680 0.490 15.840 3.160 ;
        RECT  14.880 0.490 15.680 2.590 ;
        RECT  14.720 0.490 14.880 3.160 ;
        RECT  14.480 0.490 14.720 2.590 ;
        RECT  9.240 0.490 14.480 1.290 ;
        RECT  13.920 1.790 14.480 2.590 ;
        RECT  13.760 1.790 13.920 3.160 ;
        RECT  12.960 1.790 13.760 2.590 ;
        RECT  12.800 1.790 12.960 3.160 ;
        RECT  12.000 1.790 12.800 2.590 ;
        RECT  11.840 1.790 12.000 3.160 ;
        RECT  11.040 1.790 11.840 2.590 ;
        RECT  10.880 1.790 11.040 3.160 ;
        RECT  10.080 1.790 10.880 2.590 ;
        RECT  9.920 1.790 10.080 3.160 ;
        RECT  9.120 1.790 9.920 2.590 ;
        RECT  8.960 1.790 9.120 3.160 ;
        END
        ANTENNADIFFAREA 25.684 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 2.320 2.110 2.760 ;
        RECT  1.520 2.540 1.950 2.760 ;
        RECT  1.280 2.440 1.520 2.760 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.880 -0.280 16.000 0.280 ;
        RECT  7.600 -0.280 7.880 0.340 ;
        RECT  6.820 -0.280 7.600 0.280 ;
        RECT  6.080 -0.280 6.820 0.340 ;
        RECT  5.270 -0.280 6.080 0.280 ;
        RECT  4.990 -0.280 5.270 0.340 ;
        RECT  3.090 -0.280 4.990 0.280 ;
        RECT  2.530 -0.280 3.090 0.340 ;
        RECT  1.110 -0.280 2.530 0.280 ;
        RECT  0.830 -0.280 1.110 0.340 ;
        RECT  0.000 -0.280 0.830 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.360 3.320 16.000 3.880 ;
        RECT  15.200 2.930 15.360 3.880 ;
        RECT  14.400 3.320 15.200 3.880 ;
        RECT  14.240 2.930 14.400 3.880 ;
        RECT  13.440 3.320 14.240 3.880 ;
        RECT  13.280 2.930 13.440 3.880 ;
        RECT  12.480 3.320 13.280 3.880 ;
        RECT  12.320 2.930 12.480 3.880 ;
        RECT  11.520 3.320 12.320 3.880 ;
        RECT  11.360 2.930 11.520 3.880 ;
        RECT  10.560 3.320 11.360 3.880 ;
        RECT  10.400 2.930 10.560 3.880 ;
        RECT  9.600 3.320 10.400 3.880 ;
        RECT  9.440 2.930 9.600 3.880 ;
        RECT  8.640 3.320 9.440 3.880 ;
        RECT  8.480 2.000 8.640 3.880 ;
        RECT  7.680 3.320 8.480 3.880 ;
        RECT  7.520 2.000 7.680 3.880 ;
        RECT  6.740 3.320 7.520 3.880 ;
        RECT  6.460 3.260 6.740 3.880 ;
        RECT  5.180 3.320 6.460 3.880 ;
        RECT  4.500 3.260 5.180 3.880 ;
        RECT  3.010 3.320 4.500 3.880 ;
        RECT  2.730 3.260 3.010 3.880 ;
        RECT  1.590 3.320 2.730 3.880 ;
        RECT  1.310 3.260 1.590 3.880 ;
        RECT  0.590 3.320 1.310 3.880 ;
        RECT  0.310 2.930 0.590 3.880 ;
        RECT  0.000 3.320 0.310 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.700 1.470 14.260 1.630 ;
        RECT  8.540 0.920 8.700 1.840 ;
        RECT  8.340 0.920 8.540 1.080 ;
        RECT  8.160 1.680 8.540 1.840 ;
        RECT  6.980 1.240 8.380 1.520 ;
        RECT  8.180 0.800 8.340 1.080 ;
        RECT  7.300 0.920 8.180 1.080 ;
        RECT  8.000 1.680 8.160 3.160 ;
        RECT  7.200 1.680 8.000 1.840 ;
        RECT  7.140 0.800 7.300 1.080 ;
        RECT  7.040 1.680 7.200 3.160 ;
        RECT  6.940 0.940 6.980 1.520 ;
        RECT  6.820 0.940 6.940 1.400 ;
        RECT  6.220 0.940 6.820 1.100 ;
        RECT  6.540 1.520 6.660 1.680 ;
        RECT  6.380 1.520 6.540 2.930 ;
        RECT  5.360 2.700 6.380 2.930 ;
        RECT  6.060 0.940 6.220 2.130 ;
        RECT  5.560 0.940 6.060 1.100 ;
        RECT  5.740 1.970 6.060 2.130 ;
        RECT  5.740 1.260 5.900 1.720 ;
        RECT  5.400 1.260 5.740 1.420 ;
        RECT  5.240 0.540 5.400 1.420 ;
        RECT  5.200 1.580 5.360 2.930 ;
        RECT  4.380 0.540 5.240 0.700 ;
        RECT  4.100 2.770 5.200 2.930 ;
        RECT  4.880 0.970 5.040 2.130 ;
        RECT  4.550 0.970 4.880 1.130 ;
        RECT  4.700 1.970 4.880 2.130 ;
        RECT  4.380 1.430 4.720 1.710 ;
        RECT  4.540 1.970 4.700 2.610 ;
        RECT  4.260 2.450 4.540 2.610 ;
        RECT  4.220 0.540 4.380 2.290 ;
        RECT  3.670 0.540 4.220 0.700 ;
        RECT  3.750 2.130 4.220 2.290 ;
        RECT  3.940 2.660 4.100 2.930 ;
        RECT  3.840 0.860 4.000 1.930 ;
        RECT  3.590 2.660 3.940 2.820 ;
        RECT  3.510 0.860 3.840 1.020 ;
        RECT  3.590 1.280 3.670 1.550 ;
        RECT  3.430 1.280 3.590 3.080 ;
        RECT  3.350 0.500 3.510 1.020 ;
        RECT  1.010 2.920 3.430 3.080 ;
        RECT  1.460 0.500 3.350 0.660 ;
        RECT  3.190 1.280 3.270 1.560 ;
        RECT  3.030 0.980 3.190 2.750 ;
        RECT  2.450 0.980 3.030 1.140 ;
        RECT  2.550 2.590 3.030 2.750 ;
        RECT  2.710 1.300 2.870 2.130 ;
        RECT  2.230 1.300 2.710 1.460 ;
        RECT  2.130 1.970 2.710 2.130 ;
        RECT  2.390 2.470 2.550 2.750 ;
        RECT  2.070 0.820 2.230 1.460 ;
        RECT  1.870 0.820 2.070 0.980 ;
        RECT  1.300 0.500 1.460 1.960 ;
        RECT  1.070 1.800 1.300 1.960 ;
        RECT  0.750 1.360 1.140 1.640 ;
        RECT  0.910 1.800 1.070 2.190 ;
        RECT  0.850 2.350 1.010 3.150 ;
        RECT  0.750 2.350 0.850 2.510 ;
        RECT  0.590 1.150 0.750 2.510 ;
        RECT  0.530 1.150 0.590 1.310 ;
        RECT  0.370 0.570 0.530 1.310 ;
    END
END TLATNTSCAX16TR

MACRO TLATNTSCAX12TR
    CLASS CORE ;
    FOREIGN TLATNTSCAX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 2.040 1.920 2.360 ;
        RECT  1.610 1.280 1.890 2.360 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.180 0.630 13.460 3.160 ;
        RECT  12.680 0.630 13.180 2.770 ;
        RECT  8.580 0.630 12.680 1.350 ;
        RECT  12.500 2.050 12.680 2.770 ;
        RECT  12.220 2.050 12.500 3.160 ;
        RECT  11.540 2.050 12.220 2.770 ;
        RECT  11.260 2.050 11.540 3.160 ;
        RECT  10.580 2.050 11.260 2.770 ;
        RECT  10.300 2.050 10.580 3.160 ;
        RECT  9.620 2.050 10.300 2.770 ;
        RECT  9.340 2.050 9.620 3.160 ;
        RECT  8.660 2.050 9.340 2.770 ;
        RECT  8.380 2.050 8.660 3.160 ;
        END
        ANTENNADIFFAREA 18.958 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.360 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.940 -0.280 13.600 0.280 ;
        RECT  6.480 -0.280 12.940 0.340 ;
        RECT  6.200 -0.280 6.480 0.360 ;
        RECT  5.560 -0.280 6.200 0.340 ;
        RECT  4.800 -0.280 5.560 0.360 ;
        RECT  2.680 -0.280 4.800 0.280 ;
        RECT  2.400 -0.280 2.680 0.360 ;
        RECT  0.890 -0.280 2.400 0.280 ;
        RECT  0.610 -0.280 0.890 0.760 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.980 3.320 13.600 3.880 ;
        RECT  12.700 2.930 12.980 3.880 ;
        RECT  12.020 3.320 12.700 3.880 ;
        RECT  11.740 2.930 12.020 3.880 ;
        RECT  11.060 3.320 11.740 3.880 ;
        RECT  10.780 2.930 11.060 3.880 ;
        RECT  10.100 3.320 10.780 3.880 ;
        RECT  9.820 2.930 10.100 3.880 ;
        RECT  9.140 3.320 9.820 3.880 ;
        RECT  8.860 2.930 9.140 3.880 ;
        RECT  8.180 3.320 8.860 3.880 ;
        RECT  7.900 1.830 8.180 3.880 ;
        RECT  7.220 3.320 7.900 3.880 ;
        RECT  6.940 2.310 7.220 3.880 ;
        RECT  5.560 3.320 6.940 3.880 ;
        RECT  5.280 3.180 5.560 3.880 ;
        RECT  3.240 3.260 5.280 3.880 ;
        RECT  2.960 3.200 3.240 3.880 ;
        RECT  1.370 3.320 2.960 3.880 ;
        RECT  1.070 2.950 1.370 3.880 ;
        RECT  0.370 3.320 1.070 3.880 ;
        RECT  0.090 2.990 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.900 1.510 12.260 1.670 ;
        RECT  7.740 0.900 7.900 1.670 ;
        RECT  7.620 0.900 7.740 3.160 ;
        RECT  6.980 0.900 7.620 1.060 ;
        RECT  7.580 1.510 7.620 3.160 ;
        RECT  7.420 1.780 7.580 3.160 ;
        RECT  6.900 1.250 7.420 1.530 ;
        RECT  6.740 1.990 7.420 2.150 ;
        RECT  6.700 0.780 6.980 1.060 ;
        RECT  6.740 1.250 6.900 1.830 ;
        RECT  6.400 1.670 6.740 1.830 ;
        RECT  6.580 1.990 6.740 3.160 ;
        RECT  6.460 2.370 6.580 3.160 ;
        RECT  6.440 1.230 6.560 1.510 ;
        RECT  6.280 0.520 6.440 1.510 ;
        RECT  6.120 1.670 6.400 2.060 ;
        RECT  4.440 0.520 6.280 0.680 ;
        RECT  5.960 0.900 6.120 1.830 ;
        RECT  5.800 0.900 5.960 1.180 ;
        RECT  5.580 1.450 5.800 2.980 ;
        RECT  4.320 2.820 5.580 2.980 ;
        RECT  5.260 1.000 5.420 1.950 ;
        RECT  5.080 1.000 5.260 1.160 ;
        RECT  5.080 1.790 5.260 1.950 ;
        RECT  4.440 1.340 5.100 1.620 ;
        RECT  4.800 0.910 5.080 1.160 ;
        RECT  4.880 1.790 5.080 2.070 ;
        RECT  4.600 1.790 4.880 2.490 ;
        RECT  4.280 0.520 4.440 2.280 ;
        RECT  4.040 2.820 4.320 3.100 ;
        RECT  3.640 0.520 4.280 0.800 ;
        RECT  4.080 2.120 4.280 2.280 ;
        RECT  3.960 0.960 4.120 1.960 ;
        RECT  3.800 2.120 4.080 2.400 ;
        RECT  3.600 2.820 4.040 2.980 ;
        RECT  3.480 0.960 3.960 1.120 ;
        RECT  3.840 1.680 3.960 1.960 ;
        RECT  3.600 1.280 3.720 1.560 ;
        RECT  3.440 1.280 3.600 2.980 ;
        RECT  3.320 0.520 3.480 1.120 ;
        RECT  2.800 2.820 3.440 2.980 ;
        RECT  1.450 0.520 3.320 0.680 ;
        RECT  3.160 1.600 3.280 1.880 ;
        RECT  3.000 1.000 3.160 2.660 ;
        RECT  2.400 1.000 3.000 1.160 ;
        RECT  2.480 2.500 3.000 2.660 ;
        RECT  2.680 1.320 2.840 1.600 ;
        RECT  2.640 2.820 2.800 3.120 ;
        RECT  2.520 1.320 2.680 2.340 ;
        RECT  1.820 2.960 2.640 3.120 ;
        RECT  2.210 1.320 2.520 1.480 ;
        RECT  2.160 2.120 2.520 2.340 ;
        RECT  2.200 2.500 2.480 2.800 ;
        RECT  2.050 0.840 2.210 1.480 ;
        RECT  1.840 0.840 2.050 1.120 ;
        RECT  1.660 2.630 1.820 3.120 ;
        RECT  0.850 2.630 1.660 2.790 ;
        RECT  1.170 0.520 1.450 1.960 ;
        RECT  1.060 1.800 1.170 1.960 ;
        RECT  0.840 1.800 1.060 2.190 ;
        RECT  0.680 1.230 1.010 1.510 ;
        RECT  0.680 2.630 0.850 3.070 ;
        RECT  0.570 1.230 0.680 3.070 ;
        RECT  0.520 1.230 0.570 2.790 ;
        RECT  0.370 1.230 0.520 1.390 ;
        RECT  0.210 0.900 0.370 1.390 ;
        RECT  0.090 0.900 0.210 1.180 ;
    END
END TLATNTSCAX12TR

MACRO TLATNSRXLTR
    CLASS CORE ;
    FOREIGN TLATNSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.530 2.370 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 0.840 6.720 2.360 ;
        RECT  6.150 2.120 6.430 2.360 ;
        RECT  5.870 2.120 6.150 2.400 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.830 2.560 6.110 2.860 ;
        RECT  5.830 1.640 5.960 1.960 ;
        RECT  5.710 0.950 5.830 1.960 ;
        RECT  5.710 2.560 5.830 2.720 ;
        RECT  5.550 0.950 5.710 2.720 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.440 4.250 1.720 ;
        RECT  3.640 1.240 3.960 1.720 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.720 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.470 -0.280 6.800 0.280 ;
        RECT  6.190 -0.280 6.470 0.400 ;
        RECT  5.180 -0.280 6.190 0.280 ;
        RECT  4.900 -0.280 5.180 0.400 ;
        RECT  4.050 -0.280 4.900 0.280 ;
        RECT  3.770 -0.280 4.050 0.380 ;
        RECT  1.850 -0.280 3.770 0.280 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  0.370 -0.280 1.570 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.680 3.320 6.800 3.880 ;
        RECT  6.400 2.520 6.680 3.880 ;
        RECT  5.590 3.320 6.400 3.880 ;
        RECT  5.310 2.880 5.590 3.880 ;
        RECT  2.290 3.320 5.310 3.880 ;
        RECT  2.010 3.200 2.290 3.880 ;
        RECT  0.370 3.320 2.010 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 1.170 6.270 1.450 ;
        RECT  5.990 0.630 6.150 1.450 ;
        RECT  5.830 0.630 5.990 0.790 ;
        RECT  5.550 0.490 5.830 0.790 ;
        RECT  5.390 0.630 5.550 0.790 ;
        RECT  5.230 0.630 5.390 2.510 ;
        RECT  5.150 2.350 5.230 2.510 ;
        RECT  4.990 2.350 5.150 3.030 ;
        RECT  4.850 0.660 5.070 2.190 ;
        RECT  3.930 2.810 4.990 3.030 ;
        RECT  4.610 0.660 4.850 0.820 ;
        RECT  4.550 2.350 4.830 2.650 ;
        RECT  4.610 1.510 4.690 1.790 ;
        RECT  4.330 0.540 4.610 0.820 ;
        RECT  4.410 1.000 4.610 2.190 ;
        RECT  3.130 2.480 4.550 2.650 ;
        RECT  4.330 1.000 4.410 1.280 ;
        RECT  4.330 1.880 4.410 2.190 ;
        RECT  3.290 0.540 4.330 0.700 ;
        RECT  3.290 1.880 4.330 2.040 ;
        RECT  3.650 2.810 3.930 3.090 ;
        RECT  3.130 0.540 3.290 1.520 ;
        RECT  3.010 1.700 3.290 2.040 ;
        RECT  2.930 0.540 3.130 0.760 ;
        RECT  2.730 1.360 3.130 1.520 ;
        RECT  2.690 2.480 3.130 2.720 ;
        RECT  2.690 0.920 2.970 1.200 ;
        RECT  2.530 2.880 2.810 3.160 ;
        RECT  2.570 1.360 2.730 2.320 ;
        RECT  1.270 0.920 2.690 1.080 ;
        RECT  1.130 2.560 2.690 2.720 ;
        RECT  1.470 2.160 2.570 2.320 ;
        RECT  1.010 2.880 2.530 3.040 ;
        RECT  0.810 0.600 1.500 0.760 ;
        RECT  1.290 1.700 1.470 2.320 ;
        RECT  1.130 0.920 1.270 1.200 ;
        RECT  0.970 0.920 1.130 2.720 ;
        RECT  0.730 2.880 1.010 3.160 ;
        RECT  0.850 2.370 0.970 2.720 ;
        RECT  0.690 0.600 0.810 1.310 ;
        RECT  0.690 1.910 0.810 2.190 ;
        RECT  0.690 2.880 0.730 3.040 ;
        RECT  0.530 0.600 0.690 3.040 ;
    END
END TLATNSRXLTR

MACRO TLATNSRX4TR
    CLASS CORE ;
    FOREIGN TLATNSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.610 0.530 1.890 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.320 1.240 6.380 1.400 ;
        RECT  6.030 1.240 6.320 1.610 ;
        END
        ANTENNAGATEAREA 0.432 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.310 0.440 10.630 2.190 ;
        RECT  10.080 1.440 10.310 2.190 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.390 0.440 9.670 2.190 ;
        RECT  9.280 1.310 9.390 2.190 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.420 7.200 1.700 ;
        RECT  6.600 1.420 6.760 1.960 ;
        RECT  6.480 1.640 6.600 1.960 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.390 1.500 4.380 1.720 ;
        RECT  3.230 1.500 3.390 1.840 ;
        RECT  2.360 1.680 3.230 1.840 ;
        RECT  2.040 1.240 2.360 1.840 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 -0.280 11.200 0.280 ;
        RECT  10.830 -0.280 11.110 1.310 ;
        RECT  10.150 -0.280 10.830 0.280 ;
        RECT  9.870 -0.280 10.150 1.270 ;
        RECT  9.190 -0.280 9.870 0.280 ;
        RECT  8.910 -0.280 9.190 0.780 ;
        RECT  8.330 -0.280 8.910 0.340 ;
        RECT  8.050 -0.280 8.330 0.360 ;
        RECT  6.970 -0.280 8.050 0.280 ;
        RECT  6.690 -0.280 6.970 0.400 ;
        RECT  4.430 -0.280 6.690 0.280 ;
        RECT  4.150 -0.280 4.430 0.640 ;
        RECT  2.080 -0.280 4.150 0.280 ;
        RECT  1.800 -0.280 2.080 0.400 ;
        RECT  0.850 -0.280 1.800 0.280 ;
        RECT  0.570 -0.280 0.850 0.710 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 3.320 11.200 3.880 ;
        RECT  10.830 2.910 11.110 3.880 ;
        RECT  10.150 3.320 10.830 3.880 ;
        RECT  9.870 2.910 10.150 3.880 ;
        RECT  9.150 3.320 9.870 3.880 ;
        RECT  8.870 3.200 9.150 3.880 ;
        RECT  8.330 3.320 8.870 3.880 ;
        RECT  6.800 3.260 8.330 3.880 ;
        RECT  4.900 3.320 6.800 3.880 ;
        RECT  4.620 2.900 4.900 3.880 ;
        RECT  2.610 3.320 4.620 3.880 ;
        RECT  2.330 3.020 2.610 3.880 ;
        RECT  0.890 3.320 2.330 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.790 1.580 11.070 2.510 ;
        RECT  8.970 2.350 10.790 2.510 ;
        RECT  8.850 1.150 8.970 2.510 ;
        RECT  8.810 1.030 8.850 2.510 ;
        RECT  8.570 1.030 8.810 1.310 ;
        RECT  8.730 1.960 8.810 2.510 ;
        RECT  8.570 1.960 8.730 3.100 ;
        RECT  8.410 1.520 8.650 1.800 ;
        RECT  6.640 2.940 8.570 3.100 ;
        RECT  8.370 1.520 8.410 2.780 ;
        RECT  8.250 1.640 8.370 2.780 ;
        RECT  5.700 2.620 8.250 2.780 ;
        RECT  7.930 0.520 8.090 2.340 ;
        RECT  7.590 0.520 7.930 0.800 ;
        RECT  7.650 2.180 7.930 2.460 ;
        RECT  7.490 0.980 7.770 2.020 ;
        RECT  6.060 2.300 7.650 2.460 ;
        RECT  6.700 0.980 7.490 1.260 ;
        RECT  7.470 1.860 7.490 2.020 ;
        RECT  7.190 1.860 7.470 2.140 ;
        RECT  6.540 0.920 6.700 1.260 ;
        RECT  6.480 2.940 6.640 3.160 ;
        RECT  5.390 0.920 6.540 1.080 ;
        RECT  6.360 3.000 6.480 3.160 ;
        RECT  5.220 2.940 6.200 3.160 ;
        RECT  5.900 1.940 6.060 2.460 ;
        RECT  5.870 1.940 5.900 2.100 ;
        RECT  5.590 1.240 5.870 2.100 ;
        RECT  5.580 2.500 5.700 2.780 ;
        RECT  4.750 0.480 5.630 0.760 ;
        RECT  3.710 1.880 5.590 2.100 ;
        RECT  5.420 2.260 5.580 2.780 ;
        RECT  4.100 2.260 5.420 2.420 ;
        RECT  5.230 0.920 5.390 1.520 ;
        RECT  5.110 1.180 5.230 1.520 ;
        RECT  5.060 2.580 5.220 3.160 ;
        RECT  3.070 1.180 5.110 1.340 ;
        RECT  4.420 2.580 5.060 2.740 ;
        RECT  4.590 0.480 4.750 1.020 ;
        RECT  1.410 0.800 4.590 1.020 ;
        RECT  4.260 2.580 4.420 2.860 ;
        RECT  1.240 2.700 4.260 2.860 ;
        RECT  3.940 2.260 4.100 2.540 ;
        RECT  1.450 2.320 3.940 2.540 ;
        RECT  3.550 1.880 3.710 2.160 ;
        RECT  1.770 2.000 3.550 2.160 ;
        RECT  2.790 1.180 3.070 1.520 ;
        RECT  1.610 1.240 1.770 2.160 ;
        RECT  1.450 1.240 1.610 1.520 ;
        RECT  1.290 1.910 1.450 2.540 ;
        RECT  1.290 0.440 1.410 1.080 ;
        RECT  1.130 0.440 1.290 2.540 ;
        RECT  0.970 2.700 1.240 3.040 ;
        RECT  0.810 0.920 0.970 3.040 ;
        RECT  0.690 0.920 0.810 2.740 ;
        RECT  0.370 0.920 0.690 1.080 ;
        RECT  0.370 2.520 0.690 2.740 ;
        RECT  0.090 0.440 0.370 1.080 ;
        RECT  0.090 2.520 0.370 3.160 ;
    END
END TLATNSRX4TR

MACRO TLATNSRX2TR
    CLASS CORE ;
    FOREIGN TLATNSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.320 0.410 1.620 ;
        RECT  0.080 1.320 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.670 1.240 2.720 1.560 ;
        RECT  2.430 1.240 2.670 2.120 ;
        END
        ANTENNAGATEAREA 0.2376 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.500 0.840 7.520 1.960 ;
        RECT  7.280 0.440 7.500 3.160 ;
        RECT  7.230 0.440 7.280 1.290 ;
        END
        ANTENNADIFFAREA 3.488 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.320 1.010 6.590 2.200 ;
        RECT  6.240 1.010 6.320 1.960 ;
        RECT  6.080 1.640 6.240 1.960 ;
        END
        ANTENNADIFFAREA 2.516 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.030 1.580 4.580 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.560 2.230 1.960 ;
        END
        ANTENNAGATEAREA 0.2232 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.980 -0.280 7.600 0.280 ;
        RECT  6.700 -0.280 6.980 0.300 ;
        RECT  5.600 -0.280 6.700 0.280 ;
        RECT  5.320 -0.280 5.600 0.300 ;
        RECT  4.400 -0.280 5.320 0.280 ;
        RECT  4.120 -0.280 4.400 0.300 ;
        RECT  2.130 -0.280 4.120 0.280 ;
        RECT  1.850 -0.280 2.130 0.300 ;
        RECT  0.370 -0.280 1.850 0.280 ;
        RECT  0.090 -0.280 0.370 1.040 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.030 3.320 7.600 3.880 ;
        RECT  6.740 2.920 7.030 3.880 ;
        RECT  2.530 3.320 6.740 3.880 ;
        RECT  2.250 3.260 2.530 3.880 ;
        RECT  0.410 3.320 2.250 3.880 ;
        RECT  0.130 3.260 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.990 1.470 7.120 1.760 ;
        RECT  6.830 0.600 6.990 2.760 ;
        RECT  6.060 0.600 6.830 0.760 ;
        RECT  6.140 2.600 6.830 2.760 ;
        RECT  5.980 2.380 6.140 3.160 ;
        RECT  5.900 0.480 6.060 0.760 ;
        RECT  4.260 3.000 5.980 3.160 ;
        RECT  5.820 1.440 5.880 1.790 ;
        RECT  5.660 1.440 5.820 2.840 ;
        RECT  4.580 2.680 5.660 2.840 ;
        RECT  5.340 0.660 5.500 1.960 ;
        RECT  5.000 0.660 5.340 0.820 ;
        RECT  5.220 1.800 5.340 1.960 ;
        RECT  5.060 1.800 5.220 2.120 ;
        RECT  5.020 1.020 5.180 1.640 ;
        RECT  4.900 2.360 5.070 2.520 ;
        RECT  3.870 1.020 5.020 1.180 ;
        RECT  4.900 1.480 5.020 1.640 ;
        RECT  4.720 0.540 5.000 0.820 ;
        RECT  4.740 1.480 4.900 2.520 ;
        RECT  3.550 0.660 4.720 0.820 ;
        RECT  4.420 2.390 4.580 2.840 ;
        RECT  3.330 2.390 4.420 2.550 ;
        RECT  4.040 2.760 4.260 3.160 ;
        RECT  3.720 1.020 3.870 1.900 ;
        RECT  3.710 1.020 3.720 2.040 ;
        RECT  3.360 1.740 3.710 2.040 ;
        RECT  2.850 3.000 3.580 3.160 ;
        RECT  3.390 0.660 3.550 1.580 ;
        RECT  3.250 0.660 3.390 0.820 ;
        RECT  3.050 1.420 3.390 1.580 ;
        RECT  3.310 2.390 3.330 2.760 ;
        RECT  3.150 2.220 3.310 2.760 ;
        RECT  3.070 0.980 3.230 1.260 ;
        RECT  1.370 2.600 3.150 2.760 ;
        RECT  3.060 0.980 3.070 1.140 ;
        RECT  2.890 0.920 3.060 1.140 ;
        RECT  2.990 1.420 3.050 1.890 ;
        RECT  2.890 1.420 2.990 2.440 ;
        RECT  2.210 0.920 2.890 1.080 ;
        RECT  2.830 1.720 2.890 2.440 ;
        RECT  2.690 2.940 2.850 3.160 ;
        RECT  1.520 2.280 2.830 2.440 ;
        RECT  1.690 2.940 2.690 3.100 ;
        RECT  2.020 0.920 2.210 1.200 ;
        RECT  1.180 1.040 2.020 1.200 ;
        RECT  0.850 0.520 1.740 0.680 ;
        RECT  1.530 2.940 1.690 3.160 ;
        RECT  0.850 3.000 1.530 3.160 ;
        RECT  1.350 1.680 1.520 2.440 ;
        RECT  1.180 2.600 1.370 2.840 ;
        RECT  1.020 1.040 1.180 2.840 ;
        RECT  0.690 0.520 0.850 3.160 ;
        RECT  0.580 0.830 0.690 1.080 ;
    END
END TLATNSRX2TR

MACRO TLATNSRX1TR
    CLASS CORE ;
    FOREIGN TLATNSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.570 1.960 ;
        END
        ANTENNAGATEAREA 0.1464 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.830 0.600 7.120 2.360 ;
        RECT  6.470 2.120 6.830 2.360 ;
        RECT  6.190 2.120 6.470 2.400 ;
        END
        ANTENNADIFFAREA 2.028 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.120 2.630 6.400 2.910 ;
        RECT  6.100 1.640 6.360 1.960 ;
        RECT  6.030 2.630 6.120 2.790 ;
        RECT  6.030 0.990 6.100 1.960 ;
        RECT  5.870 0.990 6.030 2.790 ;
        RECT  5.820 0.990 5.870 1.800 ;
        END
        ANTENNADIFFAREA 1.684 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.460 4.410 1.740 ;
        RECT  3.960 1.460 4.130 1.620 ;
        RECT  3.640 1.240 3.960 1.620 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.690 -0.280 7.200 0.280 ;
        RECT  6.410 -0.280 6.690 0.360 ;
        RECT  5.420 -0.280 6.410 0.280 ;
        RECT  5.120 -0.280 5.420 0.390 ;
        RECT  4.170 -0.280 5.120 0.280 ;
        RECT  3.890 -0.280 4.170 0.360 ;
        RECT  1.970 -0.280 3.890 0.280 ;
        RECT  1.690 -0.280 1.970 0.400 ;
        RECT  0.370 -0.280 1.690 0.280 ;
        RECT  0.090 -0.280 0.370 0.360 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.870 3.320 7.200 3.880 ;
        RECT  6.590 2.800 6.870 3.880 ;
        RECT  5.710 3.320 6.590 3.880 ;
        RECT  5.430 2.930 5.710 3.880 ;
        RECT  4.490 3.260 5.430 3.880 ;
        RECT  4.210 3.200 4.490 3.880 ;
        RECT  2.410 3.320 4.210 3.880 ;
        RECT  2.130 3.200 2.410 3.880 ;
        RECT  0.370 3.320 2.130 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.550 0.930 6.670 1.210 ;
        RECT  6.390 0.670 6.550 1.210 ;
        RECT  6.100 0.670 6.390 0.830 ;
        RECT  5.820 0.450 6.100 0.830 ;
        RECT  5.660 0.670 5.820 0.830 ;
        RECT  5.500 0.670 5.660 2.540 ;
        RECT  5.270 2.380 5.500 2.540 ;
        RECT  5.180 0.640 5.340 2.220 ;
        RECT  5.110 2.380 5.270 3.040 ;
        RECT  4.780 0.640 5.180 0.800 ;
        RECT  5.060 1.940 5.180 2.220 ;
        RECT  4.870 2.760 5.110 3.040 ;
        RECT  4.730 1.500 5.020 1.780 ;
        RECT  3.210 2.380 4.950 2.600 ;
        RECT  4.050 2.880 4.870 3.040 ;
        RECT  4.500 0.520 4.780 0.800 ;
        RECT  4.570 0.980 4.730 2.180 ;
        RECT  4.450 0.980 4.570 1.260 ;
        RECT  4.410 1.900 4.570 2.180 ;
        RECT  3.410 0.520 4.500 0.680 ;
        RECT  3.330 1.900 4.410 2.060 ;
        RECT  3.770 2.880 4.050 3.160 ;
        RECT  3.250 0.520 3.410 1.520 ;
        RECT  3.050 1.750 3.330 2.060 ;
        RECT  3.050 0.520 3.250 0.760 ;
        RECT  2.890 1.360 3.250 1.520 ;
        RECT  3.050 2.380 3.210 2.720 ;
        RECT  2.810 0.920 3.090 1.200 ;
        RECT  1.250 2.440 3.050 2.720 ;
        RECT  2.650 2.880 2.930 3.160 ;
        RECT  2.730 1.360 2.890 2.280 ;
        RECT  1.270 0.920 2.810 1.080 ;
        RECT  1.520 2.120 2.730 2.280 ;
        RECT  1.610 2.880 2.650 3.040 ;
        RECT  1.410 2.880 1.610 3.160 ;
        RECT  1.300 1.670 1.520 2.280 ;
        RECT  1.230 0.480 1.510 0.760 ;
        RECT  0.810 3.000 1.410 3.160 ;
        RECT  1.140 0.920 1.270 1.240 ;
        RECT  1.140 2.440 1.250 2.840 ;
        RECT  0.810 0.600 1.230 0.760 ;
        RECT  0.990 0.920 1.140 2.840 ;
        RECT  0.980 1.080 0.990 2.840 ;
        RECT  0.970 2.560 0.980 2.840 ;
        RECT  0.690 0.600 0.810 1.250 ;
        RECT  0.690 1.910 0.810 3.160 ;
        RECT  0.530 0.600 0.690 3.160 ;
    END
END TLATNSRX1TR

MACRO TLATNCAX8TR
    CLASS CORE ;
    FOREIGN TLATNCAX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.210 0.600 13.520 3.160 ;
        RECT  13.130 0.600 13.210 2.360 ;
        RECT  8.330 0.600 13.130 1.080 ;
        RECT  11.890 1.880 13.130 2.360 ;
        RECT  11.610 1.880 11.890 3.160 ;
        RECT  10.290 1.880 11.610 2.360 ;
        RECT  10.010 1.880 10.290 3.160 ;
        RECT  8.920 1.880 10.010 2.360 ;
        RECT  8.280 1.880 8.920 3.160 ;
        END
        ANTENNADIFFAREA 12.596 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.890 1.600 6.170 2.220 ;
        RECT  4.530 2.060 5.890 2.220 ;
        RECT  4.250 1.600 4.530 2.220 ;
        RECT  2.850 2.060 4.250 2.220 ;
        RECT  2.760 1.620 2.850 2.220 ;
        RECT  2.480 1.620 2.760 2.360 ;
        END
        ANTENNAGATEAREA 1.008 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.240 1.030 1.680 ;
        END
        ANTENNAGATEAREA 0.7992 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.370 -0.280 13.600 0.280 ;
        RECT  13.090 -0.280 13.370 0.400 ;
        RECT  12.330 -0.280 13.090 0.340 ;
        RECT  12.050 -0.280 12.330 0.400 ;
        RECT  11.290 -0.280 12.050 0.340 ;
        RECT  11.010 -0.280 11.290 0.400 ;
        RECT  10.250 -0.280 11.010 0.340 ;
        RECT  9.970 -0.280 10.250 0.400 ;
        RECT  9.130 -0.280 9.970 0.340 ;
        RECT  8.850 -0.280 9.130 0.400 ;
        RECT  8.090 -0.280 8.850 0.280 ;
        RECT  8.080 -0.280 8.090 0.640 ;
        RECT  7.800 -0.280 8.080 1.040 ;
        RECT  7.110 -0.280 7.800 0.640 ;
        RECT  6.050 -0.280 7.110 0.340 ;
        RECT  5.770 -0.280 6.050 0.400 ;
        RECT  4.370 -0.280 5.770 0.280 ;
        RECT  4.090 -0.280 4.370 0.400 ;
        RECT  2.650 -0.280 4.090 0.280 ;
        RECT  1.570 -0.280 2.650 0.340 ;
        RECT  0.850 -0.280 1.570 0.280 ;
        RECT  0.570 -0.280 0.850 1.080 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.690 3.320 13.600 3.880 ;
        RECT  12.410 2.930 12.690 3.880 ;
        RECT  11.090 3.320 12.410 3.880 ;
        RECT  10.810 2.520 11.090 3.880 ;
        RECT  9.490 3.320 10.810 3.880 ;
        RECT  9.210 2.520 9.490 3.880 ;
        RECT  7.850 3.320 9.210 3.880 ;
        RECT  7.100 3.180 7.850 3.880 ;
        RECT  6.010 3.260 7.100 3.880 ;
        RECT  5.730 3.200 6.010 3.880 ;
        RECT  4.330 3.320 5.730 3.880 ;
        RECT  4.050 3.200 4.330 3.880 ;
        RECT  2.650 3.320 4.050 3.880 ;
        RECT  2.370 3.200 2.650 3.880 ;
        RECT  1.850 3.260 2.370 3.880 ;
        RECT  1.570 3.200 1.850 3.880 ;
        RECT  0.850 3.320 1.570 3.880 ;
        RECT  0.570 2.160 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.590 1.240 12.970 1.400 ;
        RECT  8.030 1.560 12.490 1.720 ;
        RECT  7.870 1.560 8.030 2.980 ;
        RECT  6.610 2.820 7.870 2.980 ;
        RECT  7.430 1.240 7.590 2.660 ;
        RECT  6.490 2.500 7.430 2.660 ;
        RECT  7.110 1.020 7.270 2.300 ;
        RECT  6.650 1.850 7.110 2.010 ;
        RECT  6.730 0.650 6.890 1.690 ;
        RECT  5.730 0.650 6.730 0.930 ;
        RECT  6.490 1.530 6.730 1.690 ;
        RECT  6.330 2.820 6.610 3.100 ;
        RECT  5.730 1.090 6.570 1.370 ;
        RECT  6.330 1.530 6.490 2.660 ;
        RECT  6.090 2.380 6.330 2.660 ;
        RECT  1.350 2.820 6.330 2.980 ;
        RECT  5.170 2.380 6.090 2.540 ;
        RECT  5.570 0.640 5.730 0.930 ;
        RECT  5.570 1.090 5.730 1.900 ;
        RECT  5.210 0.640 5.570 0.800 ;
        RECT  4.970 1.740 5.570 1.900 ;
        RECT  5.130 0.960 5.410 1.560 ;
        RECT  4.930 0.520 5.210 0.800 ;
        RECT  4.890 2.380 5.170 2.660 ;
        RECT  3.730 0.960 5.130 1.120 ;
        RECT  4.850 1.620 4.970 1.900 ;
        RECT  3.530 0.640 4.930 0.800 ;
        RECT  3.490 2.380 4.890 2.540 ;
        RECT  4.690 1.280 4.850 1.900 ;
        RECT  4.050 1.280 4.690 1.440 ;
        RECT  3.890 1.280 4.050 1.900 ;
        RECT  3.290 1.740 3.890 1.900 ;
        RECT  3.450 0.960 3.730 1.560 ;
        RECT  3.250 0.520 3.530 0.800 ;
        RECT  3.210 2.380 3.490 2.660 ;
        RECT  2.630 0.960 3.450 1.120 ;
        RECT  3.010 1.300 3.290 1.900 ;
        RECT  2.310 1.300 3.010 1.460 ;
        RECT  2.470 0.500 2.630 1.120 ;
        RECT  1.350 0.500 2.470 0.660 ;
        RECT  2.250 1.040 2.310 2.320 ;
        RECT  2.150 0.920 2.250 2.320 ;
        RECT  1.970 0.920 2.150 1.200 ;
        RECT  1.970 2.040 2.150 2.320 ;
        RECT  1.770 1.360 1.990 1.880 ;
        RECT  1.350 1.360 1.770 1.520 ;
        RECT  1.330 0.500 1.350 2.980 ;
        RECT  1.190 0.500 1.330 3.160 ;
        RECT  1.050 0.500 1.190 1.080 ;
        RECT  1.050 1.840 1.190 3.160 ;
        RECT  0.370 1.840 1.050 2.000 ;
        RECT  0.250 0.440 0.370 1.080 ;
        RECT  0.250 1.840 0.370 3.160 ;
        RECT  0.090 0.440 0.250 3.160 ;
    END
END TLATNCAX8TR

MACRO TLATNCAX6TR
    CLASS CORE ;
    FOREIGN TLATNCAX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 0.780 7.920 3.160 ;
        RECT  7.360 0.780 7.640 1.120 ;
        RECT  7.630 1.840 7.640 3.160 ;
        RECT  7.080 1.840 7.630 2.560 ;
        RECT  7.080 0.440 7.360 1.120 ;
        RECT  6.400 0.780 7.080 1.120 ;
        RECT  6.310 2.040 7.080 2.560 ;
        RECT  6.120 0.440 6.400 1.120 ;
        RECT  6.030 2.040 6.310 3.160 ;
        END
        ANTENNADIFFAREA 6.368 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.640 3.960 2.260 ;
        RECT  2.210 2.100 3.600 2.260 ;
        RECT  2.050 1.660 2.210 2.260 ;
        END
        ANTENNAGATEAREA 0.504 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.560 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.880 -0.280 8.000 0.280 ;
        RECT  7.600 -0.280 7.880 0.400 ;
        RECT  6.880 -0.280 7.600 0.280 ;
        RECT  6.600 -0.280 6.880 0.620 ;
        RECT  5.920 -0.280 6.600 0.280 ;
        RECT  5.640 -0.280 5.920 0.680 ;
        RECT  3.760 -0.280 5.640 0.340 ;
        RECT  3.480 -0.280 3.760 0.370 ;
        RECT  2.080 -0.280 3.480 0.280 ;
        RECT  1.090 -0.280 2.080 0.400 ;
        RECT  0.370 -0.280 1.090 0.340 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.320 8.000 3.880 ;
        RECT  6.830 2.900 7.110 3.880 ;
        RECT  5.370 3.320 6.830 3.880 ;
        RECT  5.000 3.200 5.370 3.880 ;
        RECT  3.710 3.320 5.000 3.880 ;
        RECT  3.430 3.200 3.710 3.880 ;
        RECT  2.030 3.320 3.430 3.880 ;
        RECT  1.090 3.200 2.030 3.880 ;
        RECT  0.370 3.320 1.090 3.880 ;
        RECT  0.090 2.250 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.480 1.280 7.480 1.440 ;
        RECT  6.630 1.600 6.910 1.880 ;
        RECT  5.640 1.720 6.630 1.880 ;
        RECT  5.520 1.600 5.640 1.880 ;
        RECT  5.360 1.600 5.520 3.040 ;
        RECT  5.260 0.500 5.480 1.440 ;
        RECT  4.360 2.880 5.360 3.040 ;
        RECT  4.600 0.500 5.260 0.660 ;
        RECT  5.000 0.820 5.070 1.100 ;
        RECT  4.820 0.820 5.000 2.370 ;
        RECT  4.720 1.690 4.820 2.370 ;
        RECT  4.480 1.690 4.720 1.970 ;
        RECT  4.440 0.500 4.600 1.530 ;
        RECT  3.320 0.550 4.440 0.770 ;
        RECT  4.280 1.370 4.440 1.530 ;
        RECT  4.080 2.880 4.360 3.160 ;
        RECT  4.000 0.930 4.280 1.210 ;
        RECT  4.120 1.370 4.280 2.600 ;
        RECT  3.840 2.440 4.120 2.720 ;
        RECT  1.080 2.880 4.080 3.040 ;
        RECT  3.440 1.050 4.000 1.210 ;
        RECT  2.870 2.440 3.840 2.600 ;
        RECT  3.280 1.050 3.440 1.940 ;
        RECT  2.640 0.490 3.320 0.770 ;
        RECT  2.650 1.780 3.280 1.940 ;
        RECT  3.000 1.320 3.120 1.600 ;
        RECT  2.840 0.930 3.000 1.600 ;
        RECT  2.590 2.440 2.870 2.720 ;
        RECT  2.210 0.930 2.840 1.090 ;
        RECT  2.490 1.340 2.650 1.940 ;
        RECT  1.890 1.340 2.490 1.500 ;
        RECT  2.050 0.620 2.210 1.090 ;
        RECT  0.850 0.620 2.050 0.780 ;
        RECT  1.730 0.940 1.890 2.270 ;
        RECT  1.430 0.940 1.730 1.220 ;
        RECT  1.390 1.990 1.730 2.270 ;
        RECT  1.080 1.380 1.570 1.660 ;
        RECT  0.920 1.150 1.080 3.040 ;
        RECT  0.850 1.150 0.920 1.310 ;
        RECT  0.850 2.250 0.920 3.040 ;
        RECT  0.570 0.620 0.850 1.310 ;
        RECT  0.570 2.250 0.850 3.160 ;
    END
END TLATNCAX6TR

MACRO TLATNCAX4TR
    CLASS CORE ;
    FOREIGN TLATNCAX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.590 1.020 6.710 1.270 ;
        RECT  6.430 1.020 6.590 2.040 ;
        RECT  6.090 1.800 6.430 2.040 ;
        RECT  5.910 1.800 6.090 2.720 ;
        RECT  5.680 0.990 5.910 2.720 ;
        RECT  5.480 0.990 5.680 1.270 ;
        END
        ANTENNADIFFAREA 4.382 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.680 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.720 1.670 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 -0.280 7.200 0.280 ;
        RECT  6.830 -0.280 7.110 0.710 ;
        RECT  6.160 -0.280 6.830 0.340 ;
        RECT  5.880 -0.280 6.160 0.400 ;
        RECT  5.240 -0.280 5.880 0.340 ;
        RECT  4.430 -0.280 5.240 0.400 ;
        RECT  3.460 -0.280 4.430 0.340 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  1.780 -0.280 3.180 0.280 ;
        RECT  0.800 -0.280 1.780 0.400 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.010 3.320 7.200 3.880 ;
        RECT  6.730 2.520 7.010 3.880 ;
        RECT  5.250 3.320 6.730 3.880 ;
        RECT  4.430 3.200 5.250 3.880 ;
        RECT  3.460 3.260 4.430 3.880 ;
        RECT  3.180 3.200 3.460 3.880 ;
        RECT  1.780 3.320 3.180 3.880 ;
        RECT  0.760 2.800 1.780 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.910 1.590 7.030 1.870 ;
        RECT  6.750 1.590 6.910 2.360 ;
        RECT  6.480 2.200 6.750 2.360 ;
        RECT  6.320 2.200 6.480 3.040 ;
        RECT  5.430 2.880 6.320 3.040 ;
        RECT  6.070 0.660 6.270 1.630 ;
        RECT  4.360 0.660 6.070 0.830 ;
        RECT  5.270 1.430 5.430 3.040 ;
        RECT  4.120 2.880 5.270 3.040 ;
        RECT  4.950 1.170 5.110 2.090 ;
        RECT  4.800 1.170 4.950 1.330 ;
        RECT  4.800 1.930 4.950 2.090 ;
        RECT  4.520 1.030 4.800 1.330 ;
        RECT  4.560 1.930 4.800 2.210 ;
        RECT  4.360 1.490 4.790 1.770 ;
        RECT  4.280 1.930 4.560 2.620 ;
        RECT  4.200 0.660 4.360 1.770 ;
        RECT  3.520 0.660 4.200 0.930 ;
        RECT  3.630 1.610 4.200 1.770 ;
        RECT  3.960 2.000 4.120 3.040 ;
        RECT  3.760 1.090 4.040 1.370 ;
        RECT  3.790 2.000 3.960 2.280 ;
        RECT  2.180 2.880 3.960 3.040 ;
        RECT  3.630 2.440 3.800 2.720 ;
        RECT  3.140 1.210 3.760 1.370 ;
        RECT  3.470 1.610 3.630 2.720 ;
        RECT  2.620 0.770 3.520 0.930 ;
        RECT  2.620 2.560 3.470 2.720 ;
        RECT  2.980 1.210 3.140 1.990 ;
        RECT  2.820 1.830 2.980 1.990 ;
        RECT  2.240 1.390 2.820 1.670 ;
        RECT  2.240 1.830 2.820 2.110 ;
        RECT  2.400 0.770 2.620 1.050 ;
        RECT  2.400 2.440 2.620 2.720 ;
        RECT  2.080 0.680 2.240 1.670 ;
        RECT  2.140 1.830 2.240 2.240 ;
        RECT  2.020 2.400 2.180 3.040 ;
        RECT  2.080 1.950 2.140 2.240 ;
        RECT  1.040 0.680 2.080 0.840 ;
        RECT  1.480 2.080 2.080 2.240 ;
        RECT  1.040 2.400 2.020 2.560 ;
        RECT  1.320 1.010 1.480 2.240 ;
        RECT  1.200 1.010 1.320 1.310 ;
        RECT  1.200 1.960 1.320 2.240 ;
        RECT  1.040 1.520 1.160 1.800 ;
        RECT  0.880 0.680 1.040 2.560 ;
        RECT  0.560 0.920 0.880 1.080 ;
        RECT  0.560 1.940 0.880 2.560 ;
        RECT  0.280 0.440 0.560 1.080 ;
        RECT  0.280 1.940 0.560 3.160 ;
    END
END TLATNCAX4TR

MACRO TLATNCAX3TR
    CLASS CORE ;
    FOREIGN TLATNCAX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.600 1.910 4.880 2.720 ;
        RECT  4.440 1.030 4.600 2.720 ;
        RECT  4.320 1.030 4.440 1.310 ;
        END
        ANTENNADIFFAREA 3.296 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.620 ;
        END
        ANTENNAGATEAREA 0.2496 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.480 -0.280 6.000 0.280 ;
        RECT  5.200 -0.280 5.480 1.310 ;
        RECT  4.040 -0.280 5.200 0.340 ;
        RECT  3.330 -0.280 4.040 0.400 ;
        RECT  1.760 -0.280 3.330 0.280 ;
        RECT  1.480 -0.280 1.760 0.670 ;
        RECT  0.380 -0.280 1.480 0.340 ;
        RECT  0.100 -0.280 0.380 1.080 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.800 3.320 6.000 3.880 ;
        RECT  5.520 2.020 5.800 3.880 ;
        RECT  4.040 3.260 5.520 3.880 ;
        RECT  3.140 3.200 4.040 3.880 ;
        RECT  1.550 3.320 3.140 3.880 ;
        RECT  1.200 2.770 1.550 3.880 ;
        RECT  0.380 3.320 1.200 3.880 ;
        RECT  0.100 2.770 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.360 1.580 5.480 1.860 ;
        RECT  5.200 1.580 5.360 3.040 ;
        RECT  4.280 2.880 5.200 3.040 ;
        RECT  4.760 0.600 5.040 1.750 ;
        RECT  3.120 0.600 4.760 0.760 ;
        RECT  4.060 1.580 4.280 3.040 ;
        RECT  2.710 2.870 4.060 3.040 ;
        RECT  3.740 1.150 3.900 2.070 ;
        RECT  3.600 1.150 3.740 1.310 ;
        RECT  3.640 1.910 3.740 2.070 ;
        RECT  3.360 1.910 3.640 2.540 ;
        RECT  3.320 1.030 3.600 1.310 ;
        RECT  3.120 1.470 3.580 1.750 ;
        RECT  2.900 2.260 3.360 2.540 ;
        RECT  2.960 0.600 3.120 1.750 ;
        RECT  2.560 0.600 2.960 0.760 ;
        RECT  2.700 1.470 2.960 1.750 ;
        RECT  2.640 0.920 2.800 1.200 ;
        RECT  2.390 2.870 2.710 3.140 ;
        RECT  2.520 1.470 2.700 2.390 ;
        RECT  1.320 0.920 2.640 1.080 ;
        RECT  2.280 0.480 2.560 0.760 ;
        RECT  2.160 2.110 2.520 2.390 ;
        RECT  2.000 2.870 2.390 3.050 ;
        RECT  2.240 1.270 2.360 1.550 ;
        RECT  2.080 1.270 2.240 1.940 ;
        RECT  2.000 1.780 2.080 1.940 ;
        RECT  1.840 1.780 2.000 3.050 ;
        RECT  0.860 2.450 1.840 2.610 ;
        RECT  1.160 0.570 1.320 2.220 ;
        RECT  0.920 0.570 1.160 0.850 ;
        RECT  0.960 1.940 1.160 2.220 ;
        RECT  0.800 1.030 1.000 1.710 ;
        RECT  0.800 2.450 0.860 2.830 ;
        RECT  0.640 1.030 0.800 2.830 ;
        RECT  0.580 2.550 0.640 2.830 ;
    END
END TLATNCAX3TR

MACRO TLATNCAX2TR
    CLASS CORE ;
    FOREIGN TLATNCAX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.910 4.720 3.160 ;
        RECT  4.340 1.910 4.400 2.070 ;
        RECT  4.180 1.030 4.340 2.070 ;
        RECT  4.030 1.030 4.180 1.310 ;
        END
        ANTENNADIFFAREA 2.764 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.200 1.920 1.580 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.350 1.960 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.280 4.800 0.280 ;
        RECT  4.430 -0.280 4.710 0.400 ;
        RECT  3.790 -0.280 4.430 0.340 ;
        RECT  3.050 -0.280 3.790 0.400 ;
        RECT  1.620 -0.280 3.050 0.280 ;
        RECT  1.340 -0.280 1.620 0.710 ;
        RECT  0.370 -0.280 1.340 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 3.320 4.800 3.880 ;
        RECT  3.560 3.200 3.840 3.880 ;
        RECT  3.180 3.320 3.560 3.880 ;
        RECT  2.900 3.200 3.180 3.880 ;
        RECT  1.450 3.320 2.900 3.880 ;
        RECT  1.170 2.800 1.450 3.880 ;
        RECT  0.450 3.320 1.170 3.880 ;
        RECT  0.170 2.930 0.450 3.880 ;
        RECT  0.000 3.320 0.170 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.500 0.560 4.720 1.640 ;
        RECT  2.940 0.560 4.500 0.720 ;
        RECT  3.860 1.580 4.020 3.010 ;
        RECT  2.530 2.850 3.860 3.010 ;
        RECT  3.540 1.150 3.700 2.070 ;
        RECT  3.350 1.150 3.540 1.310 ;
        RECT  3.400 1.910 3.540 2.070 ;
        RECT  3.100 1.910 3.400 2.590 ;
        RECT  2.940 1.470 3.380 1.750 ;
        RECT  3.130 1.030 3.350 1.310 ;
        RECT  2.780 0.560 2.940 2.360 ;
        RECT  2.420 0.560 2.780 0.720 ;
        RECT  2.010 2.080 2.780 2.360 ;
        RECT  2.460 0.880 2.620 1.920 ;
        RECT  1.850 2.850 2.530 3.130 ;
        RECT  1.380 0.880 2.460 1.040 ;
        RECT  2.400 1.640 2.460 1.920 ;
        RECT  2.140 0.440 2.420 0.720 ;
        RECT  2.240 1.200 2.300 1.480 ;
        RECT  2.080 1.200 2.240 1.900 ;
        RECT  1.850 1.740 2.080 1.900 ;
        RECT  1.690 1.740 1.850 3.130 ;
        RECT  0.930 2.480 1.690 2.640 ;
        RECT  1.220 0.880 1.380 2.030 ;
        RECT  1.110 0.880 1.220 1.040 ;
        RECT  1.050 1.870 1.220 2.030 ;
        RECT  0.950 0.440 1.110 1.040 ;
        RECT  0.790 1.430 1.060 1.710 ;
        RECT  0.830 1.870 1.050 2.190 ;
        RECT  0.780 0.440 0.950 0.660 ;
        RECT  0.670 2.480 0.930 3.130 ;
        RECT  0.670 1.030 0.790 1.710 ;
        RECT  0.650 1.030 0.670 3.130 ;
        RECT  0.510 1.030 0.650 2.640 ;
    END
END TLATNCAX2TR

MACRO TLATNCAX20TR
    CLASS CORE ;
    FOREIGN TLATNCAX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.230 1.610 17.510 3.160 ;
        RECT  16.720 1.610 17.230 2.500 ;
        RECT  16.070 0.760 16.720 2.500 ;
        RECT  15.790 0.760 16.070 3.010 ;
        RECT  15.680 0.760 15.790 2.830 ;
        RECT  13.790 0.500 15.680 1.430 ;
        RECT  15.110 1.910 15.680 2.830 ;
        RECT  14.830 1.910 15.110 3.160 ;
        RECT  14.150 1.910 14.830 2.830 ;
        RECT  13.870 1.910 14.150 3.160 ;
        RECT  13.190 1.910 13.870 2.830 ;
        RECT  13.510 0.440 13.790 1.430 ;
        RECT  12.750 0.500 13.510 1.430 ;
        RECT  12.910 1.910 13.190 3.160 ;
        RECT  12.230 1.910 12.910 2.830 ;
        RECT  12.470 0.440 12.750 1.430 ;
        RECT  11.710 0.500 12.470 1.430 ;
        RECT  11.950 1.910 12.230 3.160 ;
        RECT  11.270 1.910 11.950 2.830 ;
        RECT  11.430 0.440 11.710 1.430 ;
        RECT  10.670 0.500 11.430 1.430 ;
        RECT  10.990 1.910 11.270 3.160 ;
        RECT  10.310 1.910 10.990 2.830 ;
        RECT  10.390 0.440 10.670 1.430 ;
        RECT  10.030 1.910 10.310 3.160 ;
        END
        ANTENNADIFFAREA 28.466 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.960 1.660 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.600 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.310 -0.280 17.600 0.280 ;
        RECT  14.030 -0.280 14.310 0.340 ;
        RECT  13.270 -0.280 14.030 0.280 ;
        RECT  12.990 -0.280 13.270 0.340 ;
        RECT  12.230 -0.280 12.990 0.280 ;
        RECT  11.950 -0.280 12.230 0.340 ;
        RECT  11.190 -0.280 11.950 0.280 ;
        RECT  10.910 -0.280 11.190 0.340 ;
        RECT  10.190 -0.280 10.910 0.280 ;
        RECT  9.870 -0.280 10.190 0.990 ;
        RECT  9.190 -0.280 9.870 0.340 ;
        RECT  8.910 -0.280 9.190 0.400 ;
        RECT  8.270 -0.280 8.910 0.340 ;
        RECT  7.990 -0.280 8.270 0.400 ;
        RECT  7.350 -0.280 7.990 0.340 ;
        RECT  7.070 -0.280 7.350 0.400 ;
        RECT  3.220 -0.280 7.070 0.340 ;
        RECT  1.820 -0.280 3.220 0.280 ;
        RECT  0.800 -0.280 1.820 0.400 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.030 3.320 17.600 3.880 ;
        RECT  16.270 2.730 17.030 3.880 ;
        RECT  15.590 3.320 16.270 3.880 ;
        RECT  15.310 2.990 15.590 3.880 ;
        RECT  14.630 3.320 15.310 3.880 ;
        RECT  14.350 2.990 14.630 3.880 ;
        RECT  13.670 3.320 14.350 3.880 ;
        RECT  13.390 2.990 13.670 3.880 ;
        RECT  12.710 3.320 13.390 3.880 ;
        RECT  12.430 2.990 12.710 3.880 ;
        RECT  11.750 3.320 12.430 3.880 ;
        RECT  11.470 2.990 11.750 3.880 ;
        RECT  10.790 3.320 11.470 3.880 ;
        RECT  10.510 2.990 10.790 3.880 ;
        RECT  9.830 3.320 10.510 3.880 ;
        RECT  9.550 1.930 9.830 3.880 ;
        RECT  8.870 3.320 9.550 3.880 ;
        RECT  8.590 2.250 8.870 3.880 ;
        RECT  7.910 3.320 8.590 3.880 ;
        RECT  7.630 2.250 7.910 3.880 ;
        RECT  6.950 3.320 7.630 3.880 ;
        RECT  6.670 2.420 6.950 3.880 ;
        RECT  5.250 3.320 6.670 3.880 ;
        RECT  4.970 3.200 5.250 3.880 ;
        RECT  3.500 3.260 4.970 3.880 ;
        RECT  3.220 3.200 3.500 3.880 ;
        RECT  1.820 3.320 3.220 3.880 ;
        RECT  0.760 2.800 1.820 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.390 1.590 15.310 1.750 ;
        RECT  9.390 0.990 9.710 1.270 ;
        RECT  9.230 0.990 9.390 3.160 ;
        RECT  7.590 0.990 9.230 1.270 ;
        RECT  9.070 1.930 9.230 3.160 ;
        RECT  7.350 1.490 9.070 1.770 ;
        RECT  8.390 1.930 9.070 2.090 ;
        RECT  8.110 1.930 8.390 3.160 ;
        RECT  7.430 1.930 8.110 2.090 ;
        RECT  7.150 1.930 7.430 3.160 ;
        RECT  7.190 0.780 7.350 1.770 ;
        RECT  6.590 0.780 7.190 1.060 ;
        RECT  6.910 1.220 7.030 1.500 ;
        RECT  6.750 1.220 6.910 2.260 ;
        RECT  6.410 2.100 6.750 2.260 ;
        RECT  6.430 0.780 6.590 1.940 ;
        RECT  6.090 1.780 6.430 1.940 ;
        RECT  6.250 2.100 6.410 3.040 ;
        RECT  6.050 0.500 6.270 1.620 ;
        RECT  5.570 2.880 6.250 3.040 ;
        RECT  5.890 1.780 6.090 2.720 ;
        RECT  4.360 0.500 6.050 0.660 ;
        RECT  5.810 0.820 5.890 2.720 ;
        RECT  5.730 0.820 5.810 1.940 ;
        RECT  5.590 0.820 5.730 1.100 ;
        RECT  5.290 1.260 5.570 3.040 ;
        RECT  4.160 2.880 5.290 3.040 ;
        RECT  4.970 1.050 5.130 2.090 ;
        RECT  4.520 1.050 4.970 1.330 ;
        RECT  4.800 1.930 4.970 2.090 ;
        RECT  4.360 1.490 4.810 1.770 ;
        RECT  4.600 1.930 4.800 2.190 ;
        RECT  4.320 1.930 4.600 2.610 ;
        RECT  4.200 0.500 4.360 1.770 ;
        RECT  3.840 0.500 4.200 0.660 ;
        RECT  3.650 1.610 4.200 1.770 ;
        RECT  4.000 2.000 4.160 3.040 ;
        RECT  3.180 1.090 4.040 1.370 ;
        RECT  3.810 2.000 4.000 2.280 ;
        RECT  2.140 2.880 4.000 3.040 ;
        RECT  3.560 0.500 3.840 0.930 ;
        RECT  3.650 2.440 3.840 2.720 ;
        RECT  3.490 1.610 3.650 2.720 ;
        RECT  2.660 0.500 3.560 0.660 ;
        RECT  2.660 2.560 3.490 2.720 ;
        RECT  3.020 1.090 3.180 2.100 ;
        RECT  2.280 1.820 3.020 2.100 ;
        RECT  2.280 1.380 2.860 1.660 ;
        RECT  2.440 0.500 2.660 0.990 ;
        RECT  2.440 2.440 2.660 2.720 ;
        RECT  2.120 0.680 2.280 1.660 ;
        RECT  2.120 1.820 2.280 2.210 ;
        RECT  1.980 2.370 2.140 3.040 ;
        RECT  1.040 0.680 2.120 0.840 ;
        RECT  1.480 2.050 2.120 2.210 ;
        RECT  1.040 2.370 1.980 2.530 ;
        RECT  1.320 1.000 1.480 2.210 ;
        RECT  1.200 1.000 1.320 1.310 ;
        RECT  1.200 1.930 1.320 2.210 ;
        RECT  1.040 1.470 1.160 1.750 ;
        RECT  0.880 0.680 1.040 2.530 ;
        RECT  0.560 1.170 0.880 1.330 ;
        RECT  0.560 2.370 0.880 2.530 ;
        RECT  0.280 0.500 0.560 1.330 ;
        RECT  0.280 2.120 0.560 3.160 ;
    END
END TLATNCAX20TR

MACRO TLATNCAX16TR
    CLASS CORE ;
    FOREIGN TLATNCAX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.510 0.500 14.720 2.490 ;
        RECT  13.570 0.500 14.510 2.830 ;
        RECT  9.200 0.500 13.570 1.420 ;
        RECT  13.540 1.910 13.570 2.830 ;
        RECT  13.380 1.910 13.540 3.160 ;
        RECT  12.580 1.910 13.380 2.830 ;
        RECT  12.420 1.910 12.580 3.160 ;
        RECT  11.620 1.910 12.420 2.830 ;
        RECT  11.460 1.910 11.620 3.160 ;
        RECT  10.660 1.910 11.460 2.830 ;
        RECT  10.500 1.910 10.660 3.160 ;
        RECT  9.700 1.910 10.500 2.830 ;
        RECT  9.540 1.910 9.700 3.160 ;
        RECT  8.740 1.910 9.540 2.830 ;
        RECT  8.580 1.910 8.740 3.160 ;
        END
        ANTENNADIFFAREA 23.768 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.240 1.920 1.620 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.580 1.640 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.120 -0.280 15.200 0.280 ;
        RECT  12.840 -0.280 13.120 0.340 ;
        RECT  12.080 -0.280 12.840 0.280 ;
        RECT  11.800 -0.280 12.080 0.340 ;
        RECT  11.040 -0.280 11.800 0.280 ;
        RECT  10.760 -0.280 11.040 0.340 ;
        RECT  10.000 -0.280 10.760 0.280 ;
        RECT  9.720 -0.280 10.000 0.340 ;
        RECT  8.940 -0.280 9.720 0.280 ;
        RECT  8.700 -0.280 8.940 0.990 ;
        RECT  7.920 -0.280 8.700 0.280 ;
        RECT  7.640 -0.280 7.920 0.880 ;
        RECT  6.880 -0.280 7.640 0.280 ;
        RECT  6.600 -0.280 6.880 0.880 ;
        RECT  5.890 -0.280 6.600 0.280 ;
        RECT  5.630 -0.280 5.890 1.260 ;
        RECT  4.900 -0.280 5.630 0.280 ;
        RECT  4.620 -0.280 4.900 0.340 ;
        RECT  3.860 -0.280 4.620 0.280 ;
        RECT  3.180 -0.280 3.860 0.340 ;
        RECT  1.560 -0.280 3.180 0.280 ;
        RECT  0.700 -0.280 1.560 0.760 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.970 3.320 15.200 3.880 ;
        RECT  14.720 2.880 14.970 3.880 ;
        RECT  14.120 3.320 14.720 3.880 ;
        RECT  13.840 3.260 14.120 3.880 ;
        RECT  13.120 3.320 13.840 3.880 ;
        RECT  12.840 2.990 13.120 3.880 ;
        RECT  12.160 3.320 12.840 3.880 ;
        RECT  11.880 2.990 12.160 3.880 ;
        RECT  11.200 3.320 11.880 3.880 ;
        RECT  10.920 2.990 11.200 3.880 ;
        RECT  10.240 3.320 10.920 3.880 ;
        RECT  9.960 2.990 10.240 3.880 ;
        RECT  9.280 3.320 9.960 3.880 ;
        RECT  9.000 2.990 9.280 3.880 ;
        RECT  8.340 3.320 9.000 3.880 ;
        RECT  8.030 2.130 8.340 3.880 ;
        RECT  7.370 3.320 8.030 3.880 ;
        RECT  7.070 2.130 7.370 3.880 ;
        RECT  6.410 3.320 7.070 3.880 ;
        RECT  6.100 2.310 6.410 3.880 ;
        RECT  5.630 3.320 6.100 3.880 ;
        RECT  5.260 2.610 5.630 3.880 ;
        RECT  3.910 3.320 5.260 3.880 ;
        RECT  3.360 3.220 3.910 3.880 ;
        RECT  1.510 3.320 3.360 3.880 ;
        RECT  1.510 2.730 1.660 2.950 ;
        RECT  1.100 2.730 1.510 3.880 ;
        RECT  0.960 2.730 1.100 2.950 ;
        RECT  0.000 3.320 1.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.440 1.580 13.010 1.740 ;
        RECT  8.320 1.040 8.440 1.740 ;
        RECT  8.160 1.040 8.320 1.970 ;
        RECT  6.080 1.040 8.160 1.200 ;
        RECT  7.780 1.810 8.160 1.970 ;
        RECT  5.360 1.490 8.000 1.650 ;
        RECT  7.620 1.810 7.780 3.160 ;
        RECT  6.820 1.810 7.620 1.970 ;
        RECT  6.660 1.810 6.820 3.160 ;
        RECT  5.920 1.810 6.660 1.970 ;
        RECT  5.640 1.810 5.920 2.140 ;
        RECT  5.200 0.980 5.360 1.930 ;
        RECT  4.720 1.770 5.200 1.930 ;
        RECT  4.600 0.600 4.760 1.610 ;
        RECT  4.560 1.770 4.720 2.890 ;
        RECT  2.960 0.600 4.600 0.760 ;
        RECT  4.440 1.770 4.560 1.930 ;
        RECT  4.280 1.040 4.440 1.930 ;
        RECT  4.100 1.040 4.280 1.200 ;
        RECT  3.960 1.580 4.120 2.920 ;
        RECT  2.860 2.760 3.960 2.920 ;
        RECT  3.640 1.100 3.800 2.070 ;
        RECT  3.360 1.100 3.640 1.260 ;
        RECT  3.360 1.910 3.640 2.070 ;
        RECT  2.960 1.420 3.480 1.700 ;
        RECT  3.200 0.980 3.360 1.260 ;
        RECT  3.120 1.910 3.360 2.600 ;
        RECT  2.800 0.600 2.960 2.280 ;
        RECT  2.700 2.760 2.860 3.160 ;
        RECT  2.400 0.600 2.800 0.760 ;
        RECT  2.540 2.120 2.800 2.280 ;
        RECT  2.100 3.000 2.700 3.160 ;
        RECT  2.480 0.920 2.640 1.960 ;
        RECT  2.260 2.120 2.540 2.760 ;
        RECT  1.260 0.920 2.480 1.080 ;
        RECT  2.240 0.480 2.400 0.760 ;
        RECT  2.100 1.280 2.280 1.940 ;
        RECT  2.080 1.280 2.100 3.160 ;
        RECT  1.940 1.780 2.080 3.160 ;
        RECT  0.940 2.370 1.940 2.530 ;
        RECT  1.100 0.920 1.260 2.210 ;
        RECT  0.800 0.920 0.940 2.530 ;
        RECT  0.780 0.920 0.800 2.950 ;
        RECT  0.320 0.920 0.780 1.080 ;
        RECT  0.640 2.330 0.780 2.950 ;
        RECT  0.100 2.680 0.640 2.950 ;
        RECT  0.160 0.650 0.320 1.080 ;
    END
END TLATNCAX16TR

MACRO TLATNCAX12TR
    CLASS CORE ;
    FOREIGN TLATNCAX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.040 0.500 12.280 3.160 ;
        RECT  11.480 0.500 12.040 2.550 ;
        RECT  7.010 0.500 11.480 1.220 ;
        RECT  11.350 1.830 11.480 2.550 ;
        RECT  11.040 1.830 11.350 3.160 ;
        RECT  10.410 1.830 11.040 2.550 ;
        RECT  10.100 1.830 10.410 3.160 ;
        RECT  9.430 1.830 10.100 2.550 ;
        RECT  9.140 1.830 9.430 3.160 ;
        RECT  8.490 1.830 9.140 2.550 ;
        RECT  8.190 1.830 8.490 3.160 ;
        RECT  7.520 1.830 8.190 2.550 ;
        RECT  7.230 1.830 7.520 3.160 ;
        END
        ANTENNADIFFAREA 18.944 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.320 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.2352 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.910 -0.280 12.400 0.280 ;
        RECT  11.630 -0.280 11.910 0.340 ;
        RECT  10.870 -0.280 11.630 0.280 ;
        RECT  10.590 -0.280 10.870 0.330 ;
        RECT  9.890 -0.280 10.590 0.280 ;
        RECT  9.610 -0.280 9.890 0.340 ;
        RECT  8.850 -0.280 9.610 0.280 ;
        RECT  8.570 -0.280 8.850 0.340 ;
        RECT  7.810 -0.280 8.570 0.280 ;
        RECT  7.530 -0.280 7.810 0.340 ;
        RECT  6.750 -0.280 7.530 0.280 ;
        RECT  6.590 -0.280 6.750 1.010 ;
        RECT  5.850 -0.280 6.590 0.280 ;
        RECT  5.570 -0.280 5.850 0.850 ;
        RECT  4.900 -0.280 5.570 0.280 ;
        RECT  4.620 -0.280 4.900 0.340 ;
        RECT  3.860 -0.280 4.620 0.280 ;
        RECT  3.190 -0.280 3.860 0.340 ;
        RECT  1.630 -0.280 3.190 0.280 ;
        RECT  1.350 -0.280 1.630 0.340 ;
        RECT  0.890 -0.280 1.350 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.840 3.320 12.400 3.880 ;
        RECT  11.530 2.930 11.840 3.880 ;
        RECT  10.880 3.320 11.530 3.880 ;
        RECT  10.590 2.930 10.880 3.880 ;
        RECT  9.900 3.320 10.590 3.880 ;
        RECT  9.640 2.930 9.900 3.880 ;
        RECT  8.970 3.320 9.640 3.880 ;
        RECT  8.660 2.930 8.970 3.880 ;
        RECT  8.000 3.320 8.660 3.880 ;
        RECT  7.690 2.930 8.000 3.880 ;
        RECT  7.030 3.320 7.690 3.880 ;
        RECT  6.730 2.070 7.030 3.880 ;
        RECT  6.080 3.320 6.730 3.880 ;
        RECT  5.780 2.220 6.080 3.880 ;
        RECT  5.090 3.320 5.780 3.880 ;
        RECT  4.780 2.350 5.090 3.880 ;
        RECT  3.750 3.320 4.780 3.880 ;
        RECT  3.470 3.240 3.750 3.880 ;
        RECT  1.590 3.320 3.470 3.880 ;
        RECT  0.900 2.850 1.590 3.880 ;
        RECT  0.000 3.320 0.900 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.490 1.380 11.110 1.540 ;
        RECT  6.390 1.380 6.490 3.160 ;
        RECT  6.330 1.010 6.390 3.160 ;
        RECT  6.230 1.010 6.330 2.060 ;
        RECT  5.090 1.010 6.230 1.170 ;
        RECT  5.530 1.900 6.230 2.060 ;
        RECT  4.530 1.580 6.070 1.740 ;
        RECT  5.370 1.900 5.530 3.160 ;
        RECT  4.700 1.260 4.820 1.420 ;
        RECT  4.540 0.550 4.700 1.420 ;
        RECT  2.930 0.550 4.540 0.710 ;
        RECT  4.380 1.580 4.530 3.020 ;
        RECT  4.370 0.870 4.380 3.020 ;
        RECT  4.220 0.870 4.370 1.740 ;
        RECT  4.100 0.870 4.220 1.030 ;
        RECT  3.850 1.210 4.010 2.910 ;
        RECT  2.650 2.750 3.850 2.910 ;
        RECT  3.530 0.990 3.690 2.130 ;
        RECT  3.290 0.990 3.530 1.150 ;
        RECT  3.050 1.970 3.530 2.130 ;
        RECT  2.930 1.400 3.370 1.680 ;
        RECT  3.130 0.870 3.290 1.150 ;
        RECT  2.890 1.970 3.050 2.560 ;
        RECT  2.770 0.550 2.930 1.800 ;
        RECT  2.410 0.550 2.770 0.710 ;
        RECT  2.330 1.640 2.770 1.800 ;
        RECT  2.490 2.750 2.650 3.160 ;
        RECT  2.450 0.960 2.610 1.480 ;
        RECT  2.010 3.000 2.490 3.160 ;
        RECT  1.120 0.960 2.450 1.120 ;
        RECT  2.250 0.440 2.410 0.720 ;
        RECT  2.170 1.640 2.330 2.330 ;
        RECT  2.010 1.320 2.270 1.480 ;
        RECT  1.850 1.320 2.010 3.160 ;
        RECT  0.770 2.530 1.850 2.690 ;
        RECT  1.120 2.130 1.250 2.290 ;
        RECT  0.960 0.960 1.120 2.290 ;
        RECT  0.770 0.560 1.110 0.720 ;
        RECT  0.610 0.560 0.770 2.690 ;
        RECT  0.150 0.560 0.610 0.860 ;
        RECT  0.310 2.530 0.610 2.690 ;
        RECT  0.150 2.530 0.310 2.910 ;
    END
END TLATNCAX12TR

MACRO TLATNXLTR
    CLASS CORE ;
    FOREIGN TLATNXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.560 0.920 4.720 2.760 ;
        RECT  4.320 0.920 4.560 1.200 ;
        RECT  4.480 1.640 4.560 2.760 ;
        RECT  4.260 2.440 4.480 2.760 ;
        END
        ANTENNADIFFAREA 1.202 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.360 4.320 2.280 ;
        RECT  4.100 1.360 4.160 1.520 ;
        RECT  4.080 2.120 4.160 2.280 ;
        RECT  3.940 0.690 4.100 1.520 ;
        RECT  3.920 2.120 4.080 2.880 ;
        RECT  3.840 0.690 3.940 0.850 ;
        RECT  3.640 2.720 3.920 2.880 ;
        RECT  3.560 0.570 3.840 0.850 ;
        RECT  3.280 2.720 3.640 3.160 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.470 0.490 1.750 ;
        RECT  0.320 1.470 0.360 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.420 1.450 1.960 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.510 -0.280 4.800 0.280 ;
        RECT  4.230 -0.280 4.510 0.400 ;
        RECT  3.180 -0.280 4.230 0.280 ;
        RECT  2.900 -0.280 3.180 1.230 ;
        RECT  1.390 -0.280 2.900 0.280 ;
        RECT  1.110 -0.280 1.390 0.400 ;
        RECT  0.370 -0.280 1.110 0.280 ;
        RECT  0.090 -0.280 0.370 0.650 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 3.320 4.800 3.880 ;
        RECT  3.860 3.200 4.140 3.880 ;
        RECT  3.110 3.320 3.860 3.880 ;
        RECT  2.830 2.800 3.110 3.880 ;
        RECT  1.540 3.260 2.830 3.880 ;
        RECT  1.260 2.880 1.540 3.880 ;
        RECT  0.370 3.320 1.260 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.780 1.680 4.000 1.960 ;
        RECT  3.760 1.030 3.780 1.960 ;
        RECT  3.600 1.030 3.760 2.400 ;
        RECT  2.900 2.120 3.600 2.400 ;
        RECT  3.060 1.470 3.340 1.750 ;
        RECT  2.740 1.470 3.060 1.630 ;
        RECT  2.740 1.790 2.900 2.400 ;
        RECT  2.580 0.590 2.740 1.630 ;
        RECT  2.620 1.790 2.740 2.070 ;
        RECT  1.980 0.590 2.580 0.870 ;
        RECT  2.280 1.470 2.580 1.630 ;
        RECT  2.140 1.030 2.420 1.310 ;
        RECT  2.120 1.470 2.280 2.400 ;
        RECT  1.260 1.030 2.140 1.190 ;
        RECT  1.980 2.120 2.120 2.400 ;
        RECT  1.260 2.560 2.020 2.720 ;
        RECT  1.100 0.690 1.260 2.720 ;
        RECT  0.830 0.690 1.100 0.850 ;
        RECT  0.580 2.500 1.100 2.720 ;
        RECT  0.820 2.880 1.100 3.160 ;
        RECT  0.660 1.030 0.940 2.280 ;
        RECT  0.550 0.570 0.830 0.850 ;
        RECT  0.420 2.880 0.820 3.040 ;
        RECT  0.530 1.030 0.660 1.310 ;
        RECT  0.570 1.910 0.660 2.280 ;
        RECT  0.420 2.120 0.570 2.280 ;
        RECT  0.260 2.120 0.420 3.040 ;
    END
END TLATNXLTR

MACRO TLATNX4TR
    CLASS CORE ;
    FOREIGN TLATNX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.040 6.720 1.760 ;
        RECT  6.630 1.040 6.670 2.130 ;
        RECT  6.430 0.500 6.630 3.160 ;
        RECT  6.350 0.500 6.430 1.310 ;
        RECT  6.350 1.970 6.430 3.160 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.490 5.670 2.250 ;
        RECT  5.280 1.440 5.390 2.160 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.450 2.360 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 0.790 3.400 1.590 ;
        RECT  1.920 0.790 3.180 0.950 ;
        RECT  1.740 0.790 1.920 1.620 ;
        RECT  1.620 1.240 1.740 1.620 ;
        END
        ANTENNAGATEAREA 0.5088 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 -0.280 7.200 0.280 ;
        RECT  6.880 -0.280 7.110 1.310 ;
        RECT  6.830 -0.280 6.880 0.880 ;
        RECT  6.150 -0.280 6.830 0.280 ;
        RECT  5.870 -0.280 6.150 1.310 ;
        RECT  5.150 -0.280 5.870 0.280 ;
        RECT  4.870 -0.280 5.150 0.400 ;
        RECT  3.360 -0.280 4.870 0.280 ;
        RECT  3.080 -0.280 3.360 0.310 ;
        RECT  1.720 -0.280 3.080 0.280 ;
        RECT  1.400 -0.280 1.720 0.620 ;
        RECT  0.370 -0.280 1.400 0.280 ;
        RECT  0.090 -0.280 0.370 1.050 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.320 7.200 3.880 ;
        RECT  6.830 1.970 7.110 3.880 ;
        RECT  6.150 3.320 6.830 3.880 ;
        RECT  5.870 2.930 6.150 3.880 ;
        RECT  5.150 3.320 5.870 3.880 ;
        RECT  4.870 3.180 5.150 3.880 ;
        RECT  3.360 3.320 4.870 3.880 ;
        RECT  3.080 2.860 3.360 3.880 ;
        RECT  1.660 3.320 3.080 3.880 ;
        RECT  1.380 3.200 1.660 3.880 ;
        RECT  0.370 3.320 1.380 3.880 ;
        RECT  0.090 2.750 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 1.530 6.270 1.810 ;
        RECT  5.990 1.530 6.150 2.770 ;
        RECT  4.790 2.610 5.990 2.770 ;
        RECT  4.960 1.210 5.120 2.130 ;
        RECT  4.690 1.210 4.960 1.370 ;
        RECT  4.790 1.970 4.960 2.130 ;
        RECT  4.350 1.530 4.800 1.810 ;
        RECT  4.670 1.970 4.790 2.770 ;
        RECT  4.530 0.450 4.690 1.370 ;
        RECT  4.510 1.970 4.670 3.100 ;
        RECT  4.090 0.450 4.530 0.610 ;
        RECT  4.060 2.820 4.510 3.100 ;
        RECT  4.340 1.530 4.350 2.630 ;
        RECT  4.180 0.900 4.340 2.630 ;
        RECT  3.770 0.900 4.180 1.060 ;
        RECT  2.520 2.440 4.180 2.630 ;
        RECT  3.720 2.090 4.020 2.280 ;
        RECT  3.850 1.300 4.010 1.930 ;
        RECT  3.550 1.770 3.850 1.930 ;
        RECT  3.610 0.470 3.770 1.060 ;
        RECT  2.700 2.120 3.720 2.280 ;
        RECT  2.200 0.470 3.610 0.630 ;
        RECT  3.380 1.770 3.550 1.960 ;
        RECT  3.020 1.800 3.380 1.960 ;
        RECT  2.860 1.110 3.020 1.960 ;
        RECT  2.260 1.110 2.860 1.270 ;
        RECT  2.460 1.430 2.700 2.280 ;
        RECT  2.240 2.440 2.520 3.160 ;
        RECT  1.780 2.120 2.460 2.280 ;
        RECT  2.100 1.110 2.260 1.960 ;
        RECT  1.420 1.800 2.100 1.960 ;
        RECT  1.620 2.120 1.780 2.630 ;
        RECT  0.920 2.470 1.620 2.630 ;
        RECT  1.260 0.900 1.420 2.290 ;
        RECT  1.160 0.900 1.260 1.060 ;
        RECT  1.020 2.010 1.260 2.290 ;
        RECT  1.000 0.440 1.160 1.060 ;
        RECT  0.840 1.560 1.080 1.810 ;
        RECT  0.800 2.470 0.920 2.750 ;
        RECT  0.800 0.980 0.840 1.810 ;
        RECT  0.640 0.980 0.800 2.750 ;
    END
END TLATNX4TR

MACRO TLATNX2TR
    CLASS CORE ;
    FOREIGN TLATNX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.360 0.440 5.520 3.160 ;
        RECT  5.280 0.440 5.360 1.560 ;
        RECT  5.290 1.910 5.360 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.560 1.240 4.720 1.560 ;
        RECT  4.330 1.240 4.560 3.160 ;
        RECT  4.270 1.030 4.330 3.160 ;
        RECT  4.170 1.030 4.270 1.400 ;
        END
        ANTENNADIFFAREA 3.744 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.440 0.460 1.260 ;
        RECT  0.080 0.440 0.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.720 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 -0.280 5.600 0.280 ;
        RECT  4.810 -0.280 4.970 0.670 ;
        RECT  3.380 -0.280 4.810 0.280 ;
        RECT  3.080 -0.280 3.380 1.100 ;
        RECT  1.660 -0.280 3.080 0.280 ;
        RECT  1.380 -0.280 1.660 0.340 ;
        RECT  0.000 -0.280 1.380 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.030 3.320 5.600 3.880 ;
        RECT  4.750 1.910 5.030 3.880 ;
        RECT  3.440 3.320 4.750 3.880 ;
        RECT  3.130 2.310 3.440 3.880 ;
        RECT  1.580 3.320 3.130 3.880 ;
        RECT  1.300 3.260 1.580 3.880 ;
        RECT  0.440 3.320 1.300 3.880 ;
        RECT  0.160 2.800 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.960 0.830 5.120 1.750 ;
        RECT  4.650 0.830 4.960 0.990 ;
        RECT  4.900 1.450 4.960 1.750 ;
        RECT  4.490 0.630 4.650 0.990 ;
        RECT  4.010 0.630 4.490 0.790 ;
        RECT  3.850 0.630 4.010 2.450 ;
        RECT  3.710 0.630 3.850 1.500 ;
        RECT  3.690 2.170 3.850 2.450 ;
        RECT  3.080 1.340 3.710 1.500 ;
        RECT  2.920 1.740 3.690 1.900 ;
        RECT  2.760 0.560 2.920 2.760 ;
        RECT  2.440 0.560 2.760 0.720 ;
        RECT  2.360 2.600 2.760 2.760 ;
        RECT  2.440 2.160 2.600 2.440 ;
        RECT  2.410 0.920 2.570 2.000 ;
        RECT  2.280 0.440 2.440 0.720 ;
        RECT  2.240 2.160 2.440 2.320 ;
        RECT  1.520 0.920 2.410 1.080 ;
        RECT  2.200 2.600 2.360 2.880 ;
        RECT  2.080 1.280 2.240 2.320 ;
        RECT  1.840 2.160 2.080 2.320 ;
        RECT  1.680 2.160 1.840 2.910 ;
        RECT  0.780 2.750 1.680 2.910 ;
        RECT  1.360 0.920 1.520 2.590 ;
        RECT  0.940 1.070 1.360 1.230 ;
        RECT  0.940 2.430 1.360 2.590 ;
        RECT  0.780 1.510 1.200 1.790 ;
        RECT  0.780 0.530 0.900 0.830 ;
        RECT  0.620 0.530 0.780 2.910 ;
    END
END TLATNX2TR

MACRO TLATNX1TR
    CLASS CORE ;
    FOREIGN TLATNX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 1.560 4.720 2.760 ;
        RECT  4.420 0.600 4.700 2.760 ;
        END
        ANTENNADIFFAREA 2.174 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.100 0.670 4.260 2.600 ;
        RECT  3.700 0.670 4.100 0.830 ;
        RECT  3.560 2.440 4.100 2.600 ;
        RECT  3.420 0.550 3.700 0.830 ;
        RECT  3.270 2.440 3.560 2.950 ;
        END
        ANTENNADIFFAREA 1.86 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.500 0.430 1.780 ;
        RECT  0.320 1.500 0.360 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.220 1.960 1.600 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.280 4.800 0.280 ;
        RECT  4.010 -0.280 4.290 0.360 ;
        RECT  3.160 -0.280 4.010 0.280 ;
        RECT  2.920 -0.280 3.160 0.820 ;
        RECT  1.420 -0.280 2.920 0.280 ;
        RECT  1.120 -0.280 1.420 0.590 ;
        RECT  0.370 -0.280 1.120 0.280 ;
        RECT  0.090 -0.280 0.370 0.640 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 3.320 4.800 3.880 ;
        RECT  3.840 2.910 4.170 3.880 ;
        RECT  3.080 3.320 3.840 3.880 ;
        RECT  2.780 2.800 3.080 3.880 ;
        RECT  1.540 3.320 2.780 3.880 ;
        RECT  1.260 2.930 1.540 3.880 ;
        RECT  0.370 3.320 1.260 3.880 ;
        RECT  0.090 3.240 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.700 1.410 3.940 1.690 ;
        RECT  3.580 1.010 3.700 1.690 ;
        RECT  3.420 1.010 3.580 2.270 ;
        RECT  2.820 1.990 3.420 2.270 ;
        RECT  3.040 1.380 3.260 1.660 ;
        RECT  2.760 1.380 3.040 1.540 ;
        RECT  2.660 1.720 2.820 2.270 ;
        RECT  2.600 0.580 2.760 1.540 ;
        RECT  2.540 1.720 2.660 1.940 ;
        RECT  2.260 0.580 2.600 0.740 ;
        RECT  2.280 1.340 2.600 1.540 ;
        RECT  2.220 0.900 2.440 1.180 ;
        RECT  2.120 1.340 2.280 2.170 ;
        RECT  1.980 0.460 2.260 0.740 ;
        RECT  1.220 0.900 2.220 1.060 ;
        RECT  1.900 1.890 2.120 2.170 ;
        RECT  1.860 2.660 1.980 2.940 ;
        RECT  1.700 2.540 1.860 2.940 ;
        RECT  1.220 2.540 1.700 2.750 ;
        RECT  1.060 0.750 1.220 2.750 ;
        RECT  0.820 2.920 1.100 3.160 ;
        RECT  0.830 0.750 1.060 0.910 ;
        RECT  0.620 2.480 1.060 2.750 ;
        RECT  0.620 1.070 0.900 2.290 ;
        RECT  0.550 0.550 0.830 0.910 ;
        RECT  0.420 2.920 0.820 3.080 ;
        RECT  0.530 1.070 0.620 1.290 ;
        RECT  0.510 2.030 0.620 2.290 ;
        RECT  0.420 2.130 0.510 2.290 ;
        RECT  0.260 2.130 0.420 3.080 ;
    END
END TLATNX1TR

MACRO TLATXLTR
    CLASS CORE ;
    FOREIGN TLATXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.030 1.010 4.320 3.090 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.710 0.670 3.870 2.510 ;
        RECT  3.520 0.670 3.710 0.830 ;
        RECT  3.560 2.350 3.710 2.510 ;
        RECT  3.130 2.350 3.560 2.760 ;
        RECT  3.240 0.550 3.520 0.830 ;
        END
        ANTENNADIFFAREA 1.09 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.440 0.480 1.720 ;
        RECT  0.320 1.440 0.360 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.180 1.960 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.070 -0.280 4.400 0.280 ;
        RECT  3.790 -0.280 4.070 0.400 ;
        RECT  2.950 -0.280 3.790 0.280 ;
        RECT  2.630 -0.280 2.950 0.400 ;
        RECT  1.390 -0.280 2.630 0.280 ;
        RECT  1.110 -0.280 1.390 0.400 ;
        RECT  0.370 -0.280 1.110 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 3.320 4.400 3.880 ;
        RECT  3.550 2.930 3.830 3.880 ;
        RECT  3.160 3.320 3.550 3.880 ;
        RECT  2.880 3.200 3.160 3.880 ;
        RECT  1.470 3.320 2.880 3.880 ;
        RECT  1.190 2.880 1.470 3.880 ;
        RECT  0.370 3.320 1.190 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.390 1.010 3.550 2.170 ;
        RECT  3.240 1.010 3.390 1.290 ;
        RECT  2.680 1.890 3.390 2.170 ;
        RECT  2.320 1.450 3.110 1.730 ;
        RECT  2.520 1.890 2.680 3.160 ;
        RECT  2.400 2.900 2.520 3.160 ;
        RECT  2.160 0.440 2.320 2.400 ;
        RECT  1.960 2.560 2.240 2.840 ;
        RECT  2.040 0.440 2.160 0.720 ;
        RECT  1.840 2.120 2.160 2.400 ;
        RECT  1.180 2.560 1.960 2.720 ;
        RECT  1.600 0.440 1.880 0.810 ;
        RECT  1.180 0.650 1.600 0.810 ;
        RECT  1.020 0.650 1.180 2.720 ;
        RECT  0.750 2.880 1.030 3.160 ;
        RECT  0.830 0.650 1.020 0.810 ;
        RECT  0.510 2.500 1.020 2.720 ;
        RECT  0.830 1.390 0.860 1.670 ;
        RECT  0.550 0.530 0.830 0.810 ;
        RECT  0.810 0.990 0.830 1.670 ;
        RECT  0.640 0.990 0.810 2.280 ;
        RECT  0.350 2.880 0.750 3.040 ;
        RECT  0.550 0.990 0.640 1.270 ;
        RECT  0.530 1.910 0.640 2.280 ;
        RECT  0.350 2.120 0.530 2.280 ;
        RECT  0.190 2.120 0.350 3.040 ;
    END
END TLATXLTR

MACRO TLATX4TR
    CLASS CORE ;
    FOREIGN TLATX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.040 6.720 1.760 ;
        RECT  6.630 1.040 6.670 2.130 ;
        RECT  6.430 0.540 6.630 3.160 ;
        RECT  6.350 0.540 6.430 1.310 ;
        RECT  6.350 1.970 6.430 3.160 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.540 5.670 2.250 ;
        RECT  5.280 1.440 5.390 2.160 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.480 1.950 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.440 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.432 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 -0.280 7.200 0.280 ;
        RECT  6.830 -0.280 7.110 0.750 ;
        RECT  6.150 -0.280 6.830 0.280 ;
        RECT  5.870 -0.280 6.150 1.310 ;
        RECT  5.150 -0.280 5.870 0.280 ;
        RECT  4.870 -0.280 5.150 0.400 ;
        RECT  3.460 -0.280 4.870 0.280 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  1.740 -0.280 3.180 0.280 ;
        RECT  1.460 -0.280 1.740 0.820 ;
        RECT  0.370 -0.280 1.460 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 3.320 7.200 3.880 ;
        RECT  6.830 1.970 7.110 3.880 ;
        RECT  6.150 3.320 6.830 3.880 ;
        RECT  5.870 2.930 6.150 3.880 ;
        RECT  5.150 3.320 5.870 3.880 ;
        RECT  4.870 3.180 5.150 3.880 ;
        RECT  3.370 3.320 4.870 3.880 ;
        RECT  3.090 3.200 3.370 3.880 ;
        RECT  1.690 3.320 3.090 3.880 ;
        RECT  1.410 3.200 1.690 3.880 ;
        RECT  0.370 3.320 1.410 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 1.530 6.270 1.810 ;
        RECT  5.990 1.530 6.150 2.570 ;
        RECT  5.120 2.410 5.990 2.570 ;
        RECT  4.960 1.320 5.120 2.570 ;
        RECT  4.750 1.320 4.960 1.480 ;
        RECT  4.790 2.410 4.960 2.570 ;
        RECT  4.310 1.640 4.800 1.920 ;
        RECT  4.670 2.290 4.790 2.570 ;
        RECT  4.470 0.560 4.750 1.480 ;
        RECT  4.510 2.290 4.670 3.100 ;
        RECT  4.070 2.880 4.510 3.100 ;
        RECT  3.900 0.560 4.470 0.720 ;
        RECT  4.150 0.910 4.310 2.720 ;
        RECT  2.620 0.910 4.150 1.190 ;
        RECT  2.560 2.440 4.150 2.720 ;
        RECT  3.710 1.360 3.990 2.280 ;
        RECT  3.620 0.500 3.900 0.720 ;
        RECT  2.360 2.120 3.710 2.280 ;
        RECT  2.800 1.680 3.550 1.960 ;
        RECT  2.640 1.350 2.800 1.960 ;
        RECT  2.520 1.350 2.640 1.690 ;
        RECT  2.460 0.710 2.620 1.190 ;
        RECT  2.250 2.440 2.560 3.160 ;
        RECT  2.240 1.350 2.520 1.520 ;
        RECT  2.340 0.710 2.460 0.960 ;
        RECT  2.080 1.750 2.360 2.280 ;
        RECT  2.080 1.120 2.240 1.520 ;
        RECT  1.480 1.120 2.080 1.280 ;
        RECT  1.800 2.120 2.080 2.280 ;
        RECT  1.640 2.120 1.800 2.670 ;
        RECT  0.800 2.510 1.640 2.670 ;
        RECT  1.320 1.120 1.480 2.350 ;
        RECT  1.240 1.120 1.320 1.280 ;
        RECT  1.040 2.070 1.320 2.350 ;
        RECT  1.080 0.540 1.240 1.280 ;
        RECT  0.800 1.530 1.160 1.810 ;
        RECT  0.940 0.540 1.080 0.820 ;
        RECT  0.710 1.010 0.800 2.670 ;
        RECT  0.640 1.010 0.710 2.750 ;
        RECT  0.500 1.010 0.640 1.290 ;
        RECT  0.550 2.110 0.640 2.750 ;
    END
END TLATX4TR

MACRO TLATX2TR
    CLASS CORE ;
    FOREIGN TLATX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 0.440 5.520 3.160 ;
        RECT  5.230 1.910 5.280 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.240 4.720 1.560 ;
        RECT  4.330 1.240 4.550 3.100 ;
        RECT  4.270 1.030 4.330 3.100 ;
        RECT  4.050 1.030 4.270 1.400 ;
        END
        ANTENNADIFFAREA 3.444 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.440 0.450 1.050 ;
        RECT  0.080 0.440 0.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.960 1.640 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.030 -0.280 5.600 0.280 ;
        RECT  4.810 -0.280 5.030 0.670 ;
        RECT  3.470 -0.280 4.810 0.280 ;
        RECT  3.200 -0.280 3.470 1.170 ;
        RECT  1.720 -0.280 3.200 0.280 ;
        RECT  1.440 -0.280 1.720 0.400 ;
        RECT  0.000 -0.280 1.440 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.030 3.320 5.600 3.880 ;
        RECT  4.750 1.910 5.030 3.880 ;
        RECT  3.420 3.260 4.750 3.880 ;
        RECT  3.200 2.230 3.420 3.880 ;
        RECT  1.680 3.260 3.200 3.880 ;
        RECT  1.460 2.480 1.680 3.880 ;
        RECT  0.370 3.320 1.460 3.880 ;
        RECT  0.090 1.910 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.070 1.440 5.120 1.740 ;
        RECT  4.880 0.830 5.070 1.740 ;
        RECT  4.650 0.830 4.880 0.990 ;
        RECT  4.490 0.570 4.650 0.990 ;
        RECT  3.890 0.570 4.490 0.850 ;
        RECT  3.890 2.170 3.910 2.450 ;
        RECT  3.730 0.570 3.890 2.450 ;
        RECT  3.200 1.410 3.730 1.570 ;
        RECT  3.040 1.790 3.570 2.000 ;
        RECT  2.880 0.560 3.040 2.760 ;
        RECT  2.560 0.560 2.880 0.720 ;
        RECT  2.480 2.600 2.880 2.760 ;
        RECT  2.560 0.880 2.720 2.000 ;
        RECT  2.440 2.160 2.720 2.440 ;
        RECT  2.280 0.440 2.560 0.720 ;
        RECT  1.800 0.880 2.560 1.040 ;
        RECT  2.440 1.720 2.560 2.000 ;
        RECT  2.200 2.600 2.480 2.880 ;
        RECT  2.280 2.160 2.440 2.320 ;
        RECT  2.280 1.280 2.400 1.560 ;
        RECT  2.120 1.280 2.280 2.320 ;
        RECT  1.480 2.160 2.120 2.320 ;
        RECT  1.640 0.560 1.800 1.040 ;
        RECT  0.890 0.560 1.640 0.720 ;
        RECT  1.320 1.010 1.480 2.320 ;
        RECT  0.930 1.010 1.320 1.290 ;
        RECT  1.210 2.160 1.320 2.320 ;
        RECT  1.050 2.160 1.210 3.160 ;
        RECT  0.770 1.450 1.160 1.730 ;
        RECT  0.880 2.880 1.050 3.160 ;
        RECT  0.770 0.440 0.890 0.720 ;
        RECT  0.770 1.910 0.890 2.190 ;
        RECT  0.610 0.440 0.770 2.190 ;
    END
END TLATX2TR

MACRO TLATX1TR
    CLASS CORE ;
    FOREIGN TLATX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 0.600 4.720 2.950 ;
        RECT  4.430 0.600 4.440 0.880 ;
        RECT  4.330 2.670 4.440 2.950 ;
        END
        ANTENNADIFFAREA 2.188 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.110 0.670 4.270 2.490 ;
        RECT  3.700 0.670 4.110 0.830 ;
        RECT  3.960 2.330 4.110 2.490 ;
        RECT  3.510 2.330 3.960 2.760 ;
        RECT  3.420 0.550 3.700 0.830 ;
        END
        ANTENNADIFFAREA 1.604 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.450 0.510 1.730 ;
        RECT  0.320 1.450 0.360 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 0.780 1.920 1.160 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.330 -0.280 4.800 0.280 ;
        RECT  4.050 -0.280 4.330 0.360 ;
        RECT  3.180 -0.280 4.050 0.280 ;
        RECT  2.900 -0.280 3.180 0.360 ;
        RECT  1.530 -0.280 2.900 0.280 ;
        RECT  1.230 -0.280 1.530 0.610 ;
        RECT  0.390 -0.280 1.230 0.280 ;
        RECT  0.110 -0.280 0.390 0.640 ;
        RECT  0.000 -0.280 0.110 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 3.320 4.800 3.880 ;
        RECT  3.850 2.920 4.130 3.880 ;
        RECT  3.270 3.320 3.850 3.880 ;
        RECT  2.990 3.200 3.270 3.880 ;
        RECT  1.660 3.260 2.990 3.880 ;
        RECT  1.380 2.960 1.660 3.880 ;
        RECT  0.390 3.320 1.380 3.880 ;
        RECT  0.110 3.260 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.740 1.130 3.950 2.170 ;
        RECT  3.670 1.010 3.740 2.170 ;
        RECT  3.460 1.010 3.670 1.290 ;
        RECT  3.060 1.890 3.670 2.170 ;
        RECT  2.660 1.450 3.500 1.730 ;
        RECT  2.900 1.890 3.060 2.950 ;
        RECT  2.780 2.610 2.900 2.950 ;
        RECT  2.500 0.440 2.660 2.090 ;
        RECT  2.330 2.540 2.620 3.070 ;
        RECT  2.200 0.440 2.500 0.720 ;
        RECT  2.420 1.930 2.500 2.090 ;
        RECT  2.140 1.930 2.420 2.210 ;
        RECT  1.250 2.540 2.330 2.770 ;
        RECT  1.250 1.350 2.200 1.510 ;
        RECT  1.090 0.770 1.250 2.770 ;
        RECT  0.870 2.930 1.150 3.160 ;
        RECT  1.070 0.770 1.090 0.930 ;
        RECT  0.700 2.550 1.090 2.770 ;
        RECT  0.910 0.550 1.070 0.930 ;
        RECT  0.830 1.410 0.930 1.690 ;
        RECT  0.620 0.550 0.910 0.830 ;
        RECT  0.540 2.930 0.870 3.090 ;
        RECT  0.670 1.070 0.830 2.280 ;
        RECT  0.550 1.070 0.670 1.290 ;
        RECT  0.540 1.960 0.670 2.280 ;
        RECT  0.520 1.960 0.540 3.090 ;
        RECT  0.380 2.120 0.520 3.090 ;
    END
END TLATX1TR

MACRO TIELOTR
    CLASS CORE ;
    FOREIGN TIELOTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.440 1.120 1.560 ;
        RECT  0.810 0.440 0.880 1.200 ;
        END
        ANTENNADIFFAREA 0.759 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 -0.280 1.200 0.280 ;
        RECT  0.290 -0.280 0.570 1.140 ;
        RECT  0.000 -0.280 0.290 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 3.320 1.200 3.880 ;
        RECT  0.130 1.970 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.730 1.910 1.040 2.190 ;
        RECT  0.720 1.730 0.730 2.190 ;
        RECT  0.570 1.510 0.720 2.190 ;
        RECT  0.490 1.510 0.570 1.790 ;
    END
END TIELOTR

MACRO TIEHITR
    CLASS CORE ;
    FOREIGN TIEHITR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.020 1.120 3.160 ;
        RECT  0.720 2.020 0.880 2.410 ;
        END
        ANTENNADIFFAREA 1.024 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 -0.280 1.200 0.280 ;
        RECT  0.200 -0.280 0.480 1.190 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 3.320 1.200 3.880 ;
        RECT  0.190 2.090 0.500 3.880 ;
        RECT  0.000 3.320 0.190 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 1.290 1.010 1.700 ;
        RECT  0.720 0.940 1.000 1.700 ;
        RECT  0.520 1.430 0.720 1.700 ;
    END
END TIEHITR

MACRO TBUFXLTR
    CLASS CORE ;
    FOREIGN TBUFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.590 3.120 2.750 ;
        RECT  2.860 0.590 2.880 0.870 ;
        END
        ANTENNAGATEAREA 1.144 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.470 0.610 1.630 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 2.440 2.320 2.820 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 -0.280 3.200 0.280 ;
        RECT  2.240 -0.280 2.520 0.800 ;
        RECT  0.780 -0.280 2.240 0.280 ;
        RECT  0.370 -0.280 0.780 0.390 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 3.320 3.200 3.880 ;
        RECT  2.400 3.260 2.760 3.880 ;
        RECT  1.960 3.320 2.400 3.880 ;
        RECT  1.680 3.260 1.960 3.880 ;
        RECT  0.420 3.320 1.680 3.880 ;
        RECT  0.140 2.780 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.500 0.960 2.660 1.300 ;
        RECT  2.500 2.100 2.660 2.420 ;
        RECT  1.950 0.960 2.500 1.120 ;
        RECT  1.710 2.100 2.500 2.260 ;
        RECT  1.790 0.440 1.950 1.120 ;
        RECT  1.270 0.440 1.790 0.720 ;
        RECT  1.630 1.310 1.710 3.090 ;
        RECT  1.550 1.030 1.630 3.090 ;
        RECT  1.470 1.030 1.550 1.470 ;
        RECT  0.700 2.930 1.550 3.090 ;
        RECT  1.270 2.080 1.390 2.240 ;
        RECT  1.110 0.440 1.270 2.240 ;
        RECT  0.930 2.400 1.000 2.680 ;
        RECT  0.930 0.630 0.950 0.910 ;
        RECT  0.770 0.630 0.930 2.680 ;
        RECT  0.650 2.060 0.770 2.220 ;
    END
END TBUFXLTR

MACRO TBUFX8TR
    CLASS CORE ;
    FOREIGN TBUFX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.540 0.440 4.820 3.160 ;
        RECT  3.900 1.040 4.540 1.770 ;
        RECT  3.680 0.550 3.900 3.160 ;
        RECT  3.580 0.550 3.680 1.080 ;
        RECT  3.580 2.120 3.680 3.160 ;
        END
        ANTENNAGATEAREA 7.648 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.640 0.720 1.960 ;
        RECT  0.080 1.630 0.450 1.960 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.450 2.610 1.670 ;
        RECT  2.290 1.450 2.450 2.660 ;
        RECT  2.040 1.640 2.290 1.960 ;
        RECT  1.530 2.500 2.290 2.660 ;
        RECT  1.370 2.000 1.530 2.660 ;
        RECT  1.200 2.000 1.370 2.350 ;
        END
        ANTENNAGATEAREA 0.4128 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.300 -0.280 5.600 0.280 ;
        RECT  5.020 -0.280 5.300 1.290 ;
        RECT  4.340 -0.280 5.020 0.280 ;
        RECT  4.060 -0.280 4.340 0.810 ;
        RECT  3.340 -0.280 4.060 0.280 ;
        RECT  2.370 -0.280 3.340 0.340 ;
        RECT  2.090 -0.280 2.370 0.400 ;
        RECT  0.240 -0.280 2.090 0.280 ;
        RECT  0.400 1.030 0.680 1.310 ;
        RECT  0.240 1.030 0.400 1.190 ;
        RECT  0.080 -0.280 0.240 1.190 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.300 3.320 5.600 3.880 ;
        RECT  5.020 1.950 5.300 3.880 ;
        RECT  4.340 3.320 5.020 3.880 ;
        RECT  4.060 1.950 4.340 3.880 ;
        RECT  3.370 3.320 4.060 3.880 ;
        RECT  3.090 2.120 3.370 3.880 ;
        RECT  0.890 3.260 3.090 3.880 ;
        RECT  0.610 2.930 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.420 1.240 3.520 1.520 ;
        RECT  2.930 1.680 3.430 1.960 ;
        RECT  3.260 0.810 3.420 1.520 ;
        RECT  2.890 0.810 3.260 0.970 ;
        RECT  2.770 1.130 2.930 3.100 ;
        RECT  2.610 0.690 2.890 0.970 ;
        RECT  2.070 1.130 2.770 1.290 ;
        RECT  2.610 2.060 2.770 3.100 ;
        RECT  1.630 0.690 2.610 0.850 ;
        RECT  1.210 2.820 2.610 3.100 ;
        RECT  1.850 2.120 2.130 2.340 ;
        RECT  1.790 1.030 2.070 1.310 ;
        RECT  1.690 1.470 1.850 2.340 ;
        RECT  1.630 1.470 1.690 1.630 ;
        RECT  1.470 0.690 1.630 1.630 ;
        RECT  1.310 0.850 1.470 1.130 ;
        RECT  1.150 1.360 1.310 1.640 ;
        RECT  1.050 2.610 1.210 3.100 ;
        RECT  1.040 1.320 1.150 1.640 ;
        RECT  0.410 2.610 1.050 2.770 ;
        RECT  1.000 1.320 1.040 2.400 ;
        RECT  0.880 0.590 1.000 2.400 ;
        RECT  0.840 0.590 0.880 1.480 ;
        RECT  0.130 2.120 0.880 2.400 ;
        RECT  0.680 0.590 0.840 0.750 ;
        RECT  0.400 0.470 0.680 0.750 ;
        RECT  0.130 2.610 0.410 2.890 ;
    END
END TBUFX8TR

MACRO TBUFX6TR
    CLASS CORE ;
    FOREIGN TBUFX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.450 4.280 3.110 ;
        RECT  3.360 1.030 4.000 1.770 ;
        RECT  3.140 0.450 3.360 3.070 ;
        RECT  3.100 0.450 3.140 1.180 ;
        RECT  3.060 1.810 3.140 3.070 ;
        RECT  3.040 2.180 3.060 3.070 ;
        END
        ANTENNAGATEAREA 7.097 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1824 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.490 2.240 1.770 ;
        RECT  1.760 1.490 1.920 2.730 ;
        RECT  1.670 1.490 1.760 2.020 ;
        RECT  1.160 2.570 1.760 2.730 ;
        RECT  0.890 2.440 1.160 2.730 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.800 -0.280 4.400 0.280 ;
        RECT  3.520 -0.280 3.800 0.860 ;
        RECT  2.800 -0.280 3.520 0.290 ;
        RECT  2.520 -0.280 2.800 0.410 ;
        RECT  0.240 -0.280 2.520 0.290 ;
        RECT  0.240 0.970 0.670 1.250 ;
        RECT  0.080 -0.280 0.240 1.250 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.800 3.320 4.400 3.880 ;
        RECT  3.520 2.040 3.800 3.880 ;
        RECT  2.840 3.320 3.520 3.880 ;
        RECT  2.560 2.450 2.840 3.880 ;
        RECT  0.620 3.270 2.560 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.940 1.300 2.980 1.580 ;
        RECT  2.780 0.630 2.940 1.580 ;
        RECT  2.560 1.740 2.900 2.020 ;
        RECT  2.280 0.630 2.780 0.790 ;
        RECT  2.400 1.170 2.560 2.290 ;
        RECT  1.940 1.170 2.400 1.330 ;
        RECT  2.360 2.130 2.400 2.290 ;
        RECT  2.080 2.130 2.360 3.110 ;
        RECT  2.000 0.510 2.280 0.790 ;
        RECT  0.380 2.890 2.080 3.110 ;
        RECT  1.480 0.500 2.000 0.790 ;
        RECT  1.660 0.990 1.940 1.330 ;
        RECT  1.480 2.190 1.600 2.410 ;
        RECT  1.320 0.500 1.480 2.410 ;
        RECT  1.200 0.970 1.320 1.250 ;
        RECT  1.040 1.540 1.160 1.820 ;
        RECT  0.990 1.310 1.040 2.280 ;
        RECT  0.880 0.530 0.990 2.280 ;
        RECT  0.830 0.530 0.880 1.480 ;
        RECT  0.720 2.120 0.880 2.280 ;
        RECT  0.680 0.530 0.830 0.690 ;
        RECT  0.100 2.120 0.720 2.450 ;
        RECT  0.400 0.470 0.680 0.690 ;
        RECT  0.100 2.830 0.380 3.110 ;
    END
END TBUFX6TR

MACRO TBUFX4TR
    CLASS CORE ;
    FOREIGN TBUFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.030 0.440 3.350 3.160 ;
        RECT  2.870 0.640 3.030 1.360 ;
        END
        ANTENNAGATEAREA 3.888 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.430 2.360 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.040 2.320 2.360 ;
        RECT  1.940 1.870 2.200 2.360 ;
        END
        ANTENNAGATEAREA 0.2016 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 -0.280 4.000 0.280 ;
        RECT  3.550 -0.280 3.830 1.270 ;
        RECT  2.580 -0.280 3.550 0.280 ;
        RECT  2.300 -0.280 2.580 0.800 ;
        RECT  0.460 -0.280 2.300 0.340 ;
        RECT  0.170 -0.280 0.460 0.800 ;
        RECT  0.000 -0.280 0.170 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 3.320 4.000 3.880 ;
        RECT  3.550 1.930 3.830 3.880 ;
        RECT  2.730 3.320 3.550 3.880 ;
        RECT  2.490 2.420 2.730 3.880 ;
        RECT  2.410 2.620 2.490 3.880 ;
        RECT  0.390 3.260 2.410 3.880 ;
        RECT  0.110 2.830 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.060 1.110 2.660 1.390 ;
        RECT  2.380 1.550 2.660 1.880 ;
        RECT  1.780 1.550 2.380 1.710 ;
        RECT  1.900 0.780 2.060 1.390 ;
        RECT  1.780 2.820 2.060 3.100 ;
        RECT  1.190 0.780 1.900 1.060 ;
        RECT  1.660 1.550 1.780 3.100 ;
        RECT  1.620 1.300 1.660 3.100 ;
        RECT  1.390 1.300 1.620 1.710 ;
        RECT  0.590 2.830 1.620 3.100 ;
        RECT  1.210 1.910 1.380 2.460 ;
        RECT  1.190 1.910 1.210 2.090 ;
        RECT  1.030 0.780 1.190 2.090 ;
        RECT  0.810 2.500 1.030 2.660 ;
        RECT  0.810 0.660 0.850 1.340 ;
        RECT  0.670 0.660 0.810 2.660 ;
        RECT  0.640 1.060 0.670 2.660 ;
    END
END TBUFX4TR

MACRO TBUFX3TR
    CLASS CORE ;
    FOREIGN TBUFX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.240 3.920 2.360 ;
        RECT  3.680 1.090 3.840 2.360 ;
        RECT  3.210 1.090 3.680 1.250 ;
        RECT  3.100 2.170 3.680 2.360 ;
        RECT  2.930 0.970 3.210 1.250 ;
        RECT  2.820 2.170 3.100 3.040 ;
        END
        ANTENNAGATEAREA 2.916 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.610 1.600 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.580 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 -0.280 4.000 0.280 ;
        RECT  3.410 -0.280 3.690 0.930 ;
        RECT  0.560 -0.280 3.410 0.280 ;
        RECT  0.250 -0.280 0.560 0.520 ;
        RECT  0.000 -0.280 0.250 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.580 3.320 4.000 3.880 ;
        RECT  3.300 2.760 3.580 3.880 ;
        RECT  2.620 3.320 3.300 3.880 ;
        RECT  2.400 2.170 2.620 3.880 ;
        RECT  0.450 3.320 2.400 3.880 ;
        RECT  0.170 2.570 0.450 3.880 ;
        RECT  0.000 3.320 0.170 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.680 1.410 3.410 1.580 ;
        RECT  2.240 1.810 2.910 1.970 ;
        RECT  2.520 0.450 2.680 1.580 ;
        RECT  1.290 0.450 2.520 0.610 ;
        RECT  2.080 1.150 2.240 2.800 ;
        RECT  1.610 1.150 2.080 1.310 ;
        RECT  1.360 2.640 2.080 2.800 ;
        RECT  1.450 1.030 1.610 1.310 ;
        RECT  1.340 1.470 1.500 2.300 ;
        RECT  1.290 1.470 1.340 1.630 ;
        RECT  1.130 0.450 1.290 1.630 ;
        RECT  0.970 2.400 1.200 2.560 ;
        RECT  0.810 0.630 0.970 2.560 ;
        RECT  0.780 0.630 0.810 1.310 ;
        RECT  0.750 1.940 0.810 2.220 ;
    END
END TBUFX3TR

MACRO TBUFX2TR
    CLASS CORE ;
    FOREIGN TBUFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.440 3.120 3.160 ;
        RECT  2.760 0.440 2.880 1.310 ;
        END
        ANTENNAGATEAREA 3.456 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.240 0.560 1.710 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 2.040 2.720 2.520 ;
        RECT  2.440 0.880 2.600 2.520 ;
        RECT  2.070 0.880 2.440 1.160 ;
        RECT  2.410 2.360 2.440 2.520 ;
        RECT  2.130 2.360 2.410 2.640 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.550 -0.280 3.200 0.280 ;
        RECT  2.270 -0.280 2.550 0.670 ;
        RECT  0.850 -0.280 2.270 0.280 ;
        RECT  0.450 -0.280 0.850 0.400 ;
        RECT  0.170 -0.280 0.450 0.740 ;
        RECT  0.000 -0.280 0.170 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 3.320 3.200 3.880 ;
        RECT  2.340 2.930 2.620 3.880 ;
        RECT  0.590 3.260 2.340 3.880 ;
        RECT  0.400 3.320 0.590 3.880 ;
        RECT  0.120 2.520 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 1.700 2.280 1.980 ;
        RECT  1.970 2.800 2.140 3.080 ;
        RECT  1.320 0.440 2.070 0.720 ;
        RECT  1.810 1.320 1.970 3.080 ;
        RECT  1.760 1.320 1.810 1.480 ;
        RECT  0.640 2.800 1.810 3.080 ;
        RECT  1.480 1.030 1.760 1.480 ;
        RECT  1.370 1.700 1.650 2.400 ;
        RECT  1.320 1.700 1.370 1.860 ;
        RECT  1.160 0.440 1.320 1.860 ;
        RECT  1.000 2.360 1.210 2.640 ;
        RECT  0.840 0.630 1.000 2.640 ;
        RECT  0.720 0.630 0.840 2.310 ;
        RECT  0.600 2.030 0.720 2.310 ;
    END
END TBUFX2TR

MACRO TBUFX20TR
    CLASS CORE ;
    FOREIGN TBUFX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  9.130 0.440 9.250 1.240 ;
        RECT  9.130 1.910 9.170 3.160 ;
        RECT  8.970 0.440 9.130 3.160 ;
        RECT  8.890 0.840 8.970 3.160 ;
        RECT  8.290 0.840 8.890 2.040 ;
        RECT  8.210 0.440 8.290 2.040 ;
        RECT  8.010 0.440 8.210 3.160 ;
        RECT  7.930 1.180 8.010 3.160 ;
        RECT  7.330 1.180 7.930 2.380 ;
        RECT  7.250 0.440 7.330 2.380 ;
        RECT  7.050 0.440 7.250 3.160 ;
        RECT  6.970 1.180 7.050 3.160 ;
        RECT  6.370 1.180 6.970 2.380 ;
        RECT  6.290 0.440 6.370 2.380 ;
        RECT  6.090 0.440 6.290 3.160 ;
        RECT  6.010 1.180 6.090 3.160 ;
        RECT  5.410 1.180 6.010 2.380 ;
        RECT  5.330 0.480 5.410 2.380 ;
        RECT  5.220 0.480 5.330 3.160 ;
        RECT  5.130 0.480 5.220 0.760 ;
        RECT  5.050 2.070 5.220 3.160 ;
        END
        ANTENNAGATEAREA 18.959 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.690 1.520 1.960 ;
        RECT  0.430 1.580 0.730 1.960 ;
        END
        ANTENNAGATEAREA 0.5088 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.360 4.570 1.640 ;
        RECT  3.640 1.240 4.000 1.640 ;
        RECT  3.410 1.340 3.640 1.640 ;
        END
        ANTENNAGATEAREA 0.9216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.770 -0.280 9.600 0.280 ;
        RECT  8.490 -0.280 8.770 0.680 ;
        RECT  7.810 -0.280 8.490 0.280 ;
        RECT  7.530 -0.280 7.810 1.020 ;
        RECT  6.850 -0.280 7.530 0.280 ;
        RECT  6.570 -0.280 6.850 1.010 ;
        RECT  5.890 -0.280 6.570 0.280 ;
        RECT  5.610 -0.280 5.890 1.010 ;
        RECT  4.850 -0.280 5.610 0.280 ;
        RECT  4.570 -0.280 4.850 0.760 ;
        RECT  3.890 -0.280 4.570 0.280 ;
        RECT  3.610 -0.280 3.890 0.750 ;
        RECT  1.930 -0.280 3.610 0.280 ;
        RECT  1.650 -0.280 1.930 0.740 ;
        RECT  0.890 -0.280 1.650 0.340 ;
        RECT  0.610 -0.280 0.890 0.800 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.690 3.320 9.600 3.880 ;
        RECT  8.410 2.410 8.690 3.880 ;
        RECT  7.730 3.320 8.410 3.880 ;
        RECT  7.450 2.560 7.730 3.880 ;
        RECT  6.770 3.320 7.450 3.880 ;
        RECT  6.490 2.560 6.770 3.880 ;
        RECT  5.810 3.320 6.490 3.880 ;
        RECT  5.530 2.570 5.810 3.880 ;
        RECT  4.850 3.320 5.530 3.880 ;
        RECT  4.570 2.120 4.850 3.880 ;
        RECT  3.890 3.320 4.570 3.880 ;
        RECT  3.610 2.120 3.890 3.880 ;
        RECT  1.930 3.320 3.610 3.880 ;
        RECT  1.650 3.160 1.930 3.880 ;
        RECT  0.890 3.260 1.650 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.780 0.920 5.060 1.470 ;
        RECT  4.890 1.630 5.060 1.910 ;
        RECT  4.730 1.630 4.890 1.960 ;
        RECT  4.370 0.920 4.780 1.080 ;
        RECT  4.370 1.800 4.730 1.960 ;
        RECT  4.090 0.670 4.370 1.080 ;
        RECT  4.090 1.800 4.370 3.160 ;
        RECT  3.410 0.920 4.090 1.080 ;
        RECT  3.410 1.800 4.090 1.960 ;
        RECT  3.130 0.710 3.410 1.080 ;
        RECT  3.250 1.800 3.410 3.160 ;
        RECT  3.090 1.240 3.250 3.160 ;
        RECT  2.490 0.710 3.130 0.870 ;
        RECT  2.930 1.240 3.090 1.400 ;
        RECT  2.450 3.000 3.090 3.160 ;
        RECT  2.650 1.030 2.930 1.400 ;
        RECT  2.650 1.970 2.930 2.840 ;
        RECT  2.490 1.970 2.650 2.130 ;
        RECT  2.330 0.710 2.490 2.130 ;
        RECT  2.170 2.610 2.450 3.160 ;
        RECT  2.170 0.710 2.330 1.060 ;
        RECT  1.410 0.900 2.170 1.060 ;
        RECT  2.050 1.850 2.170 2.130 ;
        RECT  1.410 2.610 2.170 2.770 ;
        RECT  1.890 1.340 2.050 2.130 ;
        RECT  1.270 1.340 1.890 1.500 ;
        RECT  1.130 0.780 1.410 1.060 ;
        RECT  1.130 2.490 1.410 2.770 ;
        RECT  1.000 1.220 1.270 1.500 ;
        RECT  0.370 1.220 1.000 1.380 ;
        RECT  0.270 0.890 0.370 1.380 ;
        RECT  0.270 2.120 0.370 2.880 ;
        RECT  0.110 0.890 0.270 2.880 ;
        RECT  0.090 0.890 0.110 1.230 ;
        RECT  0.090 2.120 0.110 2.880 ;
    END
END TBUFX20TR

MACRO TBUFX1TR
    CLASS CORE ;
    FOREIGN TBUFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.780 3.120 2.870 ;
        RECT  2.820 0.780 2.840 1.060 ;
        RECT  2.820 2.380 2.840 2.870 ;
        END
        ANTENNAGATEAREA 1.875 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.240 0.490 1.750 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 2.440 2.320 2.810 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.280 3.200 0.280 ;
        RECT  2.250 -0.280 2.530 0.830 ;
        RECT  0.770 -0.280 2.250 0.280 ;
        RECT  0.370 -0.280 0.770 0.370 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 3.320 3.200 3.880 ;
        RECT  1.820 3.260 2.620 3.880 ;
        RECT  0.370 3.320 1.820 3.880 ;
        RECT  0.090 2.700 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.400 1.160 2.680 1.440 ;
        RECT  1.750 1.940 2.680 2.220 ;
        RECT  2.090 1.160 2.400 1.320 ;
        RECT  1.930 0.440 2.090 1.320 ;
        RECT  1.330 0.440 1.930 0.720 ;
        RECT  1.750 1.030 1.770 1.310 ;
        RECT  1.590 1.030 1.750 3.100 ;
        RECT  1.490 1.030 1.590 1.310 ;
        RECT  1.370 2.940 1.590 3.100 ;
        RECT  1.330 2.120 1.410 2.280 ;
        RECT  0.650 2.940 1.370 3.160 ;
        RECT  1.170 0.440 1.330 2.280 ;
        RECT  1.130 2.120 1.170 2.280 ;
        RECT  0.870 2.480 1.080 2.640 ;
        RECT  0.930 0.630 1.010 0.910 ;
        RECT  0.870 0.630 0.930 1.310 ;
        RECT  0.730 0.630 0.870 2.640 ;
        RECT  0.710 1.030 0.730 2.640 ;
    END
END TBUFX1TR

MACRO TBUFX16TR
    CLASS CORE ;
    FOREIGN TBUFX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.890 0.440 7.170 3.100 ;
        RECT  6.810 0.440 6.890 2.360 ;
        RECT  6.210 1.240 6.810 2.360 ;
        RECT  6.130 1.240 6.210 3.100 ;
        RECT  5.930 0.440 6.130 3.100 ;
        RECT  5.850 0.440 5.930 2.360 ;
        RECT  5.250 1.240 5.850 2.360 ;
        RECT  5.170 1.240 5.250 3.100 ;
        RECT  4.970 0.440 5.170 3.100 ;
        RECT  4.890 0.440 4.970 2.830 ;
        RECT  4.590 0.770 4.890 2.830 ;
        RECT  4.210 0.770 4.590 1.440 ;
        RECT  4.290 2.110 4.590 2.830 ;
        RECT  4.010 2.110 4.290 3.130 ;
        RECT  4.040 0.550 4.210 1.440 ;
        RECT  3.930 0.550 4.040 1.190 ;
        END
        ANTENNAGATEAREA 15.248 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.450 2.360 ;
        END
        ANTENNAGATEAREA 0.4368 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.240 3.450 1.630 ;
        END
        ANTENNAGATEAREA 0.792 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.610 -0.280 7.600 0.280 ;
        RECT  6.330 -0.280 6.610 0.980 ;
        RECT  5.650 -0.280 6.330 0.280 ;
        RECT  5.370 -0.280 5.650 0.960 ;
        RECT  4.690 -0.280 5.370 0.280 ;
        RECT  4.410 -0.280 4.690 0.610 ;
        RECT  3.730 -0.280 4.410 0.280 ;
        RECT  3.450 -0.280 3.730 0.670 ;
        RECT  2.770 -0.280 3.450 0.280 ;
        RECT  2.490 -0.280 2.770 0.670 ;
        RECT  0.850 -0.280 2.490 0.340 ;
        RECT  0.570 -0.280 0.850 0.680 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.690 3.320 7.600 3.880 ;
        RECT  6.410 2.610 6.690 3.880 ;
        RECT  5.730 3.320 6.410 3.880 ;
        RECT  5.450 2.610 5.730 3.880 ;
        RECT  4.770 3.320 5.450 3.880 ;
        RECT  4.490 2.990 4.770 3.880 ;
        RECT  3.810 3.320 4.490 3.880 ;
        RECT  3.530 2.110 3.810 3.880 ;
        RECT  2.850 3.320 3.530 3.880 ;
        RECT  2.530 2.230 2.850 3.880 ;
        RECT  0.810 3.320 2.530 3.880 ;
        RECT  0.130 3.260 0.810 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.210 1.600 4.430 1.950 ;
        RECT  3.330 1.790 4.210 1.950 ;
        RECT  3.770 1.350 3.880 1.570 ;
        RECT  3.610 0.830 3.770 1.570 ;
        RECT  3.250 0.830 3.610 0.990 ;
        RECT  3.050 1.790 3.330 3.160 ;
        RECT  2.970 0.710 3.250 0.990 ;
        RECT  2.350 1.790 3.050 1.950 ;
        RECT  2.290 0.830 2.970 0.990 ;
        RECT  2.130 1.790 2.350 2.780 ;
        RECT  2.010 0.640 2.290 0.990 ;
        RECT  2.080 1.150 2.130 2.780 ;
        RECT  1.130 2.940 2.100 3.160 ;
        RECT  1.970 1.150 2.080 1.980 ;
        RECT  1.050 2.580 2.080 2.740 ;
        RECT  1.330 0.640 2.010 0.800 ;
        RECT  1.810 1.150 1.970 1.310 ;
        RECT  1.330 2.260 1.890 2.420 ;
        RECT  1.530 0.960 1.810 1.310 ;
        RECT  1.170 0.640 1.330 2.420 ;
        RECT  1.050 0.640 1.170 0.920 ;
        RECT  0.970 2.900 1.130 3.160 ;
        RECT  0.890 1.210 0.990 1.580 ;
        RECT  0.890 2.900 0.970 3.060 ;
        RECT  0.730 0.920 0.890 3.060 ;
        RECT  0.370 0.920 0.730 1.080 ;
        RECT  0.170 2.520 0.730 2.780 ;
        RECT  0.190 0.620 0.370 1.080 ;
        RECT  0.090 0.620 0.190 0.900 ;
    END
END TBUFX16TR

MACRO TBUFX12TR
    CLASS CORE ;
    FOREIGN TBUFX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.440 6.230 3.160 ;
        RECT  5.910 1.440 5.930 3.160 ;
        RECT  5.270 1.440 5.910 2.160 ;
        RECT  5.250 1.440 5.270 3.080 ;
        RECT  4.990 0.440 5.250 3.080 ;
        RECT  4.970 0.440 4.990 2.830 ;
        RECT  4.470 0.780 4.970 2.830 ;
        RECT  4.290 0.780 4.470 1.500 ;
        RECT  4.310 2.170 4.470 2.830 ;
        RECT  4.030 2.170 4.310 3.160 ;
        RECT  4.050 0.440 4.290 1.500 ;
        RECT  4.010 0.440 4.050 1.150 ;
        END
        ANTENNAGATEAREA 11.556 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.630 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.410 3.530 1.690 ;
        RECT  2.440 1.410 2.760 1.960 ;
        RECT  2.310 1.410 2.440 1.690 ;
        END
        ANTENNAGATEAREA 0.6312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.690 -0.280 6.800 0.280 ;
        RECT  6.410 -0.280 6.690 1.310 ;
        RECT  5.730 -0.280 6.410 0.280 ;
        RECT  5.450 -0.280 5.730 1.090 ;
        RECT  4.770 -0.280 5.450 0.280 ;
        RECT  4.490 -0.280 4.770 0.610 ;
        RECT  3.810 -0.280 4.490 0.280 ;
        RECT  3.530 -0.280 3.810 0.930 ;
        RECT  2.850 -0.280 3.530 0.340 ;
        RECT  2.570 -0.280 2.850 0.930 ;
        RECT  0.890 -0.280 2.570 0.340 ;
        RECT  0.610 -0.280 0.890 0.800 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.710 3.320 6.800 3.880 ;
        RECT  6.430 1.970 6.710 3.880 ;
        RECT  5.750 3.320 6.430 3.880 ;
        RECT  5.470 2.470 5.750 3.880 ;
        RECT  4.790 3.320 5.470 3.880 ;
        RECT  4.510 2.990 4.790 3.880 ;
        RECT  3.830 3.320 4.510 3.880 ;
        RECT  3.550 2.170 3.830 3.880 ;
        RECT  2.830 3.320 3.550 3.880 ;
        RECT  2.550 2.440 2.830 3.880 ;
        RECT  0.830 3.260 2.550 3.880 ;
        RECT  0.550 3.200 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.140 1.700 4.300 2.010 ;
        RECT  3.350 1.850 4.140 2.010 ;
        RECT  3.850 1.360 3.890 1.640 ;
        RECT  3.690 1.090 3.850 1.640 ;
        RECT  3.330 1.090 3.690 1.250 ;
        RECT  3.190 1.850 3.350 3.140 ;
        RECT  3.050 0.970 3.330 1.250 ;
        RECT  3.070 2.120 3.190 3.140 ;
        RECT  2.310 2.120 3.070 2.280 ;
        RECT  2.370 1.090 3.050 1.250 ;
        RECT  2.250 0.970 2.370 1.250 ;
        RECT  2.150 2.120 2.310 2.770 ;
        RECT  2.090 0.710 2.250 1.250 ;
        RECT  2.030 1.410 2.150 2.770 ;
        RECT  1.420 0.710 2.090 0.870 ;
        RECT  1.990 1.410 2.030 2.660 ;
        RECT  1.890 1.410 1.990 1.570 ;
        RECT  1.070 2.440 1.990 2.660 ;
        RECT  1.730 1.030 1.890 1.570 ;
        RECT  1.360 2.000 1.830 2.280 ;
        RECT  1.610 1.030 1.730 1.310 ;
        RECT  1.350 2.820 1.630 3.100 ;
        RECT  1.360 0.710 1.420 1.020 ;
        RECT  1.200 0.710 1.360 2.280 ;
        RECT  0.790 2.820 1.350 2.980 ;
        RECT  1.170 0.710 1.200 1.020 ;
        RECT  0.910 1.250 1.040 2.280 ;
        RECT  0.880 0.960 0.910 2.280 ;
        RECT  0.640 0.960 0.880 1.420 ;
        RECT  0.790 2.120 0.880 2.280 ;
        RECT  0.630 2.120 0.790 2.980 ;
        RECT  0.380 0.960 0.640 1.120 ;
        RECT  0.150 2.120 0.630 2.400 ;
        RECT  0.220 0.510 0.380 1.120 ;
        RECT  0.100 0.510 0.220 0.790 ;
    END
END TBUFX12TR

MACRO SMDFFHQX8TR
    CLASS CORE ;
    FOREIGN SMDFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.780 0.990 2.210 ;
        RECT  0.730 2.000 0.830 2.210 ;
        RECT  0.480 2.000 0.730 2.360 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.290 0.500 6.450 1.500 ;
        RECT  4.760 0.500 6.290 0.660 ;
        RECT  4.600 0.450 4.760 0.660 ;
        RECT  1.310 0.450 4.600 0.610 ;
        RECT  1.310 1.370 1.510 1.600 ;
        RECT  1.150 0.450 1.310 1.600 ;
        RECT  0.880 1.230 1.150 1.600 ;
        RECT  0.450 1.440 0.880 1.600 ;
        END
        ANTENNAGATEAREA 0.1824 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.690 1.540 6.850 1.820 ;
        RECT  5.920 1.660 6.690 1.820 ;
        RECT  5.690 1.640 5.920 1.960 ;
        RECT  5.680 1.270 5.690 1.960 ;
        RECT  5.530 1.270 5.680 1.800 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  20.670 0.440 20.950 3.160 ;
        RECT  20.660 0.440 20.670 1.780 ;
        RECT  19.970 1.010 20.660 1.780 ;
        RECT  19.680 0.440 19.970 3.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.640 3.120 1.960 ;
        RECT  2.880 1.480 3.040 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.720 1.410 8.750 1.690 ;
        RECT  8.590 1.240 8.720 1.690 ;
        RECT  8.480 1.240 8.590 1.560 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  10.720 1.400 10.830 1.560 ;
        RECT  10.480 1.240 10.720 1.560 ;
        RECT  10.150 1.400 10.480 1.560 ;
        END
        ANTENNAGATEAREA 0.3816 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  21.420 -0.280 21.600 0.280 ;
        RECT  21.180 -0.280 21.420 1.220 ;
        RECT  20.390 -0.280 21.180 0.280 ;
        RECT  20.230 -0.280 20.390 0.670 ;
        RECT  19.430 -0.280 20.230 0.280 ;
        RECT  19.270 -0.280 19.430 1.220 ;
        RECT  18.220 -0.280 19.270 0.280 ;
        RECT  17.900 -0.280 18.220 0.410 ;
        RECT  15.960 -0.280 17.900 0.280 ;
        RECT  15.680 -0.280 15.960 0.340 ;
        RECT  14.920 -0.280 15.680 0.280 ;
        RECT  14.640 -0.280 14.920 0.340 ;
        RECT  13.890 -0.280 14.640 0.280 ;
        RECT  13.610 -0.280 13.890 0.340 ;
        RECT  12.170 -0.280 13.610 0.280 ;
        RECT  11.890 -0.280 12.170 0.610 ;
        RECT  10.570 -0.280 11.890 0.280 ;
        RECT  10.410 -0.280 10.570 0.790 ;
        RECT  9.170 -0.280 10.410 0.280 ;
        RECT  8.890 -0.280 9.170 0.340 ;
        RECT  7.010 -0.280 8.890 0.280 ;
        RECT  6.700 -0.280 7.010 0.340 ;
        RECT  6.390 -0.280 6.700 0.280 ;
        RECT  6.110 -0.280 6.390 0.340 ;
        RECT  5.290 -0.280 6.110 0.280 ;
        RECT  5.010 -0.280 5.290 0.340 ;
        RECT  0.850 -0.280 5.010 0.280 ;
        RECT  0.570 -0.280 0.850 0.350 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  21.380 3.320 21.600 3.880 ;
        RECT  21.210 1.890 21.380 3.880 ;
        RECT  20.390 3.320 21.210 3.880 ;
        RECT  20.230 2.000 20.390 3.880 ;
        RECT  19.450 3.320 20.230 3.880 ;
        RECT  19.160 2.180 19.450 3.880 ;
        RECT  18.450 3.320 19.160 3.880 ;
        RECT  18.170 2.850 18.450 3.880 ;
        RECT  15.960 3.320 18.170 3.880 ;
        RECT  15.680 3.260 15.960 3.880 ;
        RECT  14.920 3.320 15.680 3.880 ;
        RECT  14.640 3.260 14.920 3.880 ;
        RECT  13.810 3.320 14.640 3.880 ;
        RECT  13.530 3.260 13.810 3.880 ;
        RECT  12.130 3.320 13.530 3.880 ;
        RECT  11.850 3.260 12.130 3.880 ;
        RECT  11.090 3.320 11.850 3.880 ;
        RECT  10.810 3.260 11.090 3.880 ;
        RECT  9.170 3.320 10.810 3.880 ;
        RECT  8.890 3.260 9.170 3.880 ;
        RECT  7.150 3.320 8.890 3.880 ;
        RECT  6.870 3.260 7.150 3.880 ;
        RECT  6.190 3.320 6.870 3.880 ;
        RECT  5.910 2.640 6.190 3.880 ;
        RECT  5.120 3.320 5.910 3.880 ;
        RECT  4.840 3.260 5.120 3.880 ;
        RECT  3.040 3.320 4.840 3.880 ;
        RECT  2.760 2.960 3.040 3.880 ;
        RECT  0.850 3.320 2.760 3.880 ;
        RECT  0.570 3.210 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  18.810 0.880 18.970 2.560 ;
        RECT  18.610 0.880 18.810 1.040 ;
        RECT  18.480 1.610 18.810 1.890 ;
        RECT  18.750 2.280 18.810 2.560 ;
        RECT  18.320 1.270 18.650 1.430 ;
        RECT  18.160 0.680 18.320 2.520 ;
        RECT  17.200 0.680 18.160 0.840 ;
        RECT  16.500 2.360 18.160 2.520 ;
        RECT  17.840 1.000 18.000 2.200 ;
        RECT  16.790 1.000 17.840 1.160 ;
        RECT  16.970 2.040 17.840 2.200 ;
        RECT  16.990 3.000 17.720 3.160 ;
        RECT  17.520 1.330 17.680 1.880 ;
        RECT  15.500 1.330 17.520 1.490 ;
        RECT  17.040 0.560 17.200 0.840 ;
        RECT  16.240 0.560 17.040 0.720 ;
        RECT  16.830 2.940 16.990 3.160 ;
        RECT  16.810 1.670 16.970 2.200 ;
        RECT  13.490 2.940 16.830 3.100 ;
        RECT  15.380 1.670 16.810 1.830 ;
        RECT  16.490 0.920 16.790 1.160 ;
        RECT  16.490 2.360 16.500 2.700 ;
        RECT  15.820 1.000 16.490 1.160 ;
        RECT  16.330 1.990 16.490 2.700 ;
        RECT  16.010 0.560 16.240 0.830 ;
        RECT  15.660 0.710 15.820 1.160 ;
        RECT  15.380 0.710 15.660 0.870 ;
        RECT  15.340 1.030 15.500 1.490 ;
        RECT  15.220 0.590 15.380 0.870 ;
        RECT  15.220 1.670 15.380 2.780 ;
        RECT  14.510 1.030 15.340 1.190 ;
        RECT  14.690 2.290 15.220 2.450 ;
        RECT  14.190 1.350 15.180 1.510 ;
        RECT  14.530 2.290 14.690 2.570 ;
        RECT  14.350 0.670 14.510 1.190 ;
        RECT  12.490 0.670 14.350 0.830 ;
        RECT  14.030 1.090 14.190 2.130 ;
        RECT  12.730 1.090 14.030 1.250 ;
        RECT  12.910 1.970 14.030 2.130 ;
        RECT  13.670 1.530 13.830 1.810 ;
        RECT  12.570 1.650 13.670 1.810 ;
        RECT  13.330 2.620 13.490 3.100 ;
        RECT  12.570 2.620 13.330 2.780 ;
        RECT  8.110 2.940 13.170 3.100 ;
        RECT  12.750 1.970 12.910 2.250 ;
        RECT  12.410 1.160 12.570 2.780 ;
        RECT  12.330 0.670 12.490 0.930 ;
        RECT  12.090 1.160 12.410 1.320 ;
        RECT  9.390 2.620 12.410 2.780 ;
        RECT  11.550 0.770 12.330 0.930 ;
        RECT  11.730 1.600 12.250 1.880 ;
        RECT  11.570 1.150 11.730 2.430 ;
        RECT  11.550 1.150 11.570 1.310 ;
        RECT  10.180 2.270 11.570 2.430 ;
        RECT  11.390 0.590 11.550 1.310 ;
        RECT  11.150 1.660 11.410 1.880 ;
        RECT  10.990 0.680 11.150 1.880 ;
        RECT  10.890 0.680 10.990 0.960 ;
        RECT  9.710 1.720 10.990 1.880 ;
        RECT  9.940 2.170 10.180 2.430 ;
        RECT  9.930 0.710 10.090 1.240 ;
        RECT  9.390 1.080 9.930 1.240 ;
        RECT  9.550 1.720 9.710 2.000 ;
        RECT  9.470 0.640 9.630 0.920 ;
        RECT  9.070 0.760 9.470 0.920 ;
        RECT  9.230 1.080 9.390 2.780 ;
        RECT  8.910 0.760 9.070 2.090 ;
        RECT  8.590 0.760 8.910 0.920 ;
        RECT  8.590 1.930 8.910 2.090 ;
        RECT  8.430 0.640 8.590 0.920 ;
        RECT  8.430 1.930 8.590 2.780 ;
        RECT  7.950 0.440 8.110 3.100 ;
        RECT  6.510 2.940 7.950 3.100 ;
        RECT  7.770 0.970 7.790 1.940 ;
        RECT  7.610 0.970 7.770 2.740 ;
        RECT  7.430 2.580 7.610 2.740 ;
        RECT  7.170 2.000 7.450 2.160 ;
        RECT  7.010 1.010 7.170 2.160 ;
        RECT  6.770 1.010 7.010 1.170 ;
        RECT  6.750 2.000 7.010 2.160 ;
        RECT  6.610 0.890 6.770 1.170 ;
        RECT  6.350 2.320 6.510 3.100 ;
        RECT  4.000 2.320 6.350 2.480 ;
        RECT  1.310 2.640 5.750 2.800 ;
        RECT  5.350 0.950 5.520 1.110 ;
        RECT  5.350 2.000 5.520 2.160 ;
        RECT  5.190 0.950 5.350 2.160 ;
        RECT  4.640 1.410 5.190 1.570 ;
        RECT  4.820 0.820 4.980 1.100 ;
        RECT  4.440 0.940 4.820 1.100 ;
        RECT  4.340 2.000 4.500 2.160 ;
        RECT  4.340 0.770 4.440 1.610 ;
        RECT  4.280 0.770 4.340 2.160 ;
        RECT  2.150 0.770 4.280 0.930 ;
        RECT  4.180 1.420 4.280 2.160 ;
        RECT  4.000 1.090 4.100 1.260 ;
        RECT  3.840 1.090 4.000 2.480 ;
        RECT  3.810 1.090 3.840 1.260 ;
        RECT  1.830 2.320 3.840 2.480 ;
        RECT  3.400 1.090 3.560 2.160 ;
        RECT  2.590 1.090 3.400 1.260 ;
        RECT  3.280 2.000 3.400 2.160 ;
        RECT  2.400 1.090 2.590 2.160 ;
        RECT  2.310 1.090 2.400 1.310 ;
        RECT  2.030 2.000 2.400 2.160 ;
        RECT  1.990 0.770 2.150 1.650 ;
        RECT  1.670 1.020 1.830 2.480 ;
        RECT  1.470 1.020 1.670 1.180 ;
        RECT  1.470 2.320 1.670 2.480 ;
        RECT  1.310 1.780 1.430 2.060 ;
        RECT  1.150 1.780 1.310 2.800 ;
        RECT  0.350 2.620 1.150 2.800 ;
        RECT  0.290 1.000 0.350 1.280 ;
        RECT  0.290 2.520 0.350 2.800 ;
        RECT  0.130 1.000 0.290 2.800 ;
    END
END SMDFFHQX8TR

MACRO SMDFFHQX4TR
    CLASS CORE ;
    FOREIGN SMDFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.780 0.990 2.210 ;
        RECT  0.730 2.000 0.830 2.210 ;
        RECT  0.480 2.000 0.730 2.360 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.290 0.500 6.450 1.500 ;
        RECT  4.760 0.500 6.290 0.660 ;
        RECT  4.600 0.450 4.760 0.660 ;
        RECT  1.310 0.450 4.600 0.610 ;
        RECT  1.310 1.370 1.510 1.600 ;
        RECT  1.150 0.450 1.310 1.600 ;
        RECT  0.880 1.230 1.150 1.600 ;
        RECT  0.450 1.440 0.880 1.600 ;
        END
        ANTENNAGATEAREA 0.1824 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.690 1.540 6.850 1.820 ;
        RECT  5.920 1.660 6.690 1.820 ;
        RECT  5.690 1.640 5.920 1.960 ;
        RECT  5.680 1.270 5.690 1.960 ;
        RECT  5.530 1.270 5.680 1.800 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.550 0.440 19.830 3.160 ;
        RECT  19.540 0.440 19.550 2.580 ;
        RECT  19.280 1.830 19.540 2.580 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.640 3.120 1.960 ;
        RECT  2.880 1.480 3.040 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.720 1.410 8.750 1.690 ;
        RECT  8.590 1.240 8.720 1.690 ;
        RECT  8.480 1.240 8.590 1.560 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  10.720 1.400 10.830 1.560 ;
        RECT  10.480 1.240 10.720 1.560 ;
        RECT  10.150 1.400 10.480 1.560 ;
        END
        ANTENNAGATEAREA 0.3816 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.250 -0.280 20.400 0.280 ;
        RECT  20.090 -0.280 20.250 1.220 ;
        RECT  19.290 -0.280 20.090 0.280 ;
        RECT  19.130 -0.280 19.290 1.220 ;
        RECT  18.310 -0.280 19.130 0.280 ;
        RECT  17.950 -0.280 18.310 0.410 ;
        RECT  15.960 -0.280 17.950 0.280 ;
        RECT  15.680 -0.280 15.960 0.340 ;
        RECT  14.920 -0.280 15.680 0.280 ;
        RECT  14.640 -0.280 14.920 0.340 ;
        RECT  13.890 -0.280 14.640 0.280 ;
        RECT  13.610 -0.280 13.890 0.340 ;
        RECT  12.170 -0.280 13.610 0.280 ;
        RECT  11.890 -0.280 12.170 0.610 ;
        RECT  10.570 -0.280 11.890 0.280 ;
        RECT  10.410 -0.280 10.570 0.790 ;
        RECT  9.170 -0.280 10.410 0.280 ;
        RECT  8.890 -0.280 9.170 0.340 ;
        RECT  7.010 -0.280 8.890 0.280 ;
        RECT  6.700 -0.280 7.010 0.340 ;
        RECT  6.390 -0.280 6.700 0.280 ;
        RECT  6.110 -0.280 6.390 0.340 ;
        RECT  5.290 -0.280 6.110 0.280 ;
        RECT  5.010 -0.280 5.290 0.340 ;
        RECT  0.850 -0.280 5.010 0.280 ;
        RECT  0.570 -0.280 0.850 0.350 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.250 3.320 20.400 3.880 ;
        RECT  20.090 1.820 20.250 3.880 ;
        RECT  19.310 3.320 20.090 3.880 ;
        RECT  19.030 3.260 19.310 3.880 ;
        RECT  18.450 3.320 19.030 3.880 ;
        RECT  18.170 2.790 18.450 3.880 ;
        RECT  15.960 3.320 18.170 3.880 ;
        RECT  15.680 3.260 15.960 3.880 ;
        RECT  14.920 3.320 15.680 3.880 ;
        RECT  14.640 3.260 14.920 3.880 ;
        RECT  13.810 3.320 14.640 3.880 ;
        RECT  13.530 3.260 13.810 3.880 ;
        RECT  12.130 3.320 13.530 3.880 ;
        RECT  11.850 3.260 12.130 3.880 ;
        RECT  11.090 3.320 11.850 3.880 ;
        RECT  10.810 3.260 11.090 3.880 ;
        RECT  9.170 3.320 10.810 3.880 ;
        RECT  8.890 3.260 9.170 3.880 ;
        RECT  7.150 3.320 8.890 3.880 ;
        RECT  6.870 3.260 7.150 3.880 ;
        RECT  6.190 3.320 6.870 3.880 ;
        RECT  5.910 2.640 6.190 3.880 ;
        RECT  5.120 3.320 5.910 3.880 ;
        RECT  4.840 3.260 5.120 3.880 ;
        RECT  3.040 3.320 4.840 3.880 ;
        RECT  2.760 2.960 3.040 3.880 ;
        RECT  0.850 3.320 2.760 3.880 ;
        RECT  0.570 3.210 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  18.810 0.880 18.970 2.560 ;
        RECT  18.610 0.880 18.810 1.040 ;
        RECT  18.480 1.610 18.810 1.890 ;
        RECT  18.790 2.280 18.810 2.560 ;
        RECT  18.320 1.270 18.650 1.430 ;
        RECT  18.160 0.680 18.320 2.520 ;
        RECT  17.200 0.680 18.160 0.840 ;
        RECT  16.500 2.360 18.160 2.520 ;
        RECT  17.840 1.000 18.000 2.200 ;
        RECT  16.790 1.000 17.840 1.160 ;
        RECT  16.970 2.040 17.840 2.200 ;
        RECT  16.280 3.000 17.720 3.160 ;
        RECT  17.520 1.330 17.680 1.880 ;
        RECT  15.500 1.330 17.520 1.490 ;
        RECT  17.040 0.560 17.200 0.840 ;
        RECT  16.240 0.560 17.040 0.720 ;
        RECT  16.810 1.670 16.970 2.200 ;
        RECT  15.380 1.670 16.810 1.830 ;
        RECT  16.490 0.920 16.790 1.160 ;
        RECT  16.490 2.360 16.500 2.700 ;
        RECT  15.820 1.000 16.490 1.160 ;
        RECT  16.330 1.990 16.490 2.700 ;
        RECT  16.120 2.940 16.280 3.160 ;
        RECT  16.010 0.560 16.240 0.830 ;
        RECT  13.490 2.940 16.120 3.100 ;
        RECT  15.660 0.710 15.820 1.160 ;
        RECT  15.380 0.710 15.660 0.870 ;
        RECT  15.340 1.030 15.500 1.490 ;
        RECT  15.220 0.590 15.380 0.870 ;
        RECT  15.220 1.670 15.380 2.780 ;
        RECT  14.510 1.030 15.340 1.190 ;
        RECT  14.690 2.290 15.220 2.450 ;
        RECT  14.190 1.350 15.180 1.510 ;
        RECT  14.530 2.290 14.690 2.570 ;
        RECT  14.350 0.670 14.510 1.190 ;
        RECT  12.490 0.670 14.350 0.830 ;
        RECT  14.030 1.090 14.190 2.130 ;
        RECT  12.730 1.090 14.030 1.250 ;
        RECT  12.910 1.970 14.030 2.130 ;
        RECT  13.670 1.530 13.830 1.810 ;
        RECT  12.570 1.650 13.670 1.810 ;
        RECT  13.330 2.620 13.490 3.100 ;
        RECT  12.570 2.620 13.330 2.780 ;
        RECT  8.110 2.940 13.170 3.100 ;
        RECT  12.750 1.970 12.910 2.250 ;
        RECT  12.410 1.160 12.570 2.780 ;
        RECT  12.330 0.670 12.490 0.930 ;
        RECT  12.090 1.160 12.410 1.320 ;
        RECT  9.390 2.620 12.410 2.780 ;
        RECT  11.550 0.770 12.330 0.930 ;
        RECT  11.730 1.600 12.250 1.880 ;
        RECT  11.570 1.150 11.730 2.430 ;
        RECT  11.550 1.150 11.570 1.310 ;
        RECT  10.180 2.270 11.570 2.430 ;
        RECT  11.390 0.590 11.550 1.310 ;
        RECT  11.150 1.660 11.410 1.880 ;
        RECT  10.990 0.680 11.150 1.880 ;
        RECT  10.890 0.680 10.990 0.960 ;
        RECT  9.710 1.720 10.990 1.880 ;
        RECT  9.940 2.170 10.180 2.430 ;
        RECT  9.930 0.710 10.090 1.240 ;
        RECT  9.390 1.080 9.930 1.240 ;
        RECT  9.550 1.720 9.710 2.000 ;
        RECT  9.470 0.640 9.630 0.920 ;
        RECT  9.070 0.760 9.470 0.920 ;
        RECT  9.230 1.080 9.390 2.780 ;
        RECT  8.910 0.760 9.070 2.090 ;
        RECT  8.590 0.760 8.910 0.920 ;
        RECT  8.590 1.930 8.910 2.090 ;
        RECT  8.430 0.640 8.590 0.920 ;
        RECT  8.430 1.930 8.590 2.780 ;
        RECT  7.950 0.440 8.110 3.100 ;
        RECT  6.510 2.940 7.950 3.100 ;
        RECT  7.770 0.970 7.790 1.940 ;
        RECT  7.610 0.970 7.770 2.740 ;
        RECT  7.430 2.580 7.610 2.740 ;
        RECT  7.170 2.000 7.450 2.160 ;
        RECT  7.010 1.010 7.170 2.160 ;
        RECT  6.770 1.010 7.010 1.170 ;
        RECT  6.750 2.000 7.010 2.160 ;
        RECT  6.610 0.890 6.770 1.170 ;
        RECT  6.350 2.320 6.510 3.100 ;
        RECT  3.980 2.320 6.350 2.480 ;
        RECT  1.310 2.640 5.750 2.800 ;
        RECT  5.340 0.950 5.520 1.110 ;
        RECT  5.340 2.000 5.520 2.160 ;
        RECT  5.180 0.950 5.340 2.160 ;
        RECT  4.640 1.410 5.180 1.570 ;
        RECT  4.810 0.820 4.970 1.100 ;
        RECT  4.440 0.940 4.810 1.100 ;
        RECT  4.310 2.000 4.500 2.160 ;
        RECT  4.310 0.770 4.440 1.610 ;
        RECT  4.280 0.770 4.310 2.160 ;
        RECT  2.150 0.770 4.280 0.930 ;
        RECT  4.150 1.420 4.280 2.160 ;
        RECT  3.980 1.090 4.100 1.260 ;
        RECT  3.820 1.090 3.980 2.480 ;
        RECT  3.810 1.090 3.820 1.260 ;
        RECT  1.830 2.320 3.820 2.480 ;
        RECT  3.400 1.090 3.560 2.160 ;
        RECT  2.590 1.090 3.400 1.260 ;
        RECT  3.280 2.000 3.400 2.160 ;
        RECT  2.400 1.090 2.590 2.160 ;
        RECT  2.310 1.090 2.400 1.310 ;
        RECT  2.030 2.000 2.400 2.160 ;
        RECT  1.990 0.770 2.150 1.650 ;
        RECT  1.670 1.020 1.830 2.480 ;
        RECT  1.470 1.020 1.670 1.180 ;
        RECT  1.470 2.320 1.670 2.480 ;
        RECT  1.310 1.780 1.430 2.060 ;
        RECT  1.150 1.780 1.310 2.800 ;
        RECT  0.350 2.620 1.150 2.800 ;
        RECT  0.290 1.000 0.350 1.280 ;
        RECT  0.290 2.520 0.350 2.800 ;
        RECT  0.130 1.000 0.290 2.800 ;
    END
END SMDFFHQX4TR

MACRO SMDFFHQX2TR
    CLASS CORE ;
    FOREIGN SMDFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.570 1.130 2.010 ;
        RECT  0.850 1.570 0.880 1.730 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.420 5.240 1.580 ;
        RECT  4.880 0.540 5.040 1.580 ;
        RECT  0.720 0.540 4.880 0.700 ;
        RECT  0.640 0.540 0.720 1.160 ;
        RECT  0.560 0.540 0.640 1.640 ;
        RECT  0.480 0.840 0.560 1.640 ;
        RECT  0.470 1.360 0.480 1.640 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 1.580 5.640 1.900 ;
        RECT  4.720 1.740 5.480 1.900 ;
        RECT  4.480 1.230 4.720 1.900 ;
        RECT  4.320 1.600 4.480 1.900 ;
        RECT  4.010 1.600 4.320 1.920 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.240 0.840 14.320 1.960 ;
        RECT  14.080 0.770 14.240 2.450 ;
        RECT  13.730 0.770 14.080 0.930 ;
        RECT  13.730 2.290 14.080 2.450 ;
        RECT  13.570 0.470 13.730 0.930 ;
        RECT  13.570 2.290 13.730 3.160 ;
        END
        ANTENNADIFFAREA 2.128 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.610 2.720 1.990 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.150 7.520 1.740 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.480 1.350 8.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2184 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.270 -0.280 14.400 0.280 ;
        RECT  13.990 -0.280 14.270 0.610 ;
        RECT  13.270 -0.280 13.990 0.280 ;
        RECT  12.990 -0.280 13.270 0.300 ;
        RECT  11.270 -0.280 12.990 0.280 ;
        RECT  10.990 -0.280 11.270 0.300 ;
        RECT  9.620 -0.280 10.990 0.280 ;
        RECT  8.320 -0.280 9.620 0.300 ;
        RECT  7.560 -0.280 8.320 0.280 ;
        RECT  7.400 -0.280 7.560 0.910 ;
        RECT  5.920 -0.280 7.400 0.280 ;
        RECT  5.640 -0.280 5.920 0.300 ;
        RECT  4.920 -0.280 5.640 0.280 ;
        RECT  4.640 -0.280 4.920 0.340 ;
        RECT  2.970 -0.280 4.640 0.280 ;
        RECT  2.690 -0.280 2.970 0.340 ;
        RECT  0.000 -0.280 2.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.250 3.320 14.400 3.880 ;
        RECT  14.090 2.880 14.250 3.880 ;
        RECT  13.250 3.320 14.090 3.880 ;
        RECT  13.090 2.520 13.250 3.880 ;
        RECT  11.270 3.320 13.090 3.880 ;
        RECT  10.990 3.240 11.270 3.880 ;
        RECT  9.700 3.320 10.990 3.880 ;
        RECT  9.420 3.260 9.700 3.880 ;
        RECT  7.700 3.320 9.420 3.880 ;
        RECT  7.420 3.260 7.700 3.880 ;
        RECT  5.180 3.320 7.420 3.880 ;
        RECT  4.900 2.860 5.180 3.880 ;
        RECT  3.940 3.320 4.900 3.880 ;
        RECT  3.660 3.260 3.940 3.880 ;
        RECT  2.890 3.320 3.660 3.880 ;
        RECT  2.610 2.950 2.890 3.880 ;
        RECT  0.890 3.320 2.610 3.880 ;
        RECT  0.610 2.550 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.750 1.090 13.910 2.130 ;
        RECT  13.550 1.090 13.750 1.250 ;
        RECT  13.070 1.970 13.750 2.130 ;
        RECT  13.390 1.440 13.590 1.600 ;
        RECT  13.230 0.510 13.390 1.600 ;
        RECT  12.370 0.510 13.230 0.670 ;
        RECT  12.910 1.400 13.070 2.130 ;
        RECT  12.530 1.060 12.690 3.160 ;
        RECT  11.590 3.000 12.530 3.160 ;
        RECT  12.210 0.510 12.370 1.760 ;
        RECT  12.050 1.600 12.210 2.800 ;
        RECT  11.890 0.510 12.050 1.440 ;
        RECT  9.480 0.510 11.890 0.670 ;
        RECT  11.570 0.830 11.730 2.760 ;
        RECT  11.430 2.920 11.590 3.160 ;
        RECT  10.820 2.280 11.570 2.440 ;
        RECT  10.940 2.920 11.430 3.080 ;
        RECT  11.020 1.180 11.410 1.460 ;
        RECT  10.860 0.960 11.020 2.100 ;
        RECT  10.780 2.600 10.940 3.080 ;
        RECT  10.440 0.960 10.860 1.120 ;
        RECT  10.400 1.940 10.860 2.100 ;
        RECT  10.080 2.600 10.780 2.760 ;
        RECT  10.080 1.620 10.700 1.780 ;
        RECT  10.280 0.830 10.440 1.120 ;
        RECT  10.240 1.940 10.400 2.220 ;
        RECT  9.980 2.940 10.260 3.160 ;
        RECT  9.920 1.240 10.080 2.760 ;
        RECT  6.800 2.940 9.980 3.100 ;
        RECT  9.800 1.240 9.920 1.400 ;
        RECT  7.990 2.600 9.920 2.760 ;
        RECT  9.640 1.120 9.800 1.400 ;
        RECT  9.480 1.560 9.760 1.840 ;
        RECT  9.320 0.510 9.480 2.360 ;
        RECT  8.820 0.510 9.320 0.870 ;
        RECT  8.480 2.200 9.320 2.360 ;
        RECT  9.040 1.260 9.160 1.420 ;
        RECT  8.880 1.030 9.040 1.420 ;
        RECT  8.560 1.030 8.880 1.190 ;
        RECT  8.400 0.560 8.560 1.190 ;
        RECT  8.320 2.200 8.480 2.440 ;
        RECT  8.310 1.030 8.400 1.190 ;
        RECT  8.150 1.030 8.310 1.990 ;
        RECT  7.990 0.690 8.100 0.850 ;
        RECT  7.820 0.690 7.990 2.760 ;
        RECT  7.120 2.050 7.140 2.330 ;
        RECT  6.960 0.450 7.120 2.330 ;
        RECT  6.840 0.450 6.960 0.610 ;
        RECT  6.640 0.770 6.800 3.160 ;
        RECT  6.460 0.770 6.640 0.930 ;
        RECT  6.440 2.360 6.640 2.520 ;
        RECT  5.500 3.000 6.640 3.160 ;
        RECT  6.320 1.090 6.480 1.980 ;
        RECT  6.300 0.570 6.460 0.930 ;
        RECT  6.200 1.090 6.320 1.250 ;
        RECT  6.280 1.820 6.320 1.980 ;
        RECT  6.120 1.820 6.280 2.840 ;
        RECT  5.960 1.440 6.160 1.600 ;
        RECT  5.940 2.680 6.120 2.840 ;
        RECT  5.800 1.050 5.960 2.220 ;
        RECT  5.200 1.050 5.800 1.210 ;
        RECT  5.620 2.060 5.800 2.220 ;
        RECT  5.340 2.410 5.500 3.160 ;
        RECT  3.530 2.410 5.340 2.570 ;
        RECT  3.210 2.730 4.740 2.890 ;
        RECT  3.850 2.090 4.500 2.250 ;
        RECT  3.850 1.030 3.990 1.310 ;
        RECT  3.690 1.030 3.850 2.250 ;
        RECT  3.310 1.520 3.690 1.680 ;
        RECT  3.370 2.310 3.530 2.570 ;
        RECT  3.150 1.990 3.490 2.150 ;
        RECT  3.310 0.890 3.470 1.360 ;
        RECT  1.670 2.310 3.370 2.470 ;
        RECT  3.150 1.200 3.310 1.360 ;
        RECT  3.050 2.630 3.210 2.890 ;
        RECT  2.990 1.200 3.150 2.150 ;
        RECT  1.470 2.630 3.050 2.790 ;
        RECT  2.270 1.200 2.990 1.360 ;
        RECT  1.950 0.860 2.410 1.020 ;
        RECT  2.110 1.200 2.270 1.480 ;
        RECT  2.000 1.640 2.160 2.150 ;
        RECT  1.950 1.640 2.000 1.800 ;
        RECT  1.790 0.860 1.950 1.800 ;
        RECT  1.630 2.180 1.670 2.470 ;
        RECT  1.470 0.880 1.630 2.470 ;
        RECT  1.310 2.630 1.470 2.910 ;
        RECT  1.210 2.630 1.310 2.790 ;
        RECT  1.050 2.170 1.210 2.790 ;
        RECT  0.310 2.170 1.050 2.330 ;
        RECT  0.150 1.030 0.310 2.330 ;
    END
END SMDFFHQX2TR

MACRO SMDFFHQX1TR
    CLASS CORE ;
    FOREIGN SMDFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.580 1.140 2.090 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 1.440 5.200 1.600 ;
        RECT  4.480 0.480 4.640 1.600 ;
        RECT  0.720 0.480 4.480 0.640 ;
        RECT  0.640 0.480 0.720 1.160 ;
        RECT  0.560 0.480 0.640 1.640 ;
        RECT  0.480 0.840 0.560 1.640 ;
        END
        ANTENNAGATEAREA 0.1512 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.420 1.600 5.580 1.920 ;
        RECT  4.320 1.760 5.420 1.920 ;
        RECT  4.010 1.240 4.320 1.920 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.230 1.240 14.320 2.560 ;
        RECT  14.070 0.720 14.230 2.560 ;
        RECT  13.790 0.720 14.070 0.880 ;
        RECT  13.730 2.400 14.070 2.560 ;
        RECT  13.570 0.470 13.790 0.880 ;
        RECT  13.570 2.400 13.730 3.000 ;
        END
        ANTENNADIFFAREA 1.031 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.240 7.520 1.620 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.480 1.240 8.720 1.710 ;
        RECT  8.000 1.550 8.480 1.710 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.310 -0.280 14.400 0.280 ;
        RECT  14.030 -0.280 14.310 0.340 ;
        RECT  5.880 -0.280 14.030 0.280 ;
        RECT  5.600 -0.280 5.880 0.730 ;
        RECT  4.880 -0.280 5.600 0.280 ;
        RECT  4.600 -0.280 4.880 0.320 ;
        RECT  2.980 -0.280 4.600 0.280 ;
        RECT  2.700 -0.280 2.980 0.320 ;
        RECT  0.000 -0.280 2.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.310 3.320 14.400 3.880 ;
        RECT  14.040 2.750 14.310 3.880 ;
        RECT  13.300 3.320 14.040 3.880 ;
        RECT  13.020 2.720 13.300 3.880 ;
        RECT  11.270 3.320 13.020 3.880 ;
        RECT  10.990 3.260 11.270 3.880 ;
        RECT  9.740 3.320 10.990 3.880 ;
        RECT  9.370 3.260 9.740 3.880 ;
        RECT  7.700 3.320 9.370 3.880 ;
        RECT  7.420 3.260 7.700 3.880 ;
        RECT  5.220 3.320 7.420 3.880 ;
        RECT  4.940 2.860 5.220 3.880 ;
        RECT  3.960 3.320 4.940 3.880 ;
        RECT  3.680 3.260 3.960 3.880 ;
        RECT  2.890 3.320 3.680 3.880 ;
        RECT  2.610 3.020 2.890 3.880 ;
        RECT  0.900 3.320 2.610 3.880 ;
        RECT  0.620 3.130 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.750 1.070 13.910 2.230 ;
        RECT  13.550 1.070 13.750 1.230 ;
        RECT  13.070 2.070 13.750 2.230 ;
        RECT  13.390 1.550 13.590 1.710 ;
        RECT  13.230 0.570 13.390 1.710 ;
        RECT  12.370 0.570 13.230 0.730 ;
        RECT  12.910 1.560 13.070 2.230 ;
        RECT  12.530 0.900 12.690 3.160 ;
        RECT  11.590 3.000 12.530 3.160 ;
        RECT  12.210 0.570 12.370 2.840 ;
        RECT  11.980 1.660 12.210 2.840 ;
        RECT  11.890 0.440 12.050 1.500 ;
        RECT  9.480 0.440 11.890 0.600 ;
        RECT  11.570 0.790 11.730 2.440 ;
        RECT  11.430 2.600 11.590 3.160 ;
        RECT  10.820 2.280 11.570 2.440 ;
        RECT  10.080 2.600 11.430 2.760 ;
        RECT  11.020 1.120 11.410 1.400 ;
        RECT  10.860 0.910 11.020 2.100 ;
        RECT  10.440 0.910 10.860 1.070 ;
        RECT  10.400 1.940 10.860 2.100 ;
        RECT  10.080 1.620 10.700 1.780 ;
        RECT  10.280 0.790 10.440 1.070 ;
        RECT  10.240 1.940 10.400 2.220 ;
        RECT  6.800 2.920 10.260 3.080 ;
        RECT  9.920 1.040 10.080 2.760 ;
        RECT  9.800 1.040 9.920 1.200 ;
        RECT  7.840 2.600 9.920 2.760 ;
        RECT  9.640 0.920 9.800 1.200 ;
        RECT  9.480 1.560 9.760 1.840 ;
        RECT  9.320 0.440 9.480 2.360 ;
        RECT  8.820 0.440 9.320 0.760 ;
        RECT  8.340 2.200 9.320 2.360 ;
        RECT  8.940 0.920 9.100 2.040 ;
        RECT  8.520 0.920 8.940 1.080 ;
        RECT  8.160 1.880 8.940 2.040 ;
        RECT  8.360 0.570 8.520 1.080 ;
        RECT  7.940 0.570 8.360 0.730 ;
        RECT  8.040 1.010 8.200 1.320 ;
        RECT  8.000 1.880 8.160 2.170 ;
        RECT  7.840 1.160 8.040 1.320 ;
        RECT  7.680 1.160 7.840 2.760 ;
        RECT  7.120 2.070 7.320 2.350 ;
        RECT  6.960 0.570 7.120 2.350 ;
        RECT  6.760 0.640 6.800 3.080 ;
        RECT  6.640 0.640 6.760 3.160 ;
        RECT  6.360 0.640 6.640 0.800 ;
        RECT  6.600 2.170 6.640 3.160 ;
        RECT  5.640 3.000 6.600 3.160 ;
        RECT  6.320 1.110 6.480 2.000 ;
        RECT  6.160 1.110 6.320 1.270 ;
        RECT  6.220 1.840 6.320 2.000 ;
        RECT  6.060 1.840 6.220 2.840 ;
        RECT  5.900 1.460 6.160 1.620 ;
        RECT  5.880 2.680 6.060 2.840 ;
        RECT  5.740 1.040 5.900 2.240 ;
        RECT  5.160 1.040 5.740 1.200 ;
        RECT  5.560 2.080 5.740 2.240 ;
        RECT  5.480 2.400 5.640 3.160 ;
        RECT  3.530 2.400 5.480 2.560 ;
        RECT  3.210 2.720 4.680 2.880 ;
        RECT  3.850 2.080 4.480 2.240 ;
        RECT  3.690 1.000 3.850 2.240 ;
        RECT  3.320 1.490 3.690 1.650 ;
        RECT  3.370 2.310 3.530 2.560 ;
        RECT  3.160 1.990 3.410 2.150 ;
        RECT  3.160 0.800 3.400 1.040 ;
        RECT  1.680 2.310 3.370 2.470 ;
        RECT  3.050 2.690 3.210 2.880 ;
        RECT  3.000 0.800 3.160 2.150 ;
        RECT  0.320 2.690 3.050 2.850 ;
        RECT  2.980 0.800 3.000 1.280 ;
        RECT  2.280 1.120 2.980 1.280 ;
        RECT  1.960 0.800 2.280 0.960 ;
        RECT  2.120 1.120 2.280 1.420 ;
        RECT  2.110 1.580 2.270 2.150 ;
        RECT  1.960 1.580 2.110 1.740 ;
        RECT  1.800 0.800 1.960 1.740 ;
        RECT  1.640 1.910 1.680 2.470 ;
        RECT  1.480 0.860 1.640 2.470 ;
        RECT  0.160 0.780 0.320 2.850 ;
    END
END SMDFFHQX1TR

MACRO SEDFFTRXLTR
    CLASS CORE ;
    FOREIGN SEDFFTRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.680 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.520 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.840 0.470 17.120 2.190 ;
        RECT  16.820 1.910 16.840 2.190 ;
        END
        ANTENNADIFFAREA 1.7335 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.000 0.470 16.020 1.420 ;
        RECT  15.800 0.470 16.000 2.190 ;
        RECT  15.780 1.240 15.800 2.190 ;
        RECT  15.680 1.240 15.780 1.780 ;
        END
        ANTENNADIFFAREA 1.651 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.640 6.320 2.010 ;
        RECT  5.640 1.640 6.040 1.810 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.390 4.300 1.670 ;
        RECT  3.960 1.390 4.080 1.550 ;
        RECT  3.920 1.240 3.960 1.550 ;
        RECT  3.680 1.240 3.920 1.560 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.100 1.240 8.360 1.590 ;
        RECT  8.040 1.240 8.100 1.710 ;
        RECT  7.820 1.430 8.040 1.710 ;
        END
        ANTENNAGATEAREA 0.0888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 -0.280 17.200 0.280 ;
        RECT  16.300 -0.280 16.580 0.800 ;
        RECT  15.160 -0.280 16.300 0.280 ;
        RECT  14.880 -0.280 15.160 0.520 ;
        RECT  13.980 -0.280 14.880 0.410 ;
        RECT  12.380 -0.280 13.980 0.280 ;
        RECT  12.160 -0.280 12.380 1.050 ;
        RECT  10.720 -0.280 12.160 0.280 ;
        RECT  10.440 -0.280 10.720 0.900 ;
        RECT  9.320 -0.280 10.440 0.280 ;
        RECT  9.320 1.210 9.440 1.430 ;
        RECT  9.160 -0.280 9.320 1.430 ;
        RECT  8.420 -0.280 9.160 0.280 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  6.120 -0.280 8.140 0.280 ;
        RECT  5.840 -0.280 6.120 0.350 ;
        RECT  5.040 -0.280 5.840 0.280 ;
        RECT  3.960 -0.280 5.040 0.400 ;
        RECT  1.790 -0.280 3.960 0.280 ;
        RECT  1.500 -0.280 1.790 0.400 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 3.320 17.200 3.880 ;
        RECT  16.300 3.200 16.580 3.880 ;
        RECT  15.180 3.320 16.300 3.880 ;
        RECT  13.950 3.060 15.180 3.880 ;
        RECT  12.260 3.320 13.950 3.880 ;
        RECT  11.980 3.260 12.260 3.880 ;
        RECT  10.840 3.320 11.980 3.880 ;
        RECT  10.560 3.260 10.840 3.880 ;
        RECT  8.300 3.320 10.560 3.880 ;
        RECT  8.020 2.990 8.300 3.880 ;
        RECT  6.120 3.320 8.020 3.880 ;
        RECT  5.840 2.990 6.120 3.880 ;
        RECT  4.240 3.320 5.840 3.880 ;
        RECT  3.960 2.990 4.240 3.880 ;
        RECT  1.700 3.320 3.960 3.880 ;
        RECT  1.420 3.200 1.700 3.880 ;
        RECT  0.000 3.320 1.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.380 1.580 16.660 2.510 ;
        RECT  15.480 2.350 16.380 2.510 ;
        RECT  15.480 0.470 15.620 0.750 ;
        RECT  15.480 1.910 15.540 2.190 ;
        RECT  15.320 0.470 15.480 2.510 ;
        RECT  14.880 1.580 15.160 1.960 ;
        RECT  14.680 1.800 14.880 1.960 ;
        RECT  14.520 0.860 14.680 2.590 ;
        RECT  14.400 0.860 14.520 1.140 ;
        RECT  14.350 1.800 14.520 2.590 ;
        RECT  14.240 1.320 14.360 1.540 ;
        RECT  13.900 1.800 14.350 1.960 ;
        RECT  13.900 2.430 14.350 2.590 ;
        RECT  14.080 0.630 14.240 1.540 ;
        RECT  13.380 0.630 14.080 0.790 ;
        RECT  13.740 1.580 13.900 1.960 ;
        RECT  13.790 2.430 13.900 2.830 ;
        RECT  13.740 2.430 13.790 3.160 ;
        RECT  13.630 2.670 13.740 3.160 ;
        RECT  12.540 3.000 13.630 3.160 ;
        RECT  13.420 0.980 13.580 2.510 ;
        RECT  13.320 0.980 13.420 1.200 ;
        RECT  13.150 2.350 13.420 2.510 ;
        RECT  13.140 0.520 13.380 0.790 ;
        RECT  13.140 1.910 13.260 2.190 ;
        RECT  12.880 2.350 13.150 2.840 ;
        RECT  13.100 0.520 13.140 2.190 ;
        RECT  12.980 0.630 13.100 2.190 ;
        RECT  10.400 2.350 12.880 2.630 ;
        RECT  12.660 0.770 12.820 2.190 ;
        RECT  12.580 0.770 12.660 1.050 ;
        RECT  12.500 1.910 12.660 2.190 ;
        RECT  12.400 2.940 12.540 3.160 ;
        RECT  12.380 1.280 12.500 1.560 ;
        RECT  9.320 2.940 12.400 3.100 ;
        RECT  12.220 1.210 12.380 1.560 ;
        RECT  12.000 1.210 12.220 1.370 ;
        RECT  11.840 0.450 12.000 1.370 ;
        RECT  11.680 1.910 11.860 2.190 ;
        RECT  11.300 0.450 11.840 0.610 ;
        RECT  11.460 0.770 11.680 2.190 ;
        RECT  11.140 0.450 11.300 2.190 ;
        RECT  10.900 0.450 11.140 0.730 ;
        RECT  11.080 1.910 11.140 2.190 ;
        RECT  10.600 1.910 11.080 2.070 ;
        RECT  10.760 1.220 10.980 1.750 ;
        RECT  10.080 1.220 10.760 1.380 ;
        RECT  10.320 1.540 10.600 2.070 ;
        RECT  10.240 2.350 10.400 2.780 ;
        RECT  9.640 2.600 10.240 2.780 ;
        RECT  9.960 1.220 10.080 2.430 ;
        RECT  9.800 0.740 9.960 2.430 ;
        RECT  9.760 0.740 9.800 0.900 ;
        RECT  9.480 0.620 9.760 0.900 ;
        RECT  9.480 1.870 9.640 2.780 ;
        RECT  8.680 1.870 9.480 2.070 ;
        RECT  9.160 2.350 9.320 3.100 ;
        RECT  7.400 2.350 9.160 2.510 ;
        RECT  8.720 2.670 9.000 2.950 ;
        RECT  7.720 2.670 8.720 2.830 ;
        RECT  8.520 0.920 8.680 2.190 ;
        RECT  7.880 0.920 8.520 1.080 ;
        RECT  7.780 2.030 8.520 2.190 ;
        RECT  7.600 0.920 7.880 1.270 ;
        RECT  7.560 1.910 7.780 2.190 ;
        RECT  7.560 2.670 7.720 3.150 ;
        RECT  7.400 0.480 7.560 0.760 ;
        RECT  6.440 2.990 7.560 3.150 ;
        RECT  7.240 0.480 7.400 2.830 ;
        RECT  7.080 2.670 7.240 2.830 ;
        RECT  6.920 0.520 7.080 2.510 ;
        RECT  6.800 0.520 6.920 0.800 ;
        RECT  6.880 2.350 6.920 2.510 ;
        RECT  6.600 2.350 6.880 2.730 ;
        RECT  6.640 1.570 6.760 2.190 ;
        RECT  6.480 0.440 6.640 2.190 ;
        RECT  5.160 2.350 6.600 2.510 ;
        RECT  6.300 0.440 6.480 0.790 ;
        RECT  6.280 2.670 6.440 3.150 ;
        RECT  5.680 1.210 6.320 1.440 ;
        RECT  5.200 0.510 6.300 0.790 ;
        RECT  3.600 2.670 6.280 2.830 ;
        RECT  5.480 0.960 5.680 1.440 ;
        RECT  5.480 1.970 5.680 2.190 ;
        RECT  5.400 0.960 5.480 2.190 ;
        RECT  5.320 1.270 5.400 2.190 ;
        RECT  5.160 1.550 5.320 1.830 ;
        RECT  5.000 1.990 5.160 2.510 ;
        RECT  5.000 0.950 5.120 1.230 ;
        RECT  4.880 0.630 5.000 2.510 ;
        RECT  4.840 0.630 4.880 2.150 ;
        RECT  3.680 0.630 4.840 0.790 ;
        RECT  4.460 0.950 4.680 2.190 ;
        RECT  4.360 0.950 4.460 1.230 ;
        RECT  3.560 0.440 3.680 0.790 ;
        RECT  3.520 1.910 3.680 2.190 ;
        RECT  3.440 2.670 3.600 2.970 ;
        RECT  3.400 0.440 3.560 0.930 ;
        RECT  3.240 1.090 3.520 2.190 ;
        RECT  2.760 2.810 3.440 2.970 ;
        RECT  3.080 0.770 3.400 0.930 ;
        RECT  3.080 2.370 3.280 2.650 ;
        RECT  2.760 0.450 3.160 0.610 ;
        RECT  2.920 0.770 3.080 2.650 ;
        RECT  2.600 0.450 2.760 2.970 ;
        RECT  2.480 1.910 2.600 2.190 ;
        RECT  2.280 0.520 2.440 0.800 ;
        RECT  2.160 2.380 2.440 2.660 ;
        RECT  0.700 2.820 2.320 3.040 ;
        RECT  2.120 0.520 2.280 2.220 ;
        RECT  1.080 2.380 2.160 2.540 ;
        RECT  1.920 2.060 2.120 2.220 ;
        RECT  0.920 1.030 1.080 2.540 ;
        RECT  0.700 0.570 0.990 0.850 ;
        RECT  0.860 1.910 0.920 2.540 ;
        RECT  0.540 0.570 0.700 3.040 ;
        RECT  0.420 2.580 0.540 3.040 ;
    END
END SEDFFTRXLTR

MACRO SEDFFTRX4TR
    CLASS CORE ;
    FOREIGN SEDFFTRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.680 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.520 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.680 1.040 17.940 1.760 ;
        RECT  17.400 0.590 17.680 2.990 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.560 1.440 16.740 2.160 ;
        RECT  16.320 0.560 16.560 2.570 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.640 6.320 2.010 ;
        RECT  5.640 1.640 6.040 1.810 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.390 4.300 1.670 ;
        RECT  3.960 1.390 4.080 1.550 ;
        RECT  3.920 1.240 3.960 1.550 ;
        RECT  3.680 1.240 3.920 1.560 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.100 1.240 8.360 1.590 ;
        RECT  8.040 1.240 8.100 1.710 ;
        RECT  7.820 1.430 8.040 1.710 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.180 -0.280 18.400 0.280 ;
        RECT  17.900 -0.280 18.180 0.860 ;
        RECT  17.120 -0.280 17.900 0.390 ;
        RECT  16.860 -0.280 17.120 1.310 ;
        RECT  16.120 -0.280 16.860 0.390 ;
        RECT  15.860 -0.280 16.120 1.310 ;
        RECT  15.150 -0.280 15.860 0.280 ;
        RECT  14.870 -0.280 15.150 0.420 ;
        RECT  13.860 -0.280 14.870 0.410 ;
        RECT  12.380 -0.280 13.860 0.280 ;
        RECT  12.160 -0.280 12.380 1.050 ;
        RECT  10.720 -0.280 12.160 0.280 ;
        RECT  10.440 -0.280 10.720 0.900 ;
        RECT  9.320 -0.280 10.440 0.280 ;
        RECT  9.320 1.210 9.440 1.430 ;
        RECT  9.160 -0.280 9.320 1.430 ;
        RECT  8.420 -0.280 9.160 0.280 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  6.120 -0.280 8.140 0.280 ;
        RECT  5.840 -0.280 6.120 0.350 ;
        RECT  4.240 -0.280 5.840 0.280 ;
        RECT  3.960 -0.280 4.240 0.400 ;
        RECT  1.790 -0.280 3.960 0.280 ;
        RECT  1.500 -0.280 1.790 0.890 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.180 3.320 18.400 3.880 ;
        RECT  18.140 3.200 18.180 3.880 ;
        RECT  17.880 1.930 18.140 3.880 ;
        RECT  15.140 3.200 17.880 3.880 ;
        RECT  14.890 2.210 15.140 3.880 ;
        RECT  14.010 3.200 14.890 3.880 ;
        RECT  12.260 3.320 14.010 3.880 ;
        RECT  11.980 3.260 12.260 3.880 ;
        RECT  10.840 3.320 11.980 3.880 ;
        RECT  10.560 3.260 10.840 3.880 ;
        RECT  8.300 3.320 10.560 3.880 ;
        RECT  8.020 2.990 8.300 3.880 ;
        RECT  6.120 3.320 8.020 3.880 ;
        RECT  5.840 2.990 6.120 3.880 ;
        RECT  4.240 3.320 5.840 3.880 ;
        RECT  3.960 2.990 4.240 3.880 ;
        RECT  1.700 3.320 3.960 3.880 ;
        RECT  1.420 3.200 1.700 3.880 ;
        RECT  0.000 3.320 1.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.940 1.580 17.220 2.890 ;
        RECT  15.640 2.730 16.940 2.890 ;
        RECT  15.460 0.910 15.640 2.890 ;
        RECT  15.320 0.910 15.460 1.310 ;
        RECT  15.350 2.200 15.460 2.890 ;
        RECT  15.100 1.580 15.280 2.000 ;
        RECT  14.680 1.840 15.100 2.000 ;
        RECT  14.520 0.860 14.680 2.770 ;
        RECT  14.400 0.860 14.520 1.140 ;
        RECT  14.350 1.840 14.520 2.770 ;
        RECT  14.240 1.460 14.360 1.680 ;
        RECT  13.900 1.840 14.350 2.000 ;
        RECT  13.850 2.610 14.350 2.770 ;
        RECT  14.080 0.630 14.240 1.680 ;
        RECT  13.380 0.630 14.080 0.790 ;
        RECT  13.740 1.580 13.900 2.000 ;
        RECT  13.690 2.610 13.850 3.100 ;
        RECT  9.320 2.940 13.690 3.100 ;
        RECT  13.530 1.080 13.600 1.300 ;
        RECT  13.370 1.080 13.530 2.780 ;
        RECT  13.140 0.520 13.380 0.790 ;
        RECT  13.320 1.080 13.370 1.300 ;
        RECT  10.240 2.530 13.370 2.780 ;
        RECT  13.140 2.030 13.200 2.310 ;
        RECT  13.100 0.520 13.140 2.310 ;
        RECT  12.980 0.630 13.100 2.310 ;
        RECT  12.660 0.770 12.820 2.310 ;
        RECT  12.580 0.770 12.660 1.050 ;
        RECT  12.500 2.030 12.660 2.310 ;
        RECT  12.380 1.390 12.500 1.630 ;
        RECT  12.220 1.210 12.380 1.630 ;
        RECT  12.000 1.210 12.220 1.370 ;
        RECT  11.840 0.450 12.000 1.370 ;
        RECT  11.680 2.030 11.860 2.310 ;
        RECT  11.300 0.450 11.840 0.610 ;
        RECT  11.460 0.770 11.680 2.310 ;
        RECT  11.140 0.450 11.300 2.190 ;
        RECT  10.900 0.450 11.140 0.680 ;
        RECT  11.080 1.910 11.140 2.190 ;
        RECT  10.600 1.910 11.080 2.070 ;
        RECT  10.760 1.220 10.980 1.750 ;
        RECT  10.080 1.220 10.760 1.380 ;
        RECT  10.320 1.540 10.600 2.070 ;
        RECT  9.640 2.600 10.240 2.780 ;
        RECT  9.960 1.220 10.080 2.430 ;
        RECT  9.800 0.740 9.960 2.430 ;
        RECT  9.760 0.740 9.800 0.900 ;
        RECT  9.480 0.620 9.760 0.900 ;
        RECT  9.480 1.870 9.640 2.780 ;
        RECT  8.680 1.870 9.480 2.070 ;
        RECT  9.160 2.350 9.320 3.100 ;
        RECT  7.400 2.350 9.160 2.510 ;
        RECT  8.720 2.670 9.000 2.950 ;
        RECT  7.720 2.670 8.720 2.830 ;
        RECT  8.520 0.920 8.680 2.190 ;
        RECT  7.880 0.920 8.520 1.080 ;
        RECT  7.780 2.030 8.520 2.190 ;
        RECT  7.600 0.920 7.880 1.270 ;
        RECT  7.560 1.910 7.780 2.190 ;
        RECT  7.560 2.670 7.720 3.150 ;
        RECT  6.440 2.990 7.560 3.150 ;
        RECT  7.400 0.480 7.520 0.710 ;
        RECT  7.240 0.480 7.400 2.830 ;
        RECT  7.040 2.670 7.240 2.830 ;
        RECT  6.920 0.460 7.080 2.510 ;
        RECT  6.820 0.460 6.920 0.740 ;
        RECT  6.840 2.350 6.920 2.510 ;
        RECT  6.600 2.350 6.840 2.730 ;
        RECT  6.640 1.570 6.760 2.190 ;
        RECT  6.480 0.440 6.640 2.190 ;
        RECT  5.160 2.350 6.600 2.510 ;
        RECT  6.300 0.440 6.480 0.790 ;
        RECT  6.280 2.670 6.440 3.150 ;
        RECT  5.680 1.210 6.320 1.440 ;
        RECT  5.160 0.510 6.300 0.790 ;
        RECT  3.600 2.670 6.280 2.830 ;
        RECT  5.480 0.960 5.680 1.440 ;
        RECT  5.480 1.970 5.680 2.190 ;
        RECT  5.400 0.960 5.480 2.190 ;
        RECT  5.320 1.270 5.400 2.190 ;
        RECT  5.160 1.550 5.320 1.830 ;
        RECT  5.000 1.990 5.160 2.510 ;
        RECT  5.000 0.950 5.120 1.230 ;
        RECT  4.880 0.630 5.000 2.510 ;
        RECT  4.840 0.630 4.880 2.150 ;
        RECT  3.680 0.630 4.840 0.790 ;
        RECT  4.460 0.950 4.680 2.190 ;
        RECT  4.360 0.950 4.460 1.230 ;
        RECT  3.560 0.440 3.680 0.790 ;
        RECT  3.520 1.910 3.680 2.190 ;
        RECT  3.440 2.670 3.600 2.970 ;
        RECT  3.400 0.440 3.560 0.930 ;
        RECT  3.240 1.090 3.520 2.190 ;
        RECT  2.760 2.810 3.440 2.970 ;
        RECT  3.080 0.770 3.400 0.930 ;
        RECT  3.080 2.370 3.280 2.650 ;
        RECT  2.760 0.450 3.160 0.610 ;
        RECT  2.920 0.770 3.080 2.650 ;
        RECT  2.600 0.450 2.760 2.970 ;
        RECT  2.480 1.910 2.600 2.190 ;
        RECT  2.280 0.520 2.440 0.800 ;
        RECT  2.160 2.380 2.440 2.660 ;
        RECT  0.700 2.820 2.320 3.040 ;
        RECT  2.120 0.520 2.280 2.220 ;
        RECT  1.080 2.380 2.160 2.540 ;
        RECT  1.920 2.060 2.120 2.220 ;
        RECT  0.920 1.030 1.080 2.540 ;
        RECT  0.700 0.570 1.010 0.850 ;
        RECT  0.860 1.910 0.920 2.540 ;
        RECT  0.540 0.570 0.700 3.040 ;
        RECT  0.420 2.580 0.540 3.040 ;
    END
END SEDFFTRX4TR

MACRO SEDFFTRX2TR
    CLASS CORE ;
    FOREIGN SEDFFTRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.680 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.520 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.840 0.540 17.120 3.070 ;
        RECT  16.820 1.910 16.840 3.070 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.780 1.030 16.000 2.190 ;
        RECT  15.680 1.030 15.780 1.780 ;
        END
        ANTENNADIFFAREA 3.466 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.640 6.320 2.010 ;
        RECT  5.640 1.640 6.040 1.810 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.390 4.300 1.670 ;
        RECT  3.960 1.390 4.080 1.550 ;
        RECT  3.920 1.240 3.960 1.550 ;
        RECT  3.680 1.240 3.920 1.560 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.100 1.240 8.360 1.590 ;
        RECT  8.040 1.240 8.100 1.710 ;
        RECT  7.820 1.430 8.040 1.710 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 -0.280 17.200 0.280 ;
        RECT  16.300 -0.280 16.580 1.220 ;
        RECT  15.160 -0.280 16.300 0.280 ;
        RECT  14.880 -0.280 15.160 0.520 ;
        RECT  13.860 -0.280 14.880 0.410 ;
        RECT  12.380 -0.280 13.860 0.280 ;
        RECT  12.160 -0.280 12.380 1.050 ;
        RECT  10.720 -0.280 12.160 0.280 ;
        RECT  10.440 -0.280 10.720 0.900 ;
        RECT  9.320 -0.280 10.440 0.280 ;
        RECT  9.320 1.210 9.440 1.430 ;
        RECT  9.160 -0.280 9.320 1.430 ;
        RECT  8.420 -0.280 9.160 0.280 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  6.120 -0.280 8.140 0.280 ;
        RECT  5.840 -0.280 6.120 0.350 ;
        RECT  4.240 -0.280 5.840 0.280 ;
        RECT  3.960 -0.280 4.240 0.400 ;
        RECT  1.790 -0.280 3.960 0.280 ;
        RECT  1.500 -0.280 1.790 0.910 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 3.320 17.200 3.880 ;
        RECT  16.300 2.850 16.580 3.880 ;
        RECT  15.180 3.320 16.300 3.880 ;
        RECT  14.900 2.850 15.180 3.880 ;
        RECT  14.010 3.200 14.900 3.880 ;
        RECT  12.260 3.320 14.010 3.880 ;
        RECT  11.980 3.260 12.260 3.880 ;
        RECT  10.840 3.320 11.980 3.880 ;
        RECT  10.560 3.260 10.840 3.880 ;
        RECT  8.300 3.320 10.560 3.880 ;
        RECT  8.020 2.990 8.300 3.880 ;
        RECT  6.060 3.320 8.020 3.880 ;
        RECT  5.780 2.990 6.060 3.880 ;
        RECT  4.240 3.320 5.780 3.880 ;
        RECT  3.960 2.990 4.240 3.880 ;
        RECT  1.700 3.320 3.960 3.880 ;
        RECT  1.420 3.200 1.700 3.880 ;
        RECT  0.000 3.320 1.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.380 1.580 16.660 2.510 ;
        RECT  15.480 2.350 16.380 2.510 ;
        RECT  15.480 0.470 15.620 0.750 ;
        RECT  15.480 1.910 15.540 2.190 ;
        RECT  15.320 0.470 15.480 2.510 ;
        RECT  14.880 1.580 15.160 2.000 ;
        RECT  14.680 1.840 14.880 2.000 ;
        RECT  14.520 0.860 14.680 2.770 ;
        RECT  14.400 0.860 14.520 1.140 ;
        RECT  14.350 1.840 14.520 2.770 ;
        RECT  14.240 1.460 14.360 1.680 ;
        RECT  13.900 1.840 14.350 2.000 ;
        RECT  13.850 2.610 14.350 2.770 ;
        RECT  14.080 0.630 14.240 1.680 ;
        RECT  13.380 0.630 14.080 0.790 ;
        RECT  13.740 1.580 13.900 2.000 ;
        RECT  13.690 2.610 13.850 3.100 ;
        RECT  9.320 2.940 13.690 3.100 ;
        RECT  13.530 1.080 13.600 1.300 ;
        RECT  13.370 1.080 13.530 2.780 ;
        RECT  13.140 0.520 13.380 0.790 ;
        RECT  13.320 1.080 13.370 1.300 ;
        RECT  10.240 2.530 13.370 2.780 ;
        RECT  13.140 2.030 13.200 2.310 ;
        RECT  13.100 0.520 13.140 2.310 ;
        RECT  12.980 0.630 13.100 2.310 ;
        RECT  12.660 0.770 12.820 2.310 ;
        RECT  12.580 0.770 12.660 1.050 ;
        RECT  12.500 2.030 12.660 2.310 ;
        RECT  12.380 1.390 12.500 1.630 ;
        RECT  12.220 1.210 12.380 1.630 ;
        RECT  12.000 1.210 12.220 1.370 ;
        RECT  11.840 0.450 12.000 1.370 ;
        RECT  11.680 2.030 11.860 2.310 ;
        RECT  11.300 0.450 11.840 0.610 ;
        RECT  11.460 0.770 11.680 2.310 ;
        RECT  11.140 0.450 11.300 2.190 ;
        RECT  10.900 0.450 11.140 0.730 ;
        RECT  11.080 1.910 11.140 2.190 ;
        RECT  10.600 1.910 11.080 2.070 ;
        RECT  10.760 1.220 10.980 1.750 ;
        RECT  10.080 1.220 10.760 1.380 ;
        RECT  10.320 1.540 10.600 2.070 ;
        RECT  9.640 2.600 10.240 2.780 ;
        RECT  9.960 1.220 10.080 2.430 ;
        RECT  9.800 0.740 9.960 2.430 ;
        RECT  9.760 0.740 9.800 0.900 ;
        RECT  9.480 0.620 9.760 0.900 ;
        RECT  9.480 1.870 9.640 2.780 ;
        RECT  8.680 1.870 9.480 2.070 ;
        RECT  9.160 2.350 9.320 3.100 ;
        RECT  7.400 2.350 9.160 2.510 ;
        RECT  8.720 2.670 9.000 2.950 ;
        RECT  7.720 2.670 8.720 2.830 ;
        RECT  8.520 0.920 8.680 2.190 ;
        RECT  7.880 0.920 8.520 1.080 ;
        RECT  7.780 2.030 8.520 2.190 ;
        RECT  7.600 0.920 7.880 1.270 ;
        RECT  7.560 1.910 7.780 2.190 ;
        RECT  7.560 2.670 7.720 3.150 ;
        RECT  7.400 0.480 7.560 0.700 ;
        RECT  6.440 2.990 7.560 3.150 ;
        RECT  7.240 0.480 7.400 2.830 ;
        RECT  7.080 2.670 7.240 2.830 ;
        RECT  6.920 0.520 7.080 2.510 ;
        RECT  6.800 0.520 6.920 0.800 ;
        RECT  6.880 2.350 6.920 2.510 ;
        RECT  6.600 2.350 6.880 2.730 ;
        RECT  6.640 1.570 6.760 2.190 ;
        RECT  6.480 0.440 6.640 2.190 ;
        RECT  5.160 2.350 6.600 2.510 ;
        RECT  6.300 0.440 6.480 0.790 ;
        RECT  6.280 2.670 6.440 3.150 ;
        RECT  5.680 1.210 6.320 1.440 ;
        RECT  5.160 0.510 6.300 0.790 ;
        RECT  3.600 2.670 6.280 2.830 ;
        RECT  5.480 0.960 5.680 1.440 ;
        RECT  5.480 1.970 5.680 2.190 ;
        RECT  5.400 0.960 5.480 2.190 ;
        RECT  5.320 1.270 5.400 2.190 ;
        RECT  5.160 1.550 5.320 1.830 ;
        RECT  5.000 1.990 5.160 2.510 ;
        RECT  5.000 0.950 5.120 1.230 ;
        RECT  4.880 0.630 5.000 2.510 ;
        RECT  4.840 0.630 4.880 2.150 ;
        RECT  3.680 0.630 4.840 0.790 ;
        RECT  4.460 0.950 4.680 2.190 ;
        RECT  4.360 0.950 4.460 1.230 ;
        RECT  3.560 0.440 3.680 0.790 ;
        RECT  3.520 1.910 3.680 2.190 ;
        RECT  3.440 2.670 3.600 2.970 ;
        RECT  3.400 0.440 3.560 0.930 ;
        RECT  3.240 1.090 3.520 2.190 ;
        RECT  2.760 2.810 3.440 2.970 ;
        RECT  3.080 0.770 3.400 0.930 ;
        RECT  3.080 2.370 3.280 2.650 ;
        RECT  2.760 0.450 3.160 0.610 ;
        RECT  2.920 0.770 3.080 2.650 ;
        RECT  2.600 0.450 2.760 2.970 ;
        RECT  2.480 1.910 2.600 2.190 ;
        RECT  2.280 0.520 2.440 0.800 ;
        RECT  2.160 2.380 2.440 2.660 ;
        RECT  0.700 2.820 2.320 3.040 ;
        RECT  2.120 0.520 2.280 2.220 ;
        RECT  1.080 2.380 2.160 2.540 ;
        RECT  1.920 2.060 2.120 2.220 ;
        RECT  0.920 1.030 1.080 2.540 ;
        RECT  0.700 0.570 1.060 0.850 ;
        RECT  0.860 1.910 0.920 2.540 ;
        RECT  0.540 0.570 0.700 3.040 ;
        RECT  0.420 2.580 0.540 3.040 ;
    END
END SEDFFTRX2TR

MACRO SEDFFTRX1TR
    CLASS CORE ;
    FOREIGN SEDFFTRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.680 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.520 1.520 2.090 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.840 0.840 17.120 2.190 ;
        RECT  16.820 1.910 16.840 2.190 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.780 1.030 16.000 2.190 ;
        RECT  15.680 1.030 15.780 1.780 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 1.640 6.320 2.010 ;
        RECT  5.640 1.640 5.950 1.810 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.390 4.300 1.670 ;
        RECT  3.680 1.240 4.160 1.670 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.040 1.240 8.360 1.710 ;
        RECT  7.820 1.430 8.040 1.710 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 -0.280 17.200 0.280 ;
        RECT  16.300 -0.280 16.580 0.800 ;
        RECT  15.160 -0.280 16.300 0.280 ;
        RECT  14.880 -0.280 15.160 0.520 ;
        RECT  13.960 -0.280 14.880 0.410 ;
        RECT  12.380 -0.280 13.960 0.280 ;
        RECT  12.160 -0.280 12.380 1.050 ;
        RECT  10.720 -0.280 12.160 0.280 ;
        RECT  10.440 -0.280 10.720 0.900 ;
        RECT  9.320 -0.280 10.440 0.280 ;
        RECT  9.320 1.210 9.440 1.430 ;
        RECT  9.160 -0.280 9.320 1.430 ;
        RECT  8.420 -0.280 9.160 0.280 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  6.120 -0.280 8.140 0.280 ;
        RECT  5.840 -0.280 6.120 0.350 ;
        RECT  4.240 -0.280 5.840 0.280 ;
        RECT  3.960 -0.280 4.240 0.400 ;
        RECT  1.790 -0.280 3.960 0.280 ;
        RECT  1.500 -0.280 1.790 0.850 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.580 3.320 17.200 3.880 ;
        RECT  16.300 3.200 16.580 3.880 ;
        RECT  15.180 3.320 16.300 3.880 ;
        RECT  13.950 3.060 15.180 3.880 ;
        RECT  12.260 3.320 13.950 3.880 ;
        RECT  11.980 3.260 12.260 3.880 ;
        RECT  10.840 3.320 11.980 3.880 ;
        RECT  10.560 3.260 10.840 3.880 ;
        RECT  8.300 3.320 10.560 3.880 ;
        RECT  8.020 2.990 8.300 3.880 ;
        RECT  6.120 3.320 8.020 3.880 ;
        RECT  5.840 2.990 6.120 3.880 ;
        RECT  4.240 3.320 5.840 3.880 ;
        RECT  3.960 2.990 4.240 3.880 ;
        RECT  1.700 3.320 3.960 3.880 ;
        RECT  1.420 3.200 1.700 3.880 ;
        RECT  0.000 3.320 1.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.380 1.580 16.660 2.510 ;
        RECT  15.480 2.350 16.380 2.510 ;
        RECT  15.480 0.470 15.620 0.750 ;
        RECT  15.480 1.910 15.540 2.190 ;
        RECT  15.320 0.470 15.480 2.510 ;
        RECT  14.880 1.580 15.160 1.960 ;
        RECT  14.680 1.800 14.880 1.960 ;
        RECT  14.520 0.860 14.680 2.590 ;
        RECT  14.400 0.860 14.520 1.140 ;
        RECT  14.350 1.800 14.520 2.590 ;
        RECT  14.240 1.360 14.360 1.640 ;
        RECT  13.900 1.800 14.350 1.960 ;
        RECT  13.900 2.430 14.350 2.590 ;
        RECT  14.080 0.630 14.240 1.640 ;
        RECT  13.380 0.630 14.080 0.790 ;
        RECT  13.740 1.580 13.900 1.960 ;
        RECT  13.790 2.430 13.900 2.830 ;
        RECT  13.740 2.430 13.790 3.160 ;
        RECT  13.630 2.670 13.740 3.160 ;
        RECT  12.540 3.000 13.630 3.160 ;
        RECT  13.470 0.980 13.580 2.510 ;
        RECT  13.420 0.980 13.470 2.840 ;
        RECT  13.320 0.980 13.420 1.200 ;
        RECT  13.190 2.350 13.420 2.840 ;
        RECT  13.140 0.520 13.380 0.790 ;
        RECT  13.140 1.910 13.260 2.190 ;
        RECT  10.400 2.350 13.190 2.630 ;
        RECT  13.100 0.520 13.140 2.190 ;
        RECT  12.980 0.630 13.100 2.190 ;
        RECT  12.660 0.770 12.820 2.190 ;
        RECT  12.580 0.770 12.660 1.050 ;
        RECT  12.500 1.910 12.660 2.190 ;
        RECT  12.400 2.940 12.540 3.160 ;
        RECT  12.380 1.280 12.500 1.560 ;
        RECT  9.320 2.940 12.400 3.100 ;
        RECT  12.220 1.210 12.380 1.560 ;
        RECT  12.000 1.210 12.220 1.370 ;
        RECT  11.840 0.450 12.000 1.370 ;
        RECT  11.680 1.910 11.860 2.190 ;
        RECT  11.300 0.450 11.840 0.610 ;
        RECT  11.460 0.770 11.680 2.190 ;
        RECT  11.140 0.450 11.300 2.190 ;
        RECT  10.900 0.450 11.140 0.730 ;
        RECT  11.080 1.910 11.140 2.190 ;
        RECT  10.600 1.910 11.080 2.070 ;
        RECT  10.760 1.220 10.980 1.750 ;
        RECT  10.080 1.220 10.760 1.380 ;
        RECT  10.320 1.540 10.600 2.070 ;
        RECT  10.240 2.350 10.400 2.780 ;
        RECT  9.640 2.600 10.240 2.780 ;
        RECT  9.960 1.220 10.080 2.430 ;
        RECT  9.800 0.740 9.960 2.430 ;
        RECT  9.760 0.740 9.800 0.900 ;
        RECT  9.480 0.620 9.760 0.900 ;
        RECT  9.480 1.870 9.640 2.780 ;
        RECT  8.680 1.870 9.480 2.070 ;
        RECT  9.160 2.350 9.320 3.100 ;
        RECT  7.400 2.350 9.160 2.510 ;
        RECT  8.720 2.670 9.000 2.950 ;
        RECT  7.720 2.670 8.720 2.830 ;
        RECT  8.520 0.920 8.680 2.190 ;
        RECT  7.880 0.920 8.520 1.080 ;
        RECT  7.780 2.030 8.520 2.190 ;
        RECT  7.600 0.920 7.880 1.270 ;
        RECT  7.560 1.910 7.780 2.190 ;
        RECT  7.560 2.670 7.720 3.150 ;
        RECT  7.400 0.480 7.560 0.760 ;
        RECT  6.440 2.990 7.560 3.150 ;
        RECT  7.240 0.480 7.400 2.830 ;
        RECT  7.080 2.670 7.240 2.830 ;
        RECT  6.920 0.520 7.080 2.510 ;
        RECT  6.800 0.520 6.920 0.800 ;
        RECT  6.880 2.350 6.920 2.510 ;
        RECT  6.600 2.350 6.880 2.730 ;
        RECT  6.640 1.570 6.760 2.190 ;
        RECT  6.480 0.440 6.640 2.190 ;
        RECT  5.160 2.350 6.600 2.510 ;
        RECT  6.300 0.440 6.480 0.790 ;
        RECT  6.280 2.670 6.440 3.150 ;
        RECT  5.680 1.210 6.320 1.440 ;
        RECT  5.160 0.510 6.300 0.790 ;
        RECT  3.600 2.670 6.280 2.830 ;
        RECT  5.480 0.960 5.680 1.440 ;
        RECT  5.480 1.970 5.680 2.190 ;
        RECT  5.400 0.960 5.480 2.190 ;
        RECT  5.320 1.270 5.400 2.190 ;
        RECT  5.160 1.550 5.320 1.830 ;
        RECT  5.000 1.990 5.160 2.510 ;
        RECT  5.000 0.950 5.120 1.230 ;
        RECT  4.880 0.630 5.000 2.510 ;
        RECT  4.840 0.630 4.880 2.150 ;
        RECT  3.680 0.630 4.840 0.790 ;
        RECT  4.460 0.950 4.680 2.190 ;
        RECT  4.360 0.950 4.460 1.230 ;
        RECT  3.560 0.440 3.680 0.790 ;
        RECT  3.520 1.910 3.680 2.190 ;
        RECT  3.440 2.670 3.600 2.970 ;
        RECT  3.400 0.440 3.560 0.930 ;
        RECT  3.240 1.090 3.520 2.190 ;
        RECT  2.760 2.810 3.440 2.970 ;
        RECT  3.080 0.770 3.400 0.930 ;
        RECT  3.080 2.370 3.280 2.650 ;
        RECT  2.760 0.450 3.160 0.610 ;
        RECT  2.920 0.770 3.080 2.650 ;
        RECT  2.600 0.450 2.760 2.970 ;
        RECT  2.480 1.910 2.600 2.190 ;
        RECT  2.280 0.520 2.440 0.800 ;
        RECT  2.160 2.380 2.440 2.660 ;
        RECT  0.700 2.820 2.320 3.040 ;
        RECT  2.120 0.520 2.280 2.220 ;
        RECT  1.080 2.380 2.160 2.540 ;
        RECT  1.920 2.060 2.120 2.220 ;
        RECT  0.920 1.030 1.080 2.540 ;
        RECT  0.700 0.570 1.030 0.850 ;
        RECT  0.860 1.910 0.920 2.540 ;
        RECT  0.540 0.570 0.700 3.040 ;
        RECT  0.420 2.580 0.540 3.040 ;
    END
END SEDFFTRX1TR

MACRO SEDFFHQX8TR
    CLASS CORE ;
    FOREIGN SEDFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.820 1.040 2.360 ;
        RECT  0.480 2.040 0.880 2.360 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.140 0.500 6.300 1.550 ;
        RECT  4.580 0.500 6.140 0.660 ;
        RECT  4.420 0.440 4.580 0.660 ;
        RECT  1.360 0.440 4.420 0.600 ;
        RECT  1.360 1.380 1.480 1.660 ;
        RECT  1.320 0.440 1.360 1.660 ;
        RECT  1.200 0.440 1.320 1.600 ;
        RECT  0.880 1.240 1.200 1.600 ;
        RECT  0.500 1.440 0.880 1.600 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.940 0.440 20.220 3.070 ;
        RECT  19.300 1.840 19.940 2.560 ;
        RECT  19.260 1.840 19.300 3.160 ;
        RECT  18.920 0.440 19.260 3.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.540 1.570 6.700 1.870 ;
        RECT  5.920 1.710 6.540 1.870 ;
        RECT  5.680 1.640 5.920 1.960 ;
        RECT  5.540 1.640 5.680 1.800 ;
        RECT  5.380 1.270 5.540 1.800 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.480 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  9.480 1.240 10.160 1.560 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.700 -0.280 20.800 0.280 ;
        RECT  20.420 -0.280 20.700 1.250 ;
        RECT  19.700 -0.280 20.420 0.280 ;
        RECT  19.420 -0.280 19.700 1.220 ;
        RECT  18.680 -0.280 19.420 0.280 ;
        RECT  18.520 -0.280 18.680 1.080 ;
        RECT  17.620 -0.280 18.520 0.280 ;
        RECT  17.340 -0.280 17.620 0.340 ;
        RECT  10.740 -0.280 17.340 0.280 ;
        RECT  10.460 -0.280 10.740 0.340 ;
        RECT  9.980 -0.280 10.460 0.280 ;
        RECT  9.700 -0.280 9.980 0.340 ;
        RECT  8.820 -0.280 9.700 0.280 ;
        RECT  8.540 -0.280 8.820 0.340 ;
        RECT  7.160 -0.280 8.540 0.280 ;
        RECT  6.880 -0.280 7.160 0.340 ;
        RECT  6.240 -0.280 6.880 0.280 ;
        RECT  5.960 -0.280 6.240 0.340 ;
        RECT  0.900 -0.280 5.960 0.280 ;
        RECT  0.620 -0.280 0.900 0.340 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.700 3.320 20.800 3.880 ;
        RECT  20.420 1.910 20.700 3.880 ;
        RECT  19.740 3.320 20.420 3.880 ;
        RECT  19.460 2.880 19.740 3.880 ;
        RECT  18.700 3.320 19.460 3.880 ;
        RECT  18.420 3.260 18.700 3.880 ;
        RECT  17.880 3.320 18.420 3.880 ;
        RECT  17.600 2.800 17.880 3.880 ;
        RECT  15.440 3.320 17.600 3.880 ;
        RECT  15.160 3.260 15.440 3.880 ;
        RECT  14.400 3.320 15.160 3.880 ;
        RECT  14.120 3.260 14.400 3.880 ;
        RECT  13.260 3.320 14.120 3.880 ;
        RECT  12.980 3.260 13.260 3.880 ;
        RECT  11.580 3.320 12.980 3.880 ;
        RECT  11.300 3.260 11.580 3.880 ;
        RECT  10.540 3.320 11.300 3.880 ;
        RECT  10.260 3.260 10.540 3.880 ;
        RECT  8.700 3.320 10.260 3.880 ;
        RECT  8.420 3.260 8.700 3.880 ;
        RECT  6.960 3.320 8.420 3.880 ;
        RECT  6.680 3.260 6.960 3.880 ;
        RECT  6.040 3.320 6.680 3.880 ;
        RECT  5.760 2.800 6.040 3.880 ;
        RECT  4.960 3.320 5.760 3.880 ;
        RECT  4.680 3.260 4.960 3.880 ;
        RECT  2.520 3.320 4.680 3.880 ;
        RECT  2.240 3.020 2.520 3.880 ;
        RECT  0.900 3.320 2.240 3.880 ;
        RECT  0.620 3.260 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  18.200 0.870 18.360 2.560 ;
        RECT  18.160 0.870 18.200 1.030 ;
        RECT  18.180 1.610 18.200 2.560 ;
        RECT  18.000 1.610 18.180 1.890 ;
        RECT  18.000 0.500 18.160 1.030 ;
        RECT  17.840 1.270 18.040 1.430 ;
        RECT  17.140 0.500 18.000 0.660 ;
        RECT  17.680 0.820 17.840 2.490 ;
        RECT  16.820 0.820 17.680 0.980 ;
        RECT  15.920 2.330 17.680 2.490 ;
        RECT  17.360 1.140 17.520 2.170 ;
        RECT  16.300 1.140 17.360 1.300 ;
        RECT  16.460 2.010 17.360 2.170 ;
        RECT  17.040 1.460 17.200 1.850 ;
        RECT  15.760 3.000 17.150 3.160 ;
        RECT  16.980 0.440 17.140 0.660 ;
        RECT  15.020 1.460 17.040 1.620 ;
        RECT  11.060 0.440 16.980 0.600 ;
        RECT  16.660 0.760 16.820 0.980 ;
        RECT  15.500 0.760 16.660 0.920 ;
        RECT  16.170 1.820 16.460 2.170 ;
        RECT  16.020 1.080 16.300 1.300 ;
        RECT  14.860 1.820 16.170 1.980 ;
        RECT  15.340 1.140 16.020 1.300 ;
        RECT  15.760 2.210 15.920 2.490 ;
        RECT  15.600 2.940 15.760 3.160 ;
        RECT  12.940 2.940 15.600 3.100 ;
        RECT  15.180 0.760 15.340 1.300 ;
        RECT  14.630 0.760 15.180 0.920 ;
        RECT  14.860 1.120 15.020 1.620 ;
        RECT  13.960 1.120 14.860 1.280 ;
        RECT  14.700 1.820 14.860 2.780 ;
        RECT  13.640 1.440 14.700 1.600 ;
        RECT  14.170 2.240 14.700 2.400 ;
        RECT  14.010 2.240 14.170 2.580 ;
        RECT  13.800 0.760 13.960 1.280 ;
        RECT  11.380 0.760 13.800 0.920 ;
        RECT  13.480 1.080 13.640 2.180 ;
        RECT  13.260 1.080 13.480 1.300 ;
        RECT  12.360 2.020 13.480 2.180 ;
        RECT  13.120 1.540 13.280 1.820 ;
        RECT  12.180 1.080 13.260 1.240 ;
        RECT  12.020 1.660 13.120 1.820 ;
        RECT  12.780 2.580 12.940 3.100 ;
        RECT  12.020 2.580 12.780 2.740 ;
        RECT  12.020 2.940 12.620 3.100 ;
        RECT  12.200 2.020 12.360 2.330 ;
        RECT  11.860 1.240 12.020 2.740 ;
        RECT  11.850 2.920 12.020 3.100 ;
        RECT  11.540 1.240 11.860 1.400 ;
        RECT  8.260 2.580 11.860 2.740 ;
        RECT  7.940 2.920 11.850 3.080 ;
        RECT  11.380 1.580 11.700 1.860 ;
        RECT  11.220 0.760 11.380 2.400 ;
        RECT  10.780 1.090 11.220 1.250 ;
        RECT  10.560 2.240 11.220 2.400 ;
        RECT  10.900 0.440 11.060 0.660 ;
        RECT  9.620 0.500 10.900 0.660 ;
        RECT  10.500 1.860 10.860 2.020 ;
        RECT  10.370 2.180 10.560 2.400 ;
        RECT  10.340 0.840 10.500 2.020 ;
        RECT  9.320 2.180 10.370 2.340 ;
        RECT  10.220 0.840 10.340 1.000 ;
        RECT  9.160 1.860 10.340 2.020 ;
        RECT  9.460 0.500 9.620 0.980 ;
        RECT  8.810 0.820 9.460 0.980 ;
        RECT  8.260 0.500 9.300 0.660 ;
        RECT  9.000 1.740 9.160 2.020 ;
        RECT  8.640 0.820 8.810 1.120 ;
        RECT  8.420 0.960 8.640 1.120 ;
        RECT  8.100 0.500 8.260 2.740 ;
        RECT  7.780 0.620 7.940 3.080 ;
        RECT  7.660 0.620 7.780 0.780 ;
        RECT  7.760 2.230 7.780 3.080 ;
        RECT  6.360 2.920 7.760 3.080 ;
        RECT  7.600 1.020 7.620 1.940 ;
        RECT  7.460 1.020 7.600 2.740 ;
        RECT  7.440 1.660 7.460 2.740 ;
        RECT  7.240 2.580 7.440 2.740 ;
        RECT  7.020 2.030 7.280 2.190 ;
        RECT  6.860 1.030 7.020 2.190 ;
        RECT  6.620 1.030 6.860 1.190 ;
        RECT  6.600 2.030 6.860 2.190 ;
        RECT  6.460 0.910 6.620 1.190 ;
        RECT  6.200 2.380 6.360 3.080 ;
        RECT  4.280 2.380 6.200 2.540 ;
        RECT  5.380 2.820 5.540 3.100 ;
        RECT  2.840 2.940 5.380 3.100 ;
        RECT  5.220 0.950 5.360 1.110 ;
        RECT  5.220 2.000 5.360 2.160 ;
        RECT  5.060 0.950 5.220 2.160 ;
        RECT  4.460 1.260 5.060 1.420 ;
        RECT  4.680 0.820 4.840 1.100 ;
        RECT  4.260 0.940 4.680 1.100 ;
        RECT  4.260 2.000 4.380 2.160 ;
        RECT  4.120 2.380 4.280 2.780 ;
        RECT  4.100 0.760 4.260 2.160 ;
        RECT  3.820 2.620 4.120 2.780 ;
        RECT  2.120 0.760 4.100 0.920 ;
        RECT  3.980 1.410 4.100 1.570 ;
        RECT  3.820 1.080 3.940 1.240 ;
        RECT  3.660 1.080 3.820 2.780 ;
        RECT  3.160 2.620 3.660 2.780 ;
        RECT  3.320 1.080 3.480 2.280 ;
        RECT  2.440 1.080 3.320 1.240 ;
        RECT  3.000 2.380 3.160 2.780 ;
        RECT  1.800 2.380 3.000 2.540 ;
        RECT  2.680 2.700 2.840 3.100 ;
        RECT  1.360 2.700 2.680 2.860 ;
        RECT  2.280 1.080 2.440 2.220 ;
        RECT  2.080 2.060 2.280 2.220 ;
        RECT  1.960 0.760 2.120 1.640 ;
        RECT  1.640 1.060 1.800 2.540 ;
        RECT  1.520 1.060 1.640 1.220 ;
        RECT  1.520 2.260 1.640 2.540 ;
        RECT  1.360 1.820 1.480 2.100 ;
        RECT  1.200 1.820 1.360 2.860 ;
        RECT  0.320 2.700 1.200 2.860 ;
        RECT  0.320 1.000 0.400 1.280 ;
        RECT  0.160 1.000 0.320 2.860 ;
    END
END SEDFFHQX8TR

MACRO SEDFFHQX4TR
    CLASS CORE ;
    FOREIGN SEDFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.820 1.200 2.200 ;
        RECT  1.040 1.820 1.120 2.360 ;
        RECT  0.880 2.040 1.040 2.360 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.300 0.500 6.460 1.550 ;
        RECT  4.740 0.500 6.300 0.660 ;
        RECT  4.580 0.440 4.740 0.660 ;
        RECT  1.520 0.440 4.580 0.600 ;
        RECT  1.520 1.380 1.640 1.660 ;
        RECT  1.480 0.440 1.520 1.660 ;
        RECT  1.360 0.440 1.480 1.600 ;
        RECT  1.280 1.240 1.360 1.600 ;
        RECT  0.660 1.440 1.280 1.600 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.380 1.840 19.520 2.560 ;
        RECT  19.320 0.440 19.380 2.560 ;
        RECT  19.110 0.440 19.320 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.700 1.570 6.860 1.870 ;
        RECT  5.920 1.710 6.700 1.870 ;
        RECT  5.700 1.640 5.920 1.960 ;
        RECT  5.680 1.270 5.700 1.960 ;
        RECT  5.540 1.270 5.680 1.800 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.640 3.120 1.960 ;
        RECT  2.880 1.480 3.040 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  9.640 1.240 10.320 1.560 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.850 -0.280 20.000 0.280 ;
        RECT  19.580 -0.280 19.850 1.220 ;
        RECT  18.840 -0.280 19.580 0.280 ;
        RECT  18.680 -0.280 18.840 1.080 ;
        RECT  17.780 -0.280 18.680 0.280 ;
        RECT  17.500 -0.280 17.780 0.340 ;
        RECT  10.900 -0.280 17.500 0.280 ;
        RECT  10.620 -0.280 10.900 0.340 ;
        RECT  10.140 -0.280 10.620 0.280 ;
        RECT  9.860 -0.280 10.140 0.340 ;
        RECT  8.980 -0.280 9.860 0.280 ;
        RECT  8.700 -0.280 8.980 0.340 ;
        RECT  7.320 -0.280 8.700 0.280 ;
        RECT  7.040 -0.280 7.320 0.340 ;
        RECT  6.400 -0.280 7.040 0.280 ;
        RECT  6.120 -0.280 6.400 0.340 ;
        RECT  1.060 -0.280 6.120 0.280 ;
        RECT  0.780 -0.280 1.060 0.340 ;
        RECT  0.000 -0.280 0.780 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.880 3.320 20.000 3.880 ;
        RECT  19.680 1.910 19.880 3.880 ;
        RECT  18.860 3.320 19.680 3.880 ;
        RECT  18.580 3.060 18.860 3.880 ;
        RECT  18.040 3.320 18.580 3.880 ;
        RECT  17.760 2.800 18.040 3.880 ;
        RECT  15.600 3.320 17.760 3.880 ;
        RECT  15.320 3.260 15.600 3.880 ;
        RECT  14.560 3.320 15.320 3.880 ;
        RECT  14.280 3.260 14.560 3.880 ;
        RECT  13.420 3.320 14.280 3.880 ;
        RECT  13.140 3.260 13.420 3.880 ;
        RECT  11.740 3.320 13.140 3.880 ;
        RECT  11.460 3.260 11.740 3.880 ;
        RECT  10.700 3.320 11.460 3.880 ;
        RECT  10.420 3.260 10.700 3.880 ;
        RECT  8.860 3.320 10.420 3.880 ;
        RECT  8.580 3.260 8.860 3.880 ;
        RECT  7.120 3.320 8.580 3.880 ;
        RECT  6.840 3.260 7.120 3.880 ;
        RECT  6.200 3.320 6.840 3.880 ;
        RECT  5.920 2.800 6.200 3.880 ;
        RECT  5.120 3.320 5.920 3.880 ;
        RECT  4.840 3.260 5.120 3.880 ;
        RECT  3.040 3.320 4.840 3.880 ;
        RECT  2.760 3.020 3.040 3.880 ;
        RECT  1.060 3.320 2.760 3.880 ;
        RECT  0.780 3.260 1.060 3.880 ;
        RECT  0.000 3.320 0.780 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  18.360 0.870 18.520 2.560 ;
        RECT  18.320 0.870 18.360 1.030 ;
        RECT  18.340 1.610 18.360 2.560 ;
        RECT  18.160 1.610 18.340 1.890 ;
        RECT  18.160 0.500 18.320 1.030 ;
        RECT  18.000 1.270 18.200 1.430 ;
        RECT  17.300 0.500 18.160 0.660 ;
        RECT  17.840 0.820 18.000 2.490 ;
        RECT  16.980 0.820 17.840 0.980 ;
        RECT  16.080 2.330 17.840 2.490 ;
        RECT  17.520 1.140 17.680 2.170 ;
        RECT  16.460 1.140 17.520 1.300 ;
        RECT  16.620 2.010 17.520 2.170 ;
        RECT  17.200 1.460 17.360 1.850 ;
        RECT  15.920 3.000 17.310 3.160 ;
        RECT  17.140 0.440 17.300 0.660 ;
        RECT  15.180 1.460 17.200 1.620 ;
        RECT  11.220 0.440 17.140 0.600 ;
        RECT  16.820 0.760 16.980 0.980 ;
        RECT  15.660 0.760 16.820 0.920 ;
        RECT  16.330 1.820 16.620 2.170 ;
        RECT  16.180 1.080 16.460 1.300 ;
        RECT  15.080 1.820 16.330 1.980 ;
        RECT  15.500 1.140 16.180 1.300 ;
        RECT  15.920 2.210 16.080 2.490 ;
        RECT  15.760 2.940 15.920 3.160 ;
        RECT  13.100 2.940 15.760 3.100 ;
        RECT  15.340 0.760 15.500 1.300 ;
        RECT  14.790 0.760 15.340 0.920 ;
        RECT  15.020 1.120 15.180 1.620 ;
        RECT  14.810 1.820 15.080 2.780 ;
        RECT  14.120 1.120 15.020 1.280 ;
        RECT  13.800 1.440 14.860 1.600 ;
        RECT  14.790 2.240 14.810 2.780 ;
        RECT  14.330 2.240 14.790 2.400 ;
        RECT  14.170 2.240 14.330 2.580 ;
        RECT  13.960 0.760 14.120 1.280 ;
        RECT  11.540 0.760 13.960 0.920 ;
        RECT  13.640 1.140 13.800 2.180 ;
        RECT  13.580 1.140 13.640 1.300 ;
        RECT  12.520 2.020 13.640 2.180 ;
        RECT  13.420 1.080 13.580 1.300 ;
        RECT  13.280 1.540 13.440 1.820 ;
        RECT  12.340 1.080 13.420 1.240 ;
        RECT  12.180 1.660 13.280 1.820 ;
        RECT  12.940 2.580 13.100 3.100 ;
        RECT  12.180 2.580 12.940 2.740 ;
        RECT  12.180 2.940 12.780 3.100 ;
        RECT  12.360 2.020 12.520 2.330 ;
        RECT  12.020 1.240 12.180 2.740 ;
        RECT  12.010 2.920 12.180 3.100 ;
        RECT  11.700 1.240 12.020 1.400 ;
        RECT  8.420 2.580 12.020 2.740 ;
        RECT  8.100 2.920 12.010 3.080 ;
        RECT  11.540 1.580 11.860 1.860 ;
        RECT  11.380 0.760 11.540 2.400 ;
        RECT  10.940 1.090 11.380 1.250 ;
        RECT  10.720 2.240 11.380 2.400 ;
        RECT  11.060 0.440 11.220 0.660 ;
        RECT  9.780 0.500 11.060 0.660 ;
        RECT  10.660 1.860 11.020 2.020 ;
        RECT  10.530 2.180 10.720 2.400 ;
        RECT  10.500 0.840 10.660 2.020 ;
        RECT  9.480 2.180 10.530 2.340 ;
        RECT  10.380 0.840 10.500 1.000 ;
        RECT  9.320 1.860 10.500 2.020 ;
        RECT  9.620 0.500 9.780 0.980 ;
        RECT  8.970 0.820 9.620 0.980 ;
        RECT  8.420 0.500 9.460 0.660 ;
        RECT  9.160 1.740 9.320 2.020 ;
        RECT  8.800 0.820 8.970 1.120 ;
        RECT  8.580 0.960 8.800 1.120 ;
        RECT  8.260 0.500 8.420 2.740 ;
        RECT  7.940 0.620 8.100 3.080 ;
        RECT  7.820 0.620 7.940 0.780 ;
        RECT  7.920 2.230 7.940 3.080 ;
        RECT  6.520 2.920 7.920 3.080 ;
        RECT  7.760 1.020 7.780 1.940 ;
        RECT  7.620 1.020 7.760 2.740 ;
        RECT  7.600 1.660 7.620 2.740 ;
        RECT  7.400 2.580 7.600 2.740 ;
        RECT  7.180 2.030 7.440 2.190 ;
        RECT  7.020 1.030 7.180 2.190 ;
        RECT  6.780 1.030 7.020 1.190 ;
        RECT  6.760 2.030 7.020 2.190 ;
        RECT  6.620 0.910 6.780 1.190 ;
        RECT  6.360 2.380 6.520 3.080 ;
        RECT  3.980 2.380 6.360 2.540 ;
        RECT  1.520 2.700 5.760 2.860 ;
        RECT  5.380 0.950 5.520 1.110 ;
        RECT  5.380 2.000 5.520 2.160 ;
        RECT  5.220 0.950 5.380 2.160 ;
        RECT  4.620 1.260 5.220 1.420 ;
        RECT  4.840 0.820 5.000 1.100 ;
        RECT  4.420 0.940 4.840 1.100 ;
        RECT  4.420 2.000 4.500 2.160 ;
        RECT  4.260 0.760 4.420 2.160 ;
        RECT  2.280 0.760 4.260 0.920 ;
        RECT  4.140 1.410 4.260 1.570 ;
        RECT  4.220 2.000 4.260 2.160 ;
        RECT  3.980 1.080 4.100 1.240 ;
        RECT  3.820 1.080 3.980 2.540 ;
        RECT  1.960 2.380 3.820 2.540 ;
        RECT  3.560 1.080 3.640 1.240 ;
        RECT  3.400 1.080 3.560 2.220 ;
        RECT  2.600 1.080 3.400 1.240 ;
        RECT  3.280 2.060 3.400 2.220 ;
        RECT  2.440 1.080 2.600 2.220 ;
        RECT  2.240 2.060 2.440 2.220 ;
        RECT  2.120 0.760 2.280 1.640 ;
        RECT  1.800 1.060 1.960 2.540 ;
        RECT  1.680 1.060 1.800 1.220 ;
        RECT  1.680 2.260 1.800 2.540 ;
        RECT  1.520 1.820 1.640 2.100 ;
        RECT  1.360 1.820 1.520 2.860 ;
        RECT  0.560 2.700 1.360 2.860 ;
        RECT  0.500 1.000 0.560 1.280 ;
        RECT  0.500 2.150 0.560 2.860 ;
        RECT  0.400 1.000 0.500 2.860 ;
        RECT  0.340 1.000 0.400 2.430 ;
    END
END SEDFFHQX4TR

MACRO SEDFFHQX2TR
    CLASS CORE ;
    FOREIGN SEDFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.640 1.160 1.960 ;
        RECT  0.880 1.550 1.130 1.960 ;
        RECT  0.850 1.550 0.880 1.830 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.210 4.980 1.490 ;
        RECT  4.520 0.440 4.680 1.490 ;
        RECT  1.450 0.440 4.520 0.600 ;
        RECT  1.170 0.440 1.450 0.750 ;
        RECT  0.760 0.590 1.170 0.750 ;
        RECT  0.690 0.590 0.760 1.160 ;
        RECT  0.600 0.590 0.690 1.640 ;
        RECT  0.470 0.840 0.600 1.640 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.710 0.520 14.990 3.080 ;
        RECT  14.480 1.990 14.710 2.650 ;
        RECT  13.870 2.420 14.480 2.650 ;
        RECT  13.590 2.420 13.870 2.940 ;
        END
        ANTENNADIFFAREA 3.392 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.160 1.530 5.380 1.810 ;
        RECT  4.360 1.650 5.160 1.810 ;
        RECT  3.890 1.240 4.360 1.830 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.620 2.760 2.000 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  7.480 1.240 7.960 1.560 ;
        END
        ANTENNAGATEAREA 0.2184 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.510 -0.280 15.200 0.280 ;
        RECT  14.230 -0.280 14.510 1.080 ;
        RECT  13.610 -0.280 14.230 0.280 ;
        RECT  13.330 -0.280 13.610 0.340 ;
        RECT  9.430 -0.280 13.330 0.280 ;
        RECT  9.150 -0.280 9.430 0.360 ;
        RECT  7.130 -0.280 9.150 0.340 ;
        RECT  6.850 -0.280 7.130 0.380 ;
        RECT  5.670 -0.280 6.850 0.340 ;
        RECT  5.390 -0.280 5.670 0.400 ;
        RECT  0.810 -0.280 5.390 0.280 ;
        RECT  0.530 -0.280 0.810 0.400 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.380 3.320 15.200 3.880 ;
        RECT  14.100 2.830 14.380 3.880 ;
        RECT  13.350 3.320 14.100 3.880 ;
        RECT  13.070 1.970 13.350 3.880 ;
        RECT  11.510 3.320 13.070 3.880 ;
        RECT  11.230 3.200 11.510 3.880 ;
        RECT  8.660 3.320 11.230 3.880 ;
        RECT  8.380 3.200 8.660 3.880 ;
        RECT  7.180 3.320 8.380 3.880 ;
        RECT  6.900 3.200 7.180 3.880 ;
        RECT  4.860 3.320 6.900 3.880 ;
        RECT  4.580 2.800 4.860 3.880 ;
        RECT  3.710 3.260 4.580 3.880 ;
        RECT  3.430 3.200 3.710 3.880 ;
        RECT  2.770 3.320 3.430 3.880 ;
        RECT  2.490 2.980 2.770 3.880 ;
        RECT  0.850 3.260 2.490 3.880 ;
        RECT  0.570 3.200 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.930 0.800 13.990 1.080 ;
        RECT  13.770 0.500 13.930 2.200 ;
        RECT  12.950 0.500 13.770 0.660 ;
        RECT  13.590 1.640 13.770 2.200 ;
        RECT  13.450 0.820 13.610 1.410 ;
        RECT  12.990 1.640 13.590 1.800 ;
        RECT  12.630 0.820 13.450 0.980 ;
        RECT  12.790 0.440 12.950 0.660 ;
        RECT  12.830 1.140 12.950 1.420 ;
        RECT  12.830 2.760 12.890 3.040 ;
        RECT  12.670 1.140 12.830 3.040 ;
        RECT  9.750 0.440 12.790 0.600 ;
        RECT  10.940 2.880 12.670 3.040 ;
        RECT  12.510 0.760 12.630 0.980 ;
        RECT  12.350 0.760 12.510 2.720 ;
        RECT  12.230 1.930 12.350 2.720 ;
        RECT  12.030 0.760 12.190 1.730 ;
        RECT  11.550 0.760 12.030 0.970 ;
        RECT  11.870 1.570 12.030 2.480 ;
        RECT  11.650 1.130 11.870 1.410 ;
        RECT  11.750 2.180 11.870 2.480 ;
        RECT  11.320 2.320 11.750 2.480 ;
        RECT  11.390 1.130 11.650 1.290 ;
        RECT  11.070 1.470 11.470 1.750 ;
        RECT  11.230 0.760 11.390 1.290 ;
        RECT  11.100 2.320 11.320 2.600 ;
        RECT  10.070 0.760 11.230 0.920 ;
        RECT  10.910 1.140 11.070 2.160 ;
        RECT  10.780 2.560 10.940 3.040 ;
        RECT  10.230 1.140 10.910 1.300 ;
        RECT  10.510 2.000 10.910 2.160 ;
        RECT  10.070 2.560 10.780 2.720 ;
        RECT  10.070 1.680 10.750 1.840 ;
        RECT  10.340 2.880 10.620 3.160 ;
        RECT  10.290 2.000 10.510 2.280 ;
        RECT  6.460 2.880 10.340 3.040 ;
        RECT  9.910 0.760 10.070 1.030 ;
        RECT  9.910 1.340 10.070 2.720 ;
        RECT  9.370 0.870 9.910 1.030 ;
        RECT  9.810 1.340 9.910 1.500 ;
        RECT  7.320 2.500 9.910 2.720 ;
        RECT  9.530 1.190 9.810 1.500 ;
        RECT  9.590 0.440 9.750 0.700 ;
        RECT  9.370 1.660 9.750 1.940 ;
        RECT  7.000 0.540 9.590 0.700 ;
        RECT  9.210 0.870 9.370 1.940 ;
        RECT  9.120 0.870 9.210 1.140 ;
        RECT  9.120 1.780 9.210 1.940 ;
        RECT  8.840 0.860 9.120 1.140 ;
        RECT  8.960 1.780 9.120 2.340 ;
        RECT  8.510 1.300 9.050 1.580 ;
        RECT  8.840 2.060 8.960 2.340 ;
        RECT  7.820 2.180 8.840 2.340 ;
        RECT  8.350 0.860 8.510 2.020 ;
        RECT  8.230 0.860 8.350 1.140 ;
        RECT  7.980 1.800 8.350 2.020 ;
        RECT  7.540 1.720 7.820 2.340 ;
        RECT  7.320 0.860 7.650 1.080 ;
        RECT  7.160 0.860 7.320 2.720 ;
        RECT  6.780 0.540 7.000 1.410 ;
        RECT  6.460 0.670 6.620 2.370 ;
        RECT  6.230 0.670 6.460 0.830 ;
        RECT  6.340 2.210 6.460 3.040 ;
        RECT  6.180 2.210 6.340 3.160 ;
        RECT  6.020 1.010 6.300 2.050 ;
        RECT  5.950 0.550 6.230 0.830 ;
        RECT  5.180 3.000 6.180 3.160 ;
        RECT  5.950 1.010 6.020 1.290 ;
        RECT  5.860 1.890 6.020 2.840 ;
        RECT  5.700 1.450 5.860 1.730 ;
        RECT  5.720 2.560 5.860 2.840 ;
        RECT  5.540 0.890 5.700 2.250 ;
        RECT  5.220 0.890 5.540 1.050 ;
        RECT  5.300 1.970 5.540 2.250 ;
        RECT  4.940 0.770 5.220 1.050 ;
        RECT  5.020 2.430 5.180 3.160 ;
        RECT  3.410 2.430 5.020 2.590 ;
        RECT  3.090 2.750 4.420 3.030 ;
        RECT  3.730 1.990 4.270 2.270 ;
        RECT  3.730 0.800 3.900 1.080 ;
        RECT  3.570 0.800 3.730 2.270 ;
        RECT  3.300 1.460 3.570 1.740 ;
        RECT  3.250 2.340 3.410 2.590 ;
        RECT  3.140 1.900 3.370 2.180 ;
        RECT  3.140 1.010 3.310 1.300 ;
        RECT  1.730 2.340 3.250 2.500 ;
        RECT  3.030 1.010 3.140 2.180 ;
        RECT  2.930 2.660 3.090 3.030 ;
        RECT  2.980 1.140 3.030 2.180 ;
        RECT  2.330 1.140 2.980 1.300 ;
        RECT  1.490 2.660 2.930 2.820 ;
        RECT  1.950 0.760 2.410 0.980 ;
        RECT  2.110 1.140 2.330 1.420 ;
        RECT  1.950 1.580 2.210 2.180 ;
        RECT  1.930 0.760 1.950 2.180 ;
        RECT  1.790 0.760 1.930 1.740 ;
        RECT  1.630 2.220 1.730 2.500 ;
        RECT  1.410 0.910 1.630 2.500 ;
        RECT  1.210 2.660 1.490 2.940 ;
        RECT  0.310 2.660 1.210 2.820 ;
        RECT  0.150 1.030 0.310 2.820 ;
        RECT  0.090 1.030 0.150 1.310 ;
        RECT  0.090 1.910 0.150 2.190 ;
    END
END SEDFFHQX2TR

MACRO SEDFFHQX1TR
    CLASS CORE ;
    FOREIGN SEDFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.500 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.330 4.910 1.550 ;
        RECT  4.520 0.500 4.680 1.550 ;
        RECT  1.530 0.500 4.520 0.660 ;
        RECT  1.170 0.500 1.530 0.780 ;
        RECT  0.720 0.620 1.170 0.780 ;
        RECT  0.690 0.620 0.720 1.160 ;
        RECT  0.470 0.620 0.690 1.710 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.160 1.020 14.320 2.660 ;
        RECT  14.040 1.020 14.160 1.300 ;
        RECT  13.960 2.370 14.160 2.660 ;
        RECT  13.680 2.370 13.960 3.150 ;
        END
        ANTENNADIFFAREA 2.482 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.070 1.490 5.350 1.870 ;
        RECT  4.360 1.710 5.070 1.870 ;
        RECT  3.880 1.640 4.360 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.640 2.760 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  7.420 1.240 7.960 1.680 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.470 -0.280 14.400 0.280 ;
        RECT  13.190 -0.280 13.470 0.340 ;
        RECT  9.070 -0.280 13.190 0.280 ;
        RECT  7.130 -0.280 9.070 0.340 ;
        RECT  6.850 -0.280 7.130 0.360 ;
        RECT  5.590 -0.280 6.850 0.340 ;
        RECT  5.310 -0.280 5.590 0.400 ;
        RECT  3.090 -0.280 5.310 0.340 ;
        RECT  1.270 -0.280 3.090 0.280 ;
        RECT  0.810 -0.280 1.270 0.340 ;
        RECT  0.530 -0.280 0.810 0.400 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.480 3.320 14.400 3.880 ;
        RECT  13.200 2.370 13.480 3.880 ;
        RECT  7.190 3.320 13.200 3.880 ;
        RECT  6.910 3.260 7.190 3.880 ;
        RECT  4.830 3.320 6.910 3.880 ;
        RECT  4.550 2.860 4.830 3.880 ;
        RECT  3.690 3.260 4.550 3.880 ;
        RECT  3.410 3.200 3.690 3.880 ;
        RECT  2.740 3.320 3.410 3.880 ;
        RECT  2.490 2.960 2.740 3.880 ;
        RECT  0.810 3.260 2.490 3.880 ;
        RECT  0.530 3.200 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.880 0.440 14.030 0.660 ;
        RECT  13.880 1.910 14.000 2.190 ;
        RECT  13.720 0.440 13.880 2.190 ;
        RECT  12.410 0.500 13.720 0.660 ;
        RECT  12.950 1.860 13.720 2.190 ;
        RECT  13.340 0.880 13.560 1.650 ;
        RECT  12.530 0.880 13.340 1.040 ;
        RECT  12.630 1.200 12.790 3.160 ;
        RECT  12.570 1.200 12.630 1.480 ;
        RECT  12.400 2.880 12.630 3.160 ;
        RECT  12.410 0.820 12.530 1.040 ;
        RECT  12.410 2.190 12.470 2.470 ;
        RECT  12.250 0.440 12.410 0.660 ;
        RECT  12.250 0.820 12.410 2.470 ;
        RECT  11.910 2.880 12.400 3.060 ;
        RECT  9.670 0.440 12.250 0.600 ;
        RECT  11.930 0.760 12.090 2.470 ;
        RECT  11.570 0.760 11.930 1.040 ;
        RECT  11.710 2.190 11.930 2.470 ;
        RECT  10.730 2.900 11.910 3.060 ;
        RECT  11.550 1.200 11.770 1.480 ;
        RECT  11.410 2.310 11.710 2.470 ;
        RECT  11.090 1.680 11.580 1.960 ;
        RECT  11.410 1.200 11.550 1.360 ;
        RECT  11.250 0.760 11.410 1.360 ;
        RECT  11.250 2.310 11.410 2.740 ;
        RECT  9.990 0.760 11.250 0.920 ;
        RECT  10.890 2.460 11.250 2.740 ;
        RECT  10.930 1.090 11.090 2.300 ;
        RECT  10.150 1.090 10.930 1.310 ;
        RECT  10.530 2.140 10.930 2.300 ;
        RECT  10.090 1.700 10.770 1.980 ;
        RECT  10.570 2.590 10.730 3.060 ;
        RECT  10.090 2.590 10.570 2.750 ;
        RECT  10.250 2.140 10.530 2.420 ;
        RECT  9.930 2.910 10.210 3.130 ;
        RECT  9.930 1.530 10.090 2.750 ;
        RECT  9.830 0.760 9.990 1.000 ;
        RECT  9.790 1.530 9.930 1.690 ;
        RECT  7.260 2.590 9.930 2.750 ;
        RECT  6.540 2.910 9.930 3.070 ;
        RECT  9.350 0.840 9.830 1.000 ;
        RECT  9.510 1.160 9.790 1.690 ;
        RECT  9.350 1.850 9.770 2.070 ;
        RECT  9.510 0.440 9.670 0.680 ;
        RECT  6.900 0.520 9.510 0.680 ;
        RECT  9.190 0.840 9.350 2.430 ;
        RECT  8.650 0.840 9.190 1.120 ;
        RECT  7.830 2.270 9.190 2.430 ;
        RECT  8.470 1.410 9.030 1.690 ;
        RECT  8.190 1.010 8.470 2.110 ;
        RECT  7.990 1.890 8.190 2.110 ;
        RECT  7.550 1.840 7.830 2.430 ;
        RECT  7.260 0.840 7.570 1.060 ;
        RECT  7.100 0.840 7.260 2.750 ;
        RECT  6.700 0.520 6.900 1.840 ;
        RECT  6.380 0.550 6.540 3.070 ;
        RECT  5.910 0.550 6.380 0.830 ;
        RECT  6.310 2.320 6.380 3.070 ;
        RECT  6.150 2.320 6.310 3.160 ;
        RECT  5.990 1.010 6.220 2.160 ;
        RECT  5.150 3.000 6.150 3.160 ;
        RECT  5.950 1.010 5.990 2.840 ;
        RECT  5.870 1.010 5.950 1.290 ;
        RECT  5.830 2.000 5.950 2.840 ;
        RECT  5.690 2.560 5.830 2.840 ;
        RECT  5.670 1.450 5.790 1.730 ;
        RECT  5.510 0.830 5.670 2.250 ;
        RECT  4.870 0.830 5.510 1.110 ;
        RECT  5.270 2.030 5.510 2.250 ;
        RECT  4.990 2.500 5.150 3.160 ;
        RECT  3.400 2.500 4.990 2.660 ;
        RECT  3.080 2.820 4.390 3.040 ;
        RECT  3.720 2.120 4.250 2.340 ;
        RECT  3.720 0.940 3.830 1.220 ;
        RECT  3.560 0.940 3.720 2.340 ;
        RECT  3.550 0.940 3.560 1.780 ;
        RECT  3.240 1.520 3.550 1.780 ;
        RECT  3.240 2.320 3.400 2.660 ;
        RECT  3.080 1.940 3.350 2.160 ;
        RECT  3.080 1.010 3.240 1.360 ;
        RECT  1.730 2.320 3.240 2.480 ;
        RECT  2.960 1.010 3.080 2.160 ;
        RECT  2.920 2.640 3.080 3.040 ;
        RECT  2.920 1.200 2.960 2.160 ;
        RECT  2.330 1.200 2.920 1.360 ;
        RECT  0.370 2.640 2.920 2.800 ;
        RECT  1.950 0.820 2.410 1.040 ;
        RECT  2.110 1.200 2.330 1.480 ;
        RECT  1.950 1.640 2.210 2.120 ;
        RECT  1.930 0.820 1.950 2.120 ;
        RECT  1.790 0.820 1.930 1.800 ;
        RECT  1.630 1.960 1.730 2.480 ;
        RECT  1.410 0.940 1.630 2.480 ;
        RECT  0.250 1.910 0.370 2.800 ;
        RECT  0.250 1.030 0.310 1.310 ;
        RECT  0.210 1.030 0.250 2.800 ;
        RECT  0.090 1.030 0.210 2.190 ;
    END
END SEDFFHQX1TR

MACRO SEDFFXLTR
    CLASS CORE ;
    FOREIGN SEDFFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.570 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.530 1.120 1.960 ;
        RECT  0.880 1.510 1.040 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.880 0.460 11.120 2.230 ;
        END
        ANTENNADIFFAREA 1.7195 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.560 0.640 10.720 2.760 ;
        RECT  9.940 0.640 10.560 0.800 ;
        RECT  10.480 2.420 10.560 2.760 ;
        RECT  10.080 2.600 10.480 2.760 ;
        RECT  9.920 2.600 10.080 2.880 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 2.440 0.760 2.600 ;
        RECT  0.360 2.440 0.720 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.610 3.120 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.850 6.320 2.360 ;
        RECT  5.930 1.850 6.080 2.010 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.580 -0.280 11.200 0.280 ;
        RECT  10.300 -0.280 10.580 0.340 ;
        RECT  9.700 -0.280 10.300 0.280 ;
        RECT  9.420 -0.280 9.700 0.340 ;
        RECT  7.970 -0.280 9.420 0.280 ;
        RECT  7.810 -0.280 7.970 1.050 ;
        RECT  6.400 -0.280 7.810 0.280 ;
        RECT  5.680 -0.280 6.400 0.650 ;
        RECT  2.320 -0.280 5.680 0.280 ;
        RECT  2.160 -0.280 2.320 0.740 ;
        RECT  0.880 -0.280 2.160 0.280 ;
        RECT  0.600 -0.280 0.880 0.340 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.320 11.200 3.880 ;
        RECT  10.420 3.260 10.700 3.880 ;
        RECT  9.560 3.320 10.420 3.880 ;
        RECT  9.400 2.930 9.560 3.880 ;
        RECT  7.920 3.320 9.400 3.880 ;
        RECT  7.250 3.260 7.920 3.880 ;
        RECT  6.380 3.320 7.250 3.880 ;
        RECT  5.780 3.260 6.380 3.880 ;
        RECT  1.840 3.320 5.780 3.880 ;
        RECT  1.680 2.860 1.840 3.880 ;
        RECT  0.880 3.320 1.680 3.880 ;
        RECT  0.600 2.920 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.240 1.430 10.370 1.720 ;
        RECT  10.220 1.070 10.240 1.720 ;
        RECT  10.060 1.070 10.220 2.330 ;
        RECT  9.960 1.070 10.060 1.290 ;
        RECT  9.900 2.010 10.060 2.330 ;
        RECT  9.120 2.010 9.900 2.170 ;
        RECT  9.720 1.570 9.880 1.850 ;
        RECT  8.860 1.690 9.720 1.850 ;
        RECT  8.880 0.480 9.160 0.670 ;
        RECT  8.960 2.010 9.120 3.100 ;
        RECT  4.240 2.940 8.960 3.100 ;
        RECT  8.460 0.510 8.880 0.670 ;
        RECT  8.800 0.830 8.860 1.850 ;
        RECT  8.700 0.830 8.800 2.670 ;
        RECT  8.640 1.690 8.700 2.670 ;
        RECT  8.600 2.340 8.640 2.670 ;
        RECT  8.440 0.510 8.460 1.830 ;
        RECT  8.300 0.510 8.440 2.680 ;
        RECT  8.280 1.550 8.300 2.680 ;
        RECT  5.920 2.520 8.280 2.680 ;
        RECT  7.960 1.290 8.120 2.170 ;
        RECT  7.490 1.290 7.960 1.450 ;
        RECT  7.250 2.010 7.960 2.170 ;
        RECT  7.070 1.660 7.800 1.820 ;
        RECT  7.330 0.560 7.490 1.450 ;
        RECT  6.990 0.560 7.330 0.720 ;
        RECT  6.910 0.960 7.070 1.820 ;
        RECT  6.830 0.440 6.990 0.720 ;
        RECT  6.840 1.530 6.910 1.820 ;
        RECT  6.680 1.530 6.840 2.310 ;
        RECT  5.660 1.530 6.680 1.690 ;
        RECT  6.510 0.810 6.670 1.350 ;
        RECT  5.020 0.810 6.510 0.970 ;
        RECT  5.340 1.160 5.960 1.320 ;
        RECT  5.760 2.170 5.920 2.680 ;
        RECT  5.340 2.220 5.760 2.380 ;
        RECT  5.500 1.530 5.660 1.810 ;
        RECT  5.180 1.160 5.340 2.380 ;
        RECT  5.120 1.500 5.180 2.380 ;
        RECT  4.780 1.500 5.120 1.660 ;
        RECT  4.860 2.620 5.100 2.780 ;
        RECT  4.860 0.810 5.020 1.090 ;
        RECT  4.440 0.930 4.860 1.090 ;
        RECT  4.700 1.820 4.860 2.780 ;
        RECT  4.620 1.380 4.780 1.660 ;
        RECT  4.440 1.820 4.700 1.980 ;
        RECT  4.400 0.460 4.560 0.740 ;
        RECT  2.500 2.440 4.540 2.600 ;
        RECT  4.280 0.930 4.440 1.980 ;
        RECT  2.920 0.460 4.400 0.620 ;
        RECT  4.080 2.760 4.240 3.100 ;
        RECT  3.440 1.360 3.980 1.520 ;
        RECT  2.000 0.910 3.740 1.070 ;
        RECT  2.160 2.760 3.660 2.920 ;
        RECT  3.440 2.110 3.560 2.270 ;
        RECT  3.280 1.230 3.440 2.270 ;
        RECT  1.680 1.230 3.280 1.390 ;
        RECT  2.760 0.460 2.920 0.740 ;
        RECT  2.480 1.940 2.640 2.280 ;
        RECT  1.680 2.120 2.480 2.280 ;
        RECT  2.000 2.540 2.160 2.920 ;
        RECT  1.840 0.490 2.000 1.070 ;
        RECT  1.340 2.540 2.000 2.700 ;
        RECT  1.340 0.490 1.840 0.650 ;
        RECT  1.520 0.810 1.680 1.390 ;
        RECT  1.520 1.550 1.680 2.280 ;
        RECT  0.340 0.810 1.520 0.970 ;
        RECT  1.320 1.950 1.520 2.280 ;
        RECT  1.180 2.540 1.340 2.790 ;
        RECT  0.680 1.130 1.320 1.290 ;
        RECT  0.680 2.120 1.320 2.280 ;
        RECT  1.060 2.630 1.180 2.790 ;
        RECT  0.520 1.130 0.680 2.280 ;
        RECT  0.180 0.520 0.340 2.230 ;
    END
END SEDFFXLTR

MACRO SEDFFX4TR
    CLASS CORE ;
    FOREIGN SEDFFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.570 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.530 1.160 1.960 ;
        RECT  0.840 1.510 1.040 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.680 0.520 11.920 3.070 ;
        RECT  11.610 0.520 11.680 1.360 ;
        RECT  11.610 1.910 11.680 3.070 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.290 0.500 11.450 2.730 ;
        RECT  9.940 0.500 11.290 0.720 ;
        RECT  10.320 2.570 11.290 2.730 ;
        RECT  10.150 2.240 10.320 2.960 ;
        RECT  10.070 2.210 10.150 2.960 ;
        RECT  9.910 2.210 10.070 3.030 ;
        END
        ANTENNADIFFAREA 4.18 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 2.440 0.760 2.600 ;
        RECT  0.360 2.440 0.720 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.610 3.120 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.850 6.320 2.360 ;
        RECT  5.930 1.850 6.080 2.010 ;
        END
        ANTENNAGATEAREA 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.250 -0.280 12.400 0.280 ;
        RECT  12.090 -0.280 12.250 1.310 ;
        RECT  11.250 -0.280 12.090 0.280 ;
        RECT  10.970 -0.280 11.250 0.340 ;
        RECT  9.680 -0.280 10.970 0.280 ;
        RECT  9.400 -0.280 9.680 0.340 ;
        RECT  7.990 -0.280 9.400 0.280 ;
        RECT  7.830 -0.280 7.990 1.050 ;
        RECT  6.400 -0.280 7.830 0.280 ;
        RECT  5.680 -0.280 6.400 0.650 ;
        RECT  2.320 -0.280 5.680 0.280 ;
        RECT  2.160 -0.280 2.320 0.740 ;
        RECT  0.880 -0.280 2.160 0.280 ;
        RECT  0.600 -0.280 0.880 0.340 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.250 3.320 12.400 3.880 ;
        RECT  12.090 1.930 12.250 3.880 ;
        RECT  11.250 3.320 12.090 3.880 ;
        RECT  10.480 3.260 11.250 3.880 ;
        RECT  9.590 3.320 10.480 3.880 ;
        RECT  9.430 2.930 9.590 3.880 ;
        RECT  8.000 3.320 9.430 3.880 ;
        RECT  7.720 3.260 8.000 3.880 ;
        RECT  6.380 3.320 7.720 3.880 ;
        RECT  5.780 3.260 6.380 3.880 ;
        RECT  1.840 3.320 5.780 3.880 ;
        RECT  1.680 2.860 1.840 3.880 ;
        RECT  0.880 3.320 1.680 3.880 ;
        RECT  0.600 2.920 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.950 1.170 11.130 1.970 ;
        RECT  9.950 1.170 10.950 1.330 ;
        RECT  10.670 1.810 10.950 2.260 ;
        RECT  8.910 1.490 10.750 1.650 ;
        RECT  9.230 1.810 10.670 1.970 ;
        RECT  9.070 1.810 9.230 3.100 ;
        RECT  8.840 0.480 9.120 0.670 ;
        RECT  4.240 2.940 9.070 3.100 ;
        RECT  8.750 0.830 8.910 2.670 ;
        RECT  8.460 0.510 8.840 0.670 ;
        RECT  8.660 0.830 8.750 1.130 ;
        RECT  8.620 2.340 8.750 2.670 ;
        RECT  8.460 1.850 8.580 2.140 ;
        RECT  8.300 0.510 8.460 2.780 ;
        RECT  5.920 2.620 8.300 2.780 ;
        RECT  7.800 1.500 7.960 2.410 ;
        RECT  7.510 1.500 7.800 1.660 ;
        RECT  7.290 2.250 7.800 2.410 ;
        RECT  7.070 1.820 7.640 1.980 ;
        RECT  7.350 0.560 7.510 1.660 ;
        RECT  6.990 0.560 7.350 0.720 ;
        RECT  6.910 0.960 7.070 1.980 ;
        RECT  6.830 0.440 6.990 0.720 ;
        RECT  6.840 1.530 6.910 1.980 ;
        RECT  6.680 1.530 6.840 2.310 ;
        RECT  5.660 1.530 6.680 1.690 ;
        RECT  6.510 0.810 6.670 1.350 ;
        RECT  5.020 0.810 6.510 0.970 ;
        RECT  5.340 1.160 5.960 1.320 ;
        RECT  5.760 2.170 5.920 2.780 ;
        RECT  5.340 2.220 5.760 2.380 ;
        RECT  5.500 1.530 5.660 1.810 ;
        RECT  5.180 1.160 5.340 2.380 ;
        RECT  5.120 1.500 5.180 2.380 ;
        RECT  4.780 1.500 5.120 1.660 ;
        RECT  4.860 2.620 5.100 2.780 ;
        RECT  4.860 0.810 5.020 1.090 ;
        RECT  4.440 0.930 4.860 1.090 ;
        RECT  4.700 1.820 4.860 2.780 ;
        RECT  4.620 1.380 4.780 1.660 ;
        RECT  4.440 1.820 4.700 1.980 ;
        RECT  4.400 0.460 4.560 0.740 ;
        RECT  2.500 2.440 4.540 2.600 ;
        RECT  4.280 0.930 4.440 1.980 ;
        RECT  2.920 0.460 4.400 0.620 ;
        RECT  4.080 2.760 4.240 3.100 ;
        RECT  3.440 1.360 3.980 1.520 ;
        RECT  2.000 0.910 3.740 1.070 ;
        RECT  2.160 2.760 3.660 2.920 ;
        RECT  3.440 2.110 3.560 2.270 ;
        RECT  3.280 1.230 3.440 2.270 ;
        RECT  1.680 1.230 3.280 1.390 ;
        RECT  2.760 0.460 2.920 0.740 ;
        RECT  2.480 1.940 2.640 2.280 ;
        RECT  1.680 2.120 2.480 2.280 ;
        RECT  2.000 2.540 2.160 2.920 ;
        RECT  1.840 0.490 2.000 1.070 ;
        RECT  1.340 2.540 2.000 2.700 ;
        RECT  1.310 0.490 1.840 0.650 ;
        RECT  1.520 0.810 1.680 1.390 ;
        RECT  1.520 1.550 1.680 2.280 ;
        RECT  0.340 0.810 1.520 0.970 ;
        RECT  1.320 1.950 1.520 2.280 ;
        RECT  1.180 2.540 1.340 2.790 ;
        RECT  0.680 1.130 1.320 1.290 ;
        RECT  0.680 2.120 1.320 2.280 ;
        RECT  1.060 2.630 1.180 2.790 ;
        RECT  0.520 1.130 0.680 2.280 ;
        RECT  0.180 0.520 0.340 2.230 ;
    END
END SEDFFX4TR

MACRO SEDFFX2TR
    CLASS CORE ;
    FOREIGN SEDFFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.570 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 2.030 1.120 2.360 ;
        RECT  0.880 1.620 1.040 2.360 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 0.520 11.520 3.070 ;
        END
        ANTENNADIFFAREA 3.456 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.960 0.500 11.120 2.730 ;
        RECT  9.940 0.500 10.960 0.720 ;
        RECT  10.260 2.570 10.960 2.730 ;
        RECT  10.100 2.570 10.260 3.160 ;
        RECT  9.940 2.440 10.100 3.160 ;
        RECT  9.680 2.440 9.940 2.760 ;
        END
        ANTENNADIFFAREA 3.057 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 2.440 0.720 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.610 3.120 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.850 6.320 2.360 ;
        RECT  5.930 1.850 6.080 2.010 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.920 -0.280 11.600 0.280 ;
        RECT  10.640 -0.280 10.920 0.340 ;
        RECT  9.720 -0.280 10.640 0.280 ;
        RECT  9.440 -0.280 9.720 0.340 ;
        RECT  7.990 -0.280 9.440 0.280 ;
        RECT  7.830 -0.280 7.990 1.050 ;
        RECT  6.400 -0.280 7.830 0.280 ;
        RECT  5.680 -0.280 6.400 0.650 ;
        RECT  2.320 -0.280 5.680 0.280 ;
        RECT  2.160 -0.280 2.320 0.740 ;
        RECT  0.880 -0.280 2.160 0.280 ;
        RECT  0.600 -0.280 0.880 0.340 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.980 3.320 11.600 3.880 ;
        RECT  10.700 3.260 10.980 3.880 ;
        RECT  9.690 3.320 10.700 3.880 ;
        RECT  9.400 2.930 9.690 3.880 ;
        RECT  7.970 3.320 9.400 3.880 ;
        RECT  7.270 3.260 7.970 3.880 ;
        RECT  6.380 3.320 7.270 3.880 ;
        RECT  5.780 3.260 6.380 3.880 ;
        RECT  1.840 3.320 5.780 3.880 ;
        RECT  1.680 2.860 1.840 3.880 ;
        RECT  0.880 3.320 1.680 3.880 ;
        RECT  0.600 2.920 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.640 1.200 10.800 2.170 ;
        RECT  9.980 1.200 10.640 1.360 ;
        RECT  10.560 2.010 10.640 2.170 ;
        RECT  10.340 2.010 10.560 2.390 ;
        RECT  9.140 2.010 10.340 2.170 ;
        RECT  9.740 1.570 9.900 1.850 ;
        RECT  8.880 1.690 9.740 1.850 ;
        RECT  8.900 0.480 9.180 0.670 ;
        RECT  8.980 2.010 9.140 3.100 ;
        RECT  4.240 2.940 8.980 3.100 ;
        RECT  8.480 0.510 8.900 0.670 ;
        RECT  8.820 0.830 8.880 1.850 ;
        RECT  8.720 0.830 8.820 2.670 ;
        RECT  8.660 1.690 8.720 2.670 ;
        RECT  8.620 2.340 8.660 2.670 ;
        RECT  8.460 0.510 8.480 1.830 ;
        RECT  8.320 0.510 8.460 2.680 ;
        RECT  8.300 1.550 8.320 2.680 ;
        RECT  5.920 2.520 8.300 2.680 ;
        RECT  7.980 1.290 8.140 2.170 ;
        RECT  7.510 1.290 7.980 1.450 ;
        RECT  7.270 2.010 7.980 2.170 ;
        RECT  7.070 1.660 7.820 1.820 ;
        RECT  7.350 0.560 7.510 1.450 ;
        RECT  6.990 0.560 7.350 0.720 ;
        RECT  6.910 0.960 7.070 1.820 ;
        RECT  6.830 0.440 6.990 0.720 ;
        RECT  6.840 1.530 6.910 1.820 ;
        RECT  6.680 1.530 6.840 2.310 ;
        RECT  5.660 1.530 6.680 1.690 ;
        RECT  6.510 0.810 6.670 1.350 ;
        RECT  5.020 0.810 6.510 0.970 ;
        RECT  5.340 1.160 5.960 1.320 ;
        RECT  5.760 2.170 5.920 2.680 ;
        RECT  5.340 2.220 5.760 2.380 ;
        RECT  5.500 1.530 5.660 1.810 ;
        RECT  5.180 1.160 5.340 2.380 ;
        RECT  5.120 1.500 5.180 2.380 ;
        RECT  4.780 1.500 5.120 1.660 ;
        RECT  4.860 2.620 5.100 2.780 ;
        RECT  4.860 0.810 5.020 1.090 ;
        RECT  4.440 0.930 4.860 1.090 ;
        RECT  4.700 1.820 4.860 2.780 ;
        RECT  4.620 1.380 4.780 1.660 ;
        RECT  4.440 1.820 4.700 1.980 ;
        RECT  4.400 0.460 4.560 0.740 ;
        RECT  2.500 2.440 4.540 2.600 ;
        RECT  4.280 0.930 4.440 1.980 ;
        RECT  2.920 0.460 4.400 0.620 ;
        RECT  4.080 2.760 4.240 3.100 ;
        RECT  3.440 1.360 3.980 1.520 ;
        RECT  2.000 0.910 3.740 1.070 ;
        RECT  2.160 2.760 3.660 2.920 ;
        RECT  3.440 2.110 3.560 2.270 ;
        RECT  3.280 1.230 3.440 2.270 ;
        RECT  1.680 1.230 3.280 1.390 ;
        RECT  2.760 0.460 2.920 0.740 ;
        RECT  2.480 1.940 2.640 2.280 ;
        RECT  1.520 2.120 2.480 2.280 ;
        RECT  2.000 2.540 2.160 2.920 ;
        RECT  1.840 0.490 2.000 1.070 ;
        RECT  1.340 2.540 2.000 2.700 ;
        RECT  1.310 0.490 1.840 0.650 ;
        RECT  1.520 0.810 1.680 1.390 ;
        RECT  1.520 1.550 1.680 1.820 ;
        RECT  0.340 0.810 1.520 0.970 ;
        RECT  1.360 1.550 1.520 2.280 ;
        RECT  1.320 1.130 1.360 2.280 ;
        RECT  1.180 2.540 1.340 2.790 ;
        RECT  1.200 1.130 1.320 1.810 ;
        RECT  0.520 1.130 1.200 1.290 ;
        RECT  1.060 2.630 1.180 2.790 ;
        RECT  0.180 0.520 0.340 2.230 ;
    END
END SEDFFX2TR

MACRO SEDFFX1TR
    CLASS CORE ;
    FOREIGN SEDFFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.570 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.530 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.880 0.840 11.120 2.230 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.560 0.510 10.720 2.760 ;
        RECT  10.230 0.510 10.560 0.720 ;
        RECT  10.480 2.410 10.560 2.760 ;
        RECT  10.080 2.570 10.480 2.760 ;
        RECT  9.920 0.500 10.230 0.720 ;
        RECT  9.920 2.570 10.080 2.850 ;
        END
        ANTENNADIFFAREA 1.772 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 2.440 0.760 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.610 3.120 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.820 6.320 2.360 ;
        RECT  5.910 1.820 6.080 1.980 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.700 -0.280 11.200 0.280 ;
        RECT  10.420 -0.280 10.700 0.340 ;
        RECT  9.700 -0.280 10.420 0.280 ;
        RECT  9.420 -0.280 9.700 0.340 ;
        RECT  8.030 -0.280 9.420 0.280 ;
        RECT  7.750 -0.280 8.030 1.050 ;
        RECT  6.400 -0.280 7.750 0.280 ;
        RECT  5.680 -0.280 6.400 0.650 ;
        RECT  2.320 -0.280 5.680 0.280 ;
        RECT  2.160 -0.280 2.320 0.740 ;
        RECT  0.880 -0.280 2.160 0.280 ;
        RECT  0.600 -0.280 0.880 0.340 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.700 3.320 11.200 3.880 ;
        RECT  10.420 3.260 10.700 3.880 ;
        RECT  9.600 3.320 10.420 3.880 ;
        RECT  9.440 2.930 9.600 3.880 ;
        RECT  7.930 3.320 9.440 3.880 ;
        RECT  7.250 3.260 7.930 3.880 ;
        RECT  6.380 3.320 7.250 3.880 ;
        RECT  5.780 3.260 6.380 3.880 ;
        RECT  1.840 3.320 5.780 3.880 ;
        RECT  1.680 2.860 1.840 3.880 ;
        RECT  0.880 3.320 1.680 3.880 ;
        RECT  0.600 2.920 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.240 1.430 10.370 1.720 ;
        RECT  10.220 1.070 10.240 1.720 ;
        RECT  10.060 1.070 10.220 2.330 ;
        RECT  9.960 1.070 10.060 1.290 ;
        RECT  9.900 2.010 10.060 2.330 ;
        RECT  9.120 2.010 9.900 2.170 ;
        RECT  9.720 1.570 9.880 1.850 ;
        RECT  8.860 1.690 9.720 1.850 ;
        RECT  8.810 0.480 9.160 0.670 ;
        RECT  8.960 2.010 9.120 3.100 ;
        RECT  4.240 2.940 8.960 3.100 ;
        RECT  8.800 0.830 8.860 1.850 ;
        RECT  8.460 0.510 8.810 0.670 ;
        RECT  8.700 0.830 8.800 2.670 ;
        RECT  8.640 1.690 8.700 2.670 ;
        RECT  8.600 2.340 8.640 2.670 ;
        RECT  8.440 0.510 8.460 1.830 ;
        RECT  8.300 0.510 8.440 2.680 ;
        RECT  8.280 1.550 8.300 2.680 ;
        RECT  5.920 2.520 8.280 2.680 ;
        RECT  7.960 1.290 8.120 2.170 ;
        RECT  7.490 1.290 7.960 1.450 ;
        RECT  7.530 2.010 7.960 2.170 ;
        RECT  7.070 1.660 7.800 1.820 ;
        RECT  7.250 2.010 7.530 2.230 ;
        RECT  7.330 0.560 7.490 1.450 ;
        RECT  6.990 0.560 7.330 0.720 ;
        RECT  6.910 0.960 7.070 1.820 ;
        RECT  6.830 0.440 6.990 0.720 ;
        RECT  6.840 1.500 6.910 1.820 ;
        RECT  6.680 1.500 6.840 2.310 ;
        RECT  6.670 1.080 6.730 1.340 ;
        RECT  5.660 1.500 6.680 1.660 ;
        RECT  6.450 0.810 6.670 1.340 ;
        RECT  5.020 0.810 6.450 0.970 ;
        RECT  5.340 1.160 5.960 1.320 ;
        RECT  5.760 2.170 5.920 2.680 ;
        RECT  5.340 2.220 5.760 2.380 ;
        RECT  5.500 1.500 5.660 1.810 ;
        RECT  5.180 1.160 5.340 2.380 ;
        RECT  5.050 1.380 5.180 2.380 ;
        RECT  4.860 2.620 5.100 2.780 ;
        RECT  4.690 1.380 5.050 1.660 ;
        RECT  4.860 0.810 5.020 1.090 ;
        RECT  4.440 0.930 4.860 1.090 ;
        RECT  4.700 1.820 4.860 2.780 ;
        RECT  4.440 1.820 4.700 1.980 ;
        RECT  4.340 0.460 4.630 0.740 ;
        RECT  2.500 2.440 4.540 2.600 ;
        RECT  4.280 0.930 4.440 1.980 ;
        RECT  2.920 0.460 4.340 0.620 ;
        RECT  4.080 2.760 4.240 3.100 ;
        RECT  3.440 1.300 3.910 1.580 ;
        RECT  2.000 0.910 3.740 1.070 ;
        RECT  2.160 2.760 3.660 2.920 ;
        RECT  3.440 2.110 3.560 2.270 ;
        RECT  3.280 1.230 3.440 2.270 ;
        RECT  1.680 1.230 3.280 1.390 ;
        RECT  2.760 0.460 2.920 0.740 ;
        RECT  2.480 1.870 2.640 2.280 ;
        RECT  1.680 2.120 2.480 2.280 ;
        RECT  2.000 2.540 2.160 2.920 ;
        RECT  1.840 0.490 2.000 1.070 ;
        RECT  1.340 2.540 2.000 2.700 ;
        RECT  1.340 0.490 1.840 0.650 ;
        RECT  1.520 0.810 1.680 1.390 ;
        RECT  1.520 1.550 1.680 2.280 ;
        RECT  0.340 0.810 1.520 0.970 ;
        RECT  1.320 1.950 1.520 2.280 ;
        RECT  1.060 2.540 1.340 2.790 ;
        RECT  0.680 1.130 1.320 1.290 ;
        RECT  0.680 2.120 1.320 2.280 ;
        RECT  0.520 1.130 0.680 2.280 ;
        RECT  0.180 0.520 0.340 2.230 ;
    END
END SEDFFX1TR

MACRO SDFFTRXLTR
    CLASS CORE ;
    FOREIGN SDFFTRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.940 2.760 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.640 0.720 2.020 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.120 1.780 ;
        RECT  2.600 1.240 2.840 1.400 ;
        RECT  2.440 0.440 2.600 1.400 ;
        RECT  0.890 0.440 2.440 0.600 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.030 1.010 10.320 2.360 ;
        END
        ANTENNADIFFAREA 1.128 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.840 1.010 9.120 2.250 ;
        END
        ANTENNADIFFAREA 1.128 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 2.360 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 3.920 1.640 ;
        RECT  3.600 1.240 3.760 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.750 -0.280 10.400 0.280 ;
        RECT  9.400 -0.280 9.750 0.400 ;
        RECT  8.100 -0.280 9.400 0.280 ;
        RECT  7.820 -0.280 8.100 0.670 ;
        RECT  6.440 -0.280 7.820 0.280 ;
        RECT  6.100 -0.280 6.440 0.400 ;
        RECT  4.040 -0.280 6.100 0.280 ;
        RECT  3.760 -0.280 4.040 0.760 ;
        RECT  3.040 -0.280 3.760 0.280 ;
        RECT  2.760 -0.280 3.040 0.800 ;
        RECT  0.730 -0.280 2.760 0.280 ;
        RECT  0.730 0.780 0.930 1.060 ;
        RECT  0.530 -0.280 0.730 1.060 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.750 3.320 10.400 3.880 ;
        RECT  9.400 3.230 9.750 3.880 ;
        RECT  8.100 3.320 9.400 3.880 ;
        RECT  7.820 2.850 8.100 3.880 ;
        RECT  6.260 3.320 7.820 3.880 ;
        RECT  5.980 2.290 6.260 3.880 ;
        RECT  4.080 3.320 5.980 3.880 ;
        RECT  3.800 2.670 4.080 3.880 ;
        RECT  2.640 3.260 3.800 3.880 ;
        RECT  2.360 2.840 2.640 3.880 ;
        RECT  0.960 3.320 2.360 3.880 ;
        RECT  0.680 2.610 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.590 0.570 9.870 3.010 ;
        RECT  8.980 0.570 9.590 0.730 ;
        RECT  8.620 2.850 9.590 3.010 ;
        RECT  8.700 0.450 8.980 0.730 ;
        RECT  8.660 1.400 8.680 1.680 ;
        RECT  8.460 1.000 8.660 2.190 ;
        RECT  8.340 2.850 8.620 3.130 ;
        RECT  8.380 1.000 8.460 1.280 ;
        RECT  8.380 1.910 8.460 2.190 ;
        RECT  7.860 1.910 8.380 2.070 ;
        RECT  8.020 1.440 8.300 1.720 ;
        RECT  7.340 1.440 8.020 1.600 ;
        RECT  7.580 1.910 7.860 2.190 ;
        RECT  7.340 0.440 7.460 0.670 ;
        RECT  7.220 0.440 7.340 2.450 ;
        RECT  7.180 0.440 7.220 2.570 ;
        RECT  6.940 2.290 7.180 2.570 ;
        RECT  6.740 0.520 7.020 0.800 ;
        RECT  6.740 1.360 7.020 1.660 ;
        RECT  5.940 0.640 6.740 0.800 ;
        RECT  6.580 1.500 6.740 1.660 ;
        RECT  6.580 2.290 6.740 2.570 ;
        RECT  6.420 1.500 6.580 2.570 ;
        RECT  5.940 1.500 6.420 1.660 ;
        RECT  5.980 1.820 6.260 2.100 ;
        RECT  5.500 1.820 5.980 1.980 ;
        RECT  5.780 0.440 5.940 0.800 ;
        RECT  5.660 1.380 5.940 1.660 ;
        RECT  4.680 0.440 5.780 0.600 ;
        RECT  5.500 0.760 5.620 1.040 ;
        RECT  5.340 0.760 5.500 2.770 ;
        RECT  5.300 2.610 5.340 2.770 ;
        RECT  5.020 2.610 5.300 2.870 ;
        RECT  5.000 0.760 5.060 1.040 ;
        RECT  4.840 0.760 5.000 2.450 ;
        RECT  4.780 2.290 4.840 2.450 ;
        RECT  4.500 2.290 4.780 2.650 ;
        RECT  4.520 0.440 4.680 2.130 ;
        RECT  4.460 0.480 4.520 2.130 ;
        RECT  3.520 2.290 4.500 2.450 ;
        RECT  4.320 0.480 4.460 0.760 ;
        RECT  4.360 1.910 4.460 2.130 ;
        RECT  4.080 0.920 4.300 1.310 ;
        RECT  3.480 0.920 4.080 1.080 ;
        RECT  3.440 1.910 3.640 2.130 ;
        RECT  3.360 2.290 3.520 2.890 ;
        RECT  3.440 0.500 3.480 1.080 ;
        RECT  3.280 0.500 3.440 2.130 ;
        RECT  3.240 2.520 3.360 2.890 ;
        RECT  3.200 0.500 3.280 0.780 ;
        RECT  2.280 2.520 3.240 2.680 ;
        RECT  2.130 0.880 2.280 2.680 ;
        RECT  2.120 0.760 2.130 2.680 ;
        RECT  1.850 0.760 2.120 1.040 ;
        RECT  1.760 2.520 2.120 2.680 ;
        RECT  1.680 1.200 1.960 2.360 ;
        RECT  1.480 2.520 1.760 2.810 ;
        RECT  1.570 1.200 1.680 1.480 ;
        RECT  0.250 1.320 1.570 1.480 ;
        RECT  0.250 2.530 0.400 2.810 ;
        RECT  0.250 0.790 0.370 1.070 ;
        RECT  0.090 0.790 0.250 2.810 ;
    END
END SDFFTRXLTR

MACRO SDFFTRX4TR
    CLASS CORE ;
    FOREIGN SDFFTRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.940 2.760 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.640 0.720 2.020 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.120 1.780 ;
        RECT  2.600 1.240 2.840 1.400 ;
        RECT  2.440 0.440 2.600 1.400 ;
        RECT  0.890 0.440 2.440 0.600 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.480 0.600 10.720 3.140 ;
        RECT  10.410 0.600 10.480 1.280 ;
        RECT  10.410 2.060 10.480 3.140 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.680 1.090 9.920 2.420 ;
        RECT  9.390 1.090 9.680 1.310 ;
        RECT  9.390 2.140 9.680 2.420 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 2.360 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 3.920 1.640 ;
        RECT  3.600 1.240 3.760 1.560 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 -0.280 11.200 0.280 ;
        RECT  10.880 -0.280 11.110 1.220 ;
        RECT  10.150 -0.280 10.880 0.280 ;
        RECT  9.870 -0.280 10.150 0.610 ;
        RECT  9.190 -0.280 9.870 0.280 ;
        RECT  8.910 -0.280 9.190 0.610 ;
        RECT  8.100 -0.280 8.910 0.280 ;
        RECT  7.820 -0.280 8.100 0.670 ;
        RECT  6.440 -0.280 7.820 0.280 ;
        RECT  6.100 -0.280 6.440 0.400 ;
        RECT  4.040 -0.280 6.100 0.280 ;
        RECT  3.760 -0.280 4.040 0.760 ;
        RECT  3.040 -0.280 3.760 0.280 ;
        RECT  2.760 -0.280 3.040 0.800 ;
        RECT  0.730 -0.280 2.760 0.280 ;
        RECT  0.730 0.780 0.930 1.060 ;
        RECT  0.530 -0.280 0.730 1.060 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 3.320 11.200 3.880 ;
        RECT  10.880 2.060 11.110 3.880 ;
        RECT  10.150 3.320 10.880 3.880 ;
        RECT  9.870 2.910 10.150 3.880 ;
        RECT  9.190 3.320 9.870 3.880 ;
        RECT  8.910 2.910 9.190 3.880 ;
        RECT  7.890 3.320 8.910 3.880 ;
        RECT  7.610 2.500 7.890 3.880 ;
        RECT  6.040 3.320 7.610 3.880 ;
        RECT  5.760 2.290 6.040 3.880 ;
        RECT  4.080 3.320 5.760 3.880 ;
        RECT  3.800 2.670 4.080 3.880 ;
        RECT  2.640 3.260 3.800 3.880 ;
        RECT  2.360 2.840 2.640 3.880 ;
        RECT  0.960 3.320 2.360 3.880 ;
        RECT  0.680 2.610 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.250 1.440 10.320 1.720 ;
        RECT  10.080 0.770 10.250 2.740 ;
        RECT  8.670 0.770 10.080 0.930 ;
        RECT  8.710 2.580 10.080 2.740 ;
        RECT  8.660 1.660 9.520 1.940 ;
        RECT  8.550 2.580 8.710 3.150 ;
        RECT  8.390 0.450 8.670 0.930 ;
        RECT  8.460 1.090 8.660 2.060 ;
        RECT  8.430 2.930 8.550 3.150 ;
        RECT  8.380 1.090 8.460 1.280 ;
        RECT  8.370 1.840 8.460 2.060 ;
        RECT  8.090 1.840 8.370 2.710 ;
        RECT  7.980 1.440 8.260 1.680 ;
        RECT  7.720 1.840 8.090 2.040 ;
        RECT  7.340 1.440 7.980 1.600 ;
        RECT  7.500 1.760 7.720 2.040 ;
        RECT  7.340 0.440 7.460 0.670 ;
        RECT  7.180 0.440 7.340 2.660 ;
        RECT  7.070 2.500 7.180 2.660 ;
        RECT  6.790 2.500 7.070 2.780 ;
        RECT  6.740 0.500 7.020 0.800 ;
        RECT  6.740 1.360 7.020 1.660 ;
        RECT  5.940 0.640 6.740 0.800 ;
        RECT  6.520 1.500 6.740 1.660 ;
        RECT  6.360 1.500 6.520 2.570 ;
        RECT  5.840 1.500 6.360 1.660 ;
        RECT  6.240 2.290 6.360 2.570 ;
        RECT  5.880 1.820 6.160 2.100 ;
        RECT  5.780 0.440 5.940 0.800 ;
        RECT  5.320 1.820 5.880 1.980 ;
        RECT  5.560 1.380 5.840 1.660 ;
        RECT  4.680 0.440 5.780 0.600 ;
        RECT  5.320 0.760 5.620 1.040 ;
        RECT  5.200 0.760 5.320 2.770 ;
        RECT  5.160 0.760 5.200 2.870 ;
        RECT  4.920 2.610 5.160 2.870 ;
        RECT  4.840 0.760 5.000 2.450 ;
        RECT  4.640 2.290 4.840 2.450 ;
        RECT  4.520 0.440 4.680 2.130 ;
        RECT  4.360 2.290 4.640 2.650 ;
        RECT  4.460 0.480 4.520 2.130 ;
        RECT  4.320 0.480 4.460 0.760 ;
        RECT  4.360 1.910 4.460 2.130 ;
        RECT  3.520 2.290 4.360 2.450 ;
        RECT  4.080 0.920 4.300 1.310 ;
        RECT  3.480 0.920 4.080 1.080 ;
        RECT  3.440 1.910 3.640 2.130 ;
        RECT  3.360 2.290 3.520 2.890 ;
        RECT  3.440 0.500 3.480 1.080 ;
        RECT  3.280 0.500 3.440 2.130 ;
        RECT  3.240 2.520 3.360 2.890 ;
        RECT  3.200 0.500 3.280 0.780 ;
        RECT  2.280 2.520 3.240 2.680 ;
        RECT  2.130 0.880 2.280 2.680 ;
        RECT  2.120 0.760 2.130 2.680 ;
        RECT  1.850 0.760 2.120 1.040 ;
        RECT  1.760 2.520 2.120 2.680 ;
        RECT  1.680 1.200 1.960 2.360 ;
        RECT  1.480 2.520 1.760 2.810 ;
        RECT  1.570 1.200 1.680 1.480 ;
        RECT  0.250 1.320 1.570 1.480 ;
        RECT  0.250 2.530 0.400 2.810 ;
        RECT  0.250 0.790 0.370 1.070 ;
        RECT  0.090 0.790 0.250 2.810 ;
    END
END SDFFTRX4TR

MACRO SDFFTRX2TR
    CLASS CORE ;
    FOREIGN SDFFTRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.940 2.760 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.640 0.720 2.020 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.120 1.780 ;
        RECT  2.600 1.240 2.840 1.400 ;
        RECT  2.440 0.440 2.600 1.400 ;
        RECT  0.890 0.440 2.440 0.600 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.080 0.600 10.320 3.140 ;
        RECT  10.010 0.600 10.080 1.280 ;
        RECT  10.010 2.060 10.080 3.140 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.090 9.520 2.420 ;
        RECT  9.070 1.090 9.280 1.310 ;
        RECT  9.070 2.140 9.280 2.420 ;
        END
        ANTENNADIFFAREA 3.025 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 2.360 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 3.920 1.640 ;
        RECT  3.600 1.240 3.760 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 -0.280 10.400 0.280 ;
        RECT  9.550 -0.280 9.830 0.610 ;
        RECT  8.100 -0.280 9.550 0.280 ;
        RECT  7.820 -0.280 8.100 0.670 ;
        RECT  6.440 -0.280 7.820 0.280 ;
        RECT  6.100 -0.280 6.440 0.400 ;
        RECT  4.040 -0.280 6.100 0.280 ;
        RECT  3.760 -0.280 4.040 0.760 ;
        RECT  3.040 -0.280 3.760 0.280 ;
        RECT  2.760 -0.280 3.040 0.800 ;
        RECT  0.730 -0.280 2.760 0.280 ;
        RECT  0.730 0.780 0.930 1.060 ;
        RECT  0.530 -0.280 0.730 1.060 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 3.320 10.400 3.880 ;
        RECT  9.550 2.910 9.830 3.880 ;
        RECT  8.490 3.320 9.550 3.880 ;
        RECT  7.630 3.200 8.490 3.880 ;
        RECT  6.040 3.320 7.630 3.880 ;
        RECT  5.760 2.290 6.040 3.880 ;
        RECT  4.080 3.320 5.760 3.880 ;
        RECT  3.800 2.670 4.080 3.880 ;
        RECT  2.640 3.260 3.800 3.880 ;
        RECT  2.360 2.840 2.640 3.880 ;
        RECT  0.960 3.320 2.360 3.880 ;
        RECT  0.680 2.610 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.850 1.440 9.890 1.720 ;
        RECT  9.680 0.770 9.850 2.740 ;
        RECT  8.980 0.770 9.680 0.930 ;
        RECT  9.010 2.580 9.680 2.740 ;
        RECT  8.660 1.500 9.110 1.780 ;
        RECT  8.850 2.580 9.010 3.150 ;
        RECT  8.700 0.450 8.980 0.930 ;
        RECT  8.730 2.930 8.850 3.150 ;
        RECT  8.460 1.090 8.660 2.060 ;
        RECT  8.380 1.090 8.460 1.280 ;
        RECT  8.320 1.840 8.460 2.060 ;
        RECT  8.040 1.840 8.320 2.630 ;
        RECT  7.980 1.440 8.260 1.680 ;
        RECT  7.720 1.840 8.040 2.040 ;
        RECT  7.340 1.440 7.980 1.600 ;
        RECT  7.500 1.760 7.720 2.040 ;
        RECT  7.340 0.440 7.460 0.670 ;
        RECT  7.180 0.440 7.340 2.660 ;
        RECT  7.070 2.500 7.180 2.660 ;
        RECT  6.790 2.500 7.070 2.780 ;
        RECT  6.740 0.500 7.020 0.800 ;
        RECT  6.740 1.360 7.020 1.660 ;
        RECT  5.940 0.640 6.740 0.800 ;
        RECT  6.520 1.500 6.740 1.660 ;
        RECT  6.360 1.500 6.520 2.570 ;
        RECT  5.840 1.500 6.360 1.660 ;
        RECT  6.240 2.290 6.360 2.570 ;
        RECT  5.880 1.820 6.160 2.100 ;
        RECT  5.780 0.440 5.940 0.800 ;
        RECT  5.320 1.820 5.880 1.980 ;
        RECT  5.560 1.380 5.840 1.660 ;
        RECT  4.680 0.440 5.780 0.600 ;
        RECT  5.320 0.760 5.620 1.040 ;
        RECT  5.200 0.760 5.320 2.770 ;
        RECT  5.160 0.760 5.200 2.870 ;
        RECT  4.920 2.610 5.160 2.870 ;
        RECT  4.840 0.760 5.000 2.450 ;
        RECT  4.640 2.290 4.840 2.450 ;
        RECT  4.520 0.440 4.680 2.130 ;
        RECT  4.360 2.290 4.640 2.650 ;
        RECT  4.460 0.480 4.520 2.130 ;
        RECT  4.320 0.480 4.460 0.760 ;
        RECT  4.360 1.910 4.460 2.130 ;
        RECT  3.520 2.290 4.360 2.450 ;
        RECT  4.080 0.920 4.300 1.310 ;
        RECT  3.480 0.920 4.080 1.080 ;
        RECT  3.440 1.910 3.640 2.130 ;
        RECT  3.360 2.290 3.520 2.890 ;
        RECT  3.440 0.500 3.480 1.080 ;
        RECT  3.280 0.500 3.440 2.130 ;
        RECT  3.240 2.520 3.360 2.890 ;
        RECT  3.200 0.500 3.280 0.780 ;
        RECT  2.280 2.520 3.240 2.680 ;
        RECT  2.130 0.880 2.280 2.680 ;
        RECT  2.120 0.760 2.130 2.680 ;
        RECT  1.850 0.760 2.120 1.040 ;
        RECT  1.760 2.520 2.120 2.680 ;
        RECT  1.680 1.200 1.960 2.360 ;
        RECT  1.480 2.520 1.760 2.810 ;
        RECT  1.570 1.200 1.680 1.480 ;
        RECT  0.250 1.320 1.570 1.480 ;
        RECT  0.250 2.530 0.400 2.810 ;
        RECT  0.250 0.790 0.370 1.070 ;
        RECT  0.090 0.790 0.250 2.810 ;
    END
END SDFFTRX2TR

MACRO SDFFTRX1TR
    CLASS CORE ;
    FOREIGN SDFFTRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.940 2.760 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.640 0.720 2.020 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.120 1.780 ;
        RECT  2.600 1.240 2.840 1.400 ;
        RECT  2.440 0.440 2.600 1.400 ;
        RECT  0.890 0.440 2.440 0.600 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.030 1.000 10.320 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.840 1.000 9.160 2.330 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 2.360 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 3.920 1.640 ;
        RECT  3.600 1.240 3.760 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.790 -0.280 10.400 0.280 ;
        RECT  9.360 -0.280 9.790 0.400 ;
        RECT  8.100 -0.280 9.360 0.280 ;
        RECT  7.820 -0.280 8.100 0.670 ;
        RECT  6.440 -0.280 7.820 0.280 ;
        RECT  6.100 -0.280 6.440 0.400 ;
        RECT  4.040 -0.280 6.100 0.280 ;
        RECT  3.760 -0.280 4.040 0.760 ;
        RECT  3.040 -0.280 3.760 0.280 ;
        RECT  2.760 -0.280 3.040 0.800 ;
        RECT  0.730 -0.280 2.760 0.280 ;
        RECT  0.730 0.780 0.930 1.060 ;
        RECT  0.530 -0.280 0.730 1.060 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.790 3.320 10.400 3.880 ;
        RECT  9.360 3.230 9.790 3.880 ;
        RECT  8.100 3.320 9.360 3.880 ;
        RECT  7.820 2.850 8.100 3.880 ;
        RECT  6.260 3.320 7.820 3.880 ;
        RECT  5.980 2.290 6.260 3.880 ;
        RECT  4.080 3.320 5.980 3.880 ;
        RECT  3.800 2.670 4.080 3.880 ;
        RECT  2.640 3.260 3.800 3.880 ;
        RECT  2.360 2.840 2.640 3.880 ;
        RECT  0.960 3.320 2.360 3.880 ;
        RECT  0.680 2.610 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.590 0.570 9.870 3.010 ;
        RECT  8.980 0.570 9.590 0.730 ;
        RECT  9.070 2.850 9.590 3.010 ;
        RECT  8.780 2.850 9.070 3.130 ;
        RECT  8.700 0.450 8.980 0.730 ;
        RECT  8.660 1.400 8.680 1.680 ;
        RECT  8.460 1.000 8.660 2.190 ;
        RECT  8.380 1.000 8.460 1.280 ;
        RECT  8.380 1.910 8.460 2.190 ;
        RECT  7.860 1.910 8.380 2.070 ;
        RECT  8.020 1.440 8.300 1.720 ;
        RECT  7.340 1.440 8.020 1.600 ;
        RECT  7.580 1.910 7.860 2.190 ;
        RECT  7.340 0.440 7.460 0.670 ;
        RECT  7.220 0.440 7.340 2.450 ;
        RECT  7.180 0.440 7.220 2.570 ;
        RECT  6.940 2.290 7.180 2.570 ;
        RECT  6.740 0.520 7.020 0.800 ;
        RECT  6.740 1.360 7.020 1.660 ;
        RECT  5.940 0.640 6.740 0.800 ;
        RECT  6.580 1.500 6.740 1.660 ;
        RECT  6.580 2.290 6.740 2.570 ;
        RECT  6.420 1.500 6.580 2.570 ;
        RECT  5.940 1.500 6.420 1.660 ;
        RECT  5.980 1.820 6.260 2.100 ;
        RECT  5.500 1.820 5.980 1.980 ;
        RECT  5.780 0.440 5.940 0.800 ;
        RECT  5.660 1.380 5.940 1.660 ;
        RECT  4.680 0.440 5.780 0.600 ;
        RECT  5.500 0.760 5.620 1.040 ;
        RECT  5.340 0.760 5.500 2.770 ;
        RECT  5.300 2.610 5.340 2.770 ;
        RECT  5.020 2.610 5.300 2.870 ;
        RECT  5.000 0.760 5.060 1.040 ;
        RECT  4.840 0.760 5.000 2.450 ;
        RECT  4.780 2.290 4.840 2.450 ;
        RECT  4.500 2.290 4.780 2.650 ;
        RECT  4.520 0.440 4.680 2.130 ;
        RECT  4.460 0.480 4.520 2.130 ;
        RECT  3.520 2.290 4.500 2.450 ;
        RECT  4.320 0.480 4.460 0.760 ;
        RECT  4.360 1.910 4.460 2.130 ;
        RECT  4.080 0.920 4.300 1.310 ;
        RECT  3.480 0.920 4.080 1.080 ;
        RECT  3.440 1.910 3.640 2.130 ;
        RECT  3.360 2.290 3.520 2.890 ;
        RECT  3.440 0.500 3.480 1.080 ;
        RECT  3.280 0.500 3.440 2.130 ;
        RECT  3.240 2.520 3.360 2.890 ;
        RECT  3.200 0.500 3.280 0.780 ;
        RECT  2.280 2.520 3.240 2.680 ;
        RECT  2.130 0.880 2.280 2.680 ;
        RECT  2.120 0.760 2.130 2.680 ;
        RECT  1.850 0.760 2.120 1.040 ;
        RECT  1.760 2.520 2.120 2.680 ;
        RECT  1.680 1.200 1.960 2.360 ;
        RECT  1.480 2.520 1.760 2.810 ;
        RECT  1.570 1.200 1.680 1.480 ;
        RECT  0.250 1.320 1.570 1.480 ;
        RECT  0.250 2.530 0.400 2.810 ;
        RECT  0.250 0.790 0.370 1.070 ;
        RECT  0.090 0.790 0.250 2.810 ;
    END
END SDFFTRX1TR

MACRO SDFFSRHQX8TR
    CLASS CORE ;
    FOREIGN SDFFSRHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.120 1.640 7.690 2.040 ;
        END
        ANTENNAGATEAREA 0.2448 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.000 1.200 6.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.360 1.590 5.520 2.520 ;
        RECT  2.760 2.360 5.360 2.520 ;
        RECT  2.600 1.360 2.760 2.520 ;
        RECT  2.480 1.640 2.600 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.730 1.960 14.850 2.180 ;
        RECT  14.570 1.660 14.730 2.180 ;
        RECT  13.520 1.660 14.570 1.820 ;
        RECT  13.280 1.640 13.520 2.060 ;
        RECT  12.770 1.900 13.280 2.060 ;
        END
        ANTENNAGATEAREA 0.3072 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  18.420 0.630 18.730 3.160 ;
        RECT  17.660 1.440 18.420 2.160 ;
        RECT  17.380 0.630 17.660 3.160 ;
        END
        ANTENNADIFFAREA 8.88 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.220 4.220 1.740 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.390 1.770 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.220 -0.280 19.600 0.280 ;
        RECT  18.940 -0.280 19.220 1.130 ;
        RECT  18.180 -0.280 18.940 0.280 ;
        RECT  17.900 -0.280 18.180 1.190 ;
        RECT  17.100 -0.280 17.900 0.280 ;
        RECT  16.820 -0.280 17.100 0.400 ;
        RECT  15.470 -0.280 16.820 0.280 ;
        RECT  15.190 -0.280 15.470 0.400 ;
        RECT  12.240 -0.280 15.190 0.280 ;
        RECT  11.960 -0.280 12.240 0.400 ;
        RECT  10.080 -0.280 11.960 0.280 ;
        RECT  9.800 -0.280 10.080 0.400 ;
        RECT  7.900 -0.280 9.800 0.280 ;
        RECT  7.620 -0.280 7.900 0.400 ;
        RECT  6.520 -0.280 7.620 0.280 ;
        RECT  5.880 -0.280 6.520 0.400 ;
        RECT  4.100 -0.280 5.880 0.280 ;
        RECT  3.460 -0.280 4.100 0.400 ;
        RECT  0.960 -0.280 3.460 0.280 ;
        RECT  0.320 -0.280 0.960 0.400 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.220 3.320 19.600 3.880 ;
        RECT  18.940 2.100 19.220 3.880 ;
        RECT  18.180 3.320 18.940 3.880 ;
        RECT  17.900 2.320 18.180 3.880 ;
        RECT  17.130 3.320 17.900 3.880 ;
        RECT  16.490 2.740 17.130 3.880 ;
        RECT  15.070 3.320 16.490 3.880 ;
        RECT  14.790 3.200 15.070 3.880 ;
        RECT  12.460 3.320 14.790 3.880 ;
        RECT  12.180 3.200 12.460 3.880 ;
        RECT  11.340 3.320 12.180 3.880 ;
        RECT  11.060 3.200 11.340 3.880 ;
        RECT  9.680 3.320 11.060 3.880 ;
        RECT  9.400 2.590 9.680 3.880 ;
        RECT  6.930 3.320 9.400 3.880 ;
        RECT  6.650 3.200 6.930 3.880 ;
        RECT  1.260 3.320 6.650 3.880 ;
        RECT  0.580 3.200 1.260 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  17.130 0.720 17.160 1.770 ;
        RECT  17.000 0.720 17.130 2.580 ;
        RECT  16.100 0.720 17.000 0.880 ;
        RECT  16.970 1.490 17.000 2.580 ;
        RECT  16.820 1.490 16.970 1.770 ;
        RECT  16.190 2.420 16.970 2.580 ;
        RECT  16.420 1.050 16.670 1.330 ;
        RECT  16.420 1.910 16.670 2.190 ;
        RECT  16.260 1.050 16.420 2.190 ;
        RECT  16.070 1.640 16.260 1.920 ;
        RECT  16.030 2.420 16.190 2.880 ;
        RECT  15.820 0.720 16.100 1.000 ;
        RECT  14.130 2.720 16.030 2.880 ;
        RECT  15.810 1.160 15.880 1.440 ;
        RECT  14.150 0.840 15.820 1.000 ;
        RECT  15.690 1.160 15.810 2.240 ;
        RECT  15.650 1.160 15.690 2.560 ;
        RECT  15.600 1.160 15.650 1.440 ;
        RECT  15.530 1.960 15.650 2.560 ;
        RECT  14.370 2.400 15.530 2.560 ;
        RECT  15.210 2.020 15.330 2.180 ;
        RECT  15.050 1.220 15.210 2.180 ;
        RECT  13.430 1.220 15.050 1.380 ;
        RECT  14.210 1.980 14.370 2.560 ;
        RECT  14.090 1.980 14.210 2.380 ;
        RECT  13.630 0.780 14.150 1.060 ;
        RECT  13.850 2.720 14.130 3.000 ;
        RECT  12.560 2.220 14.090 2.380 ;
        RECT  13.430 0.440 14.010 0.600 ;
        RECT  11.080 2.540 13.620 2.700 ;
        RECT  13.270 0.440 13.430 1.380 ;
        RECT  12.780 3.000 13.410 3.160 ;
        RECT  12.560 0.440 13.270 0.600 ;
        RECT  13.000 0.880 13.100 1.680 ;
        RECT  12.940 0.760 13.000 1.680 ;
        RECT  12.720 0.760 12.940 1.040 ;
        RECT  12.560 1.520 12.940 1.680 ;
        RECT  12.620 2.880 12.780 3.160 ;
        RECT  11.160 1.200 12.730 1.360 ;
        RECT  11.480 0.880 12.720 1.040 ;
        RECT  10.900 2.880 12.620 3.040 ;
        RECT  12.400 0.440 12.560 0.720 ;
        RECT  12.400 1.520 12.560 2.380 ;
        RECT  11.800 0.560 12.400 0.720 ;
        RECT  11.640 0.440 11.800 0.720 ;
        RECT  10.400 0.440 11.640 0.600 ;
        RECT  11.320 0.810 11.480 1.040 ;
        RECT  10.720 0.810 11.320 0.970 ;
        RECT  11.080 1.130 11.160 1.360 ;
        RECT  10.920 1.130 11.080 2.700 ;
        RECT  10.880 1.130 10.920 1.360 ;
        RECT  10.800 1.840 10.920 2.000 ;
        RECT  10.740 2.880 10.900 3.160 ;
        RECT  10.060 3.000 10.740 3.160 ;
        RECT  10.560 0.810 10.720 1.100 ;
        RECT  10.520 1.320 10.680 1.650 ;
        RECT  7.300 0.940 10.560 1.100 ;
        RECT  10.460 2.510 10.540 2.820 ;
        RECT  10.460 1.490 10.520 1.650 ;
        RECT  10.300 1.490 10.460 2.820 ;
        RECT  10.240 0.440 10.400 0.720 ;
        RECT  9.340 1.490 10.300 1.650 ;
        RECT  9.510 0.560 10.240 0.720 ;
        RECT  9.900 2.170 10.060 3.160 ;
        RECT  8.960 2.170 9.900 2.330 ;
        RECT  9.230 0.560 9.510 0.780 ;
        RECT  9.180 1.260 9.340 1.650 ;
        RECT  3.910 0.560 9.230 0.720 ;
        RECT  8.010 1.260 9.180 1.420 ;
        RECT  8.800 1.930 8.960 3.160 ;
        RECT  8.540 1.930 8.800 2.090 ;
        RECT  7.260 3.000 8.800 3.160 ;
        RECT  8.010 2.260 8.640 2.420 ;
        RECT  7.620 2.680 8.600 2.840 ;
        RECT  8.380 1.580 8.540 2.090 ;
        RECT  7.850 1.260 8.010 2.420 ;
        RECT  7.460 2.560 7.620 2.840 ;
        RECT  6.960 2.240 7.460 2.400 ;
        RECT  6.640 2.560 7.460 2.720 ;
        RECT  7.020 0.920 7.300 1.200 ;
        RECT  7.100 2.880 7.260 3.160 ;
        RECT  6.160 2.880 7.100 3.040 ;
        RECT  6.960 1.040 7.020 1.200 ;
        RECT  6.800 1.040 6.960 2.400 ;
        RECT  6.480 0.880 6.640 2.720 ;
        RECT  5.000 0.880 6.480 1.040 ;
        RECT  6.000 2.440 6.480 2.720 ;
        RECT  5.840 1.740 6.310 2.020 ;
        RECT  6.000 2.880 6.160 3.160 ;
        RECT  1.720 3.000 6.000 3.160 ;
        RECT  5.680 1.200 5.840 2.840 ;
        RECT  5.040 1.200 5.680 1.360 ;
        RECT  2.240 2.680 5.680 2.840 ;
        RECT  4.720 2.040 5.120 2.200 ;
        RECT  4.880 1.200 5.040 1.590 ;
        RECT  4.560 0.880 4.720 2.200 ;
        RECT  4.430 0.880 4.560 1.040 ;
        RECT  3.300 2.040 4.120 2.200 ;
        RECT  3.750 0.560 3.910 0.920 ;
        RECT  3.300 0.760 3.750 0.920 ;
        RECT  3.140 0.760 3.300 2.200 ;
        RECT  2.900 0.760 3.140 1.020 ;
        RECT  1.640 0.760 2.900 0.920 ;
        RECT  1.320 0.440 2.800 0.600 ;
        RECT  2.080 1.080 2.240 2.840 ;
        RECT  1.800 1.080 2.080 1.240 ;
        RECT  1.640 1.550 1.900 1.830 ;
        RECT  1.560 2.110 1.720 3.160 ;
        RECT  1.480 0.760 1.640 1.830 ;
        RECT  1.440 2.110 1.560 2.390 ;
        RECT  1.260 1.550 1.480 1.830 ;
        RECT  1.090 2.110 1.440 2.270 ;
        RECT  1.160 0.440 1.320 0.800 ;
        RECT  1.160 0.960 1.320 1.330 ;
        RECT  0.740 0.640 1.160 0.800 ;
        RECT  1.090 1.170 1.160 1.330 ;
        RECT  0.930 1.170 1.090 2.270 ;
        RECT  0.580 0.640 0.740 2.950 ;
        RECT  0.100 0.880 0.580 1.040 ;
        RECT  0.100 2.790 0.580 2.950 ;
    END
END SDFFSRHQX8TR

MACRO SDFFSRHQX4TR
    CLASS CORE ;
    FOREIGN SDFFSRHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.120 1.640 7.690 2.040 ;
        END
        ANTENNAGATEAREA 0.2448 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.000 1.200 6.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.360 1.590 5.520 2.520 ;
        RECT  2.760 2.360 5.360 2.520 ;
        RECT  2.600 1.360 2.760 2.520 ;
        RECT  2.480 1.640 2.600 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.730 1.960 14.850 2.180 ;
        RECT  14.570 1.660 14.730 2.180 ;
        RECT  13.520 1.660 14.570 1.820 ;
        RECT  13.280 1.640 13.520 2.060 ;
        RECT  12.770 1.900 13.280 2.060 ;
        END
        ANTENNAGATEAREA 0.3072 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.380 0.630 17.660 3.160 ;
        RECT  17.280 1.440 17.380 2.160 ;
        END
        ANTENNADIFFAREA 4.44 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.220 4.220 1.740 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.390 1.770 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.180 -0.280 18.400 0.280 ;
        RECT  17.900 -0.280 18.180 1.190 ;
        RECT  17.100 -0.280 17.900 0.280 ;
        RECT  16.820 -0.280 17.100 0.400 ;
        RECT  15.470 -0.280 16.820 0.280 ;
        RECT  15.190 -0.280 15.470 0.400 ;
        RECT  12.240 -0.280 15.190 0.280 ;
        RECT  11.960 -0.280 12.240 0.400 ;
        RECT  10.080 -0.280 11.960 0.280 ;
        RECT  9.800 -0.280 10.080 0.400 ;
        RECT  7.900 -0.280 9.800 0.280 ;
        RECT  7.620 -0.280 7.900 0.400 ;
        RECT  6.520 -0.280 7.620 0.280 ;
        RECT  5.880 -0.280 6.520 0.400 ;
        RECT  4.100 -0.280 5.880 0.280 ;
        RECT  3.460 -0.280 4.100 0.400 ;
        RECT  0.960 -0.280 3.460 0.280 ;
        RECT  0.320 -0.280 0.960 0.400 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.180 3.320 18.400 3.880 ;
        RECT  17.900 2.320 18.180 3.880 ;
        RECT  17.130 3.320 17.900 3.880 ;
        RECT  16.490 2.740 17.130 3.880 ;
        RECT  15.070 3.320 16.490 3.880 ;
        RECT  14.790 3.200 15.070 3.880 ;
        RECT  12.460 3.320 14.790 3.880 ;
        RECT  12.180 3.200 12.460 3.880 ;
        RECT  11.340 3.320 12.180 3.880 ;
        RECT  11.060 3.200 11.340 3.880 ;
        RECT  9.680 3.320 11.060 3.880 ;
        RECT  9.400 2.590 9.680 3.880 ;
        RECT  6.930 3.320 9.400 3.880 ;
        RECT  6.650 3.200 6.930 3.880 ;
        RECT  1.260 3.320 6.650 3.880 ;
        RECT  0.580 3.200 1.260 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.820 0.720 16.980 2.580 ;
        RECT  16.100 0.720 16.820 0.880 ;
        RECT  16.190 2.420 16.820 2.580 ;
        RECT  16.420 1.050 16.600 1.330 ;
        RECT  16.420 1.910 16.600 2.190 ;
        RECT  16.260 1.050 16.420 2.190 ;
        RECT  16.070 1.640 16.260 1.920 ;
        RECT  16.030 2.420 16.190 2.880 ;
        RECT  15.820 0.720 16.100 1.000 ;
        RECT  14.130 2.720 16.030 2.880 ;
        RECT  15.810 1.160 15.880 1.440 ;
        RECT  14.150 0.840 15.820 1.000 ;
        RECT  15.690 1.160 15.810 2.240 ;
        RECT  15.650 1.160 15.690 2.560 ;
        RECT  15.600 1.160 15.650 1.440 ;
        RECT  15.530 1.960 15.650 2.560 ;
        RECT  14.370 2.400 15.530 2.560 ;
        RECT  15.210 2.020 15.330 2.180 ;
        RECT  15.050 1.220 15.210 2.180 ;
        RECT  13.430 1.220 15.050 1.380 ;
        RECT  14.210 1.980 14.370 2.560 ;
        RECT  14.090 1.980 14.210 2.380 ;
        RECT  13.630 0.780 14.150 1.060 ;
        RECT  13.850 2.720 14.130 3.000 ;
        RECT  12.560 2.220 14.090 2.380 ;
        RECT  13.430 0.440 14.010 0.600 ;
        RECT  11.080 2.540 13.620 2.700 ;
        RECT  13.270 0.440 13.430 1.380 ;
        RECT  12.780 3.000 13.410 3.160 ;
        RECT  12.560 0.440 13.270 0.600 ;
        RECT  13.000 0.880 13.100 1.680 ;
        RECT  12.940 0.760 13.000 1.680 ;
        RECT  12.720 0.760 12.940 1.040 ;
        RECT  12.560 1.520 12.940 1.680 ;
        RECT  12.620 2.880 12.780 3.160 ;
        RECT  11.160 1.200 12.730 1.360 ;
        RECT  11.480 0.880 12.720 1.040 ;
        RECT  10.900 2.880 12.620 3.040 ;
        RECT  12.400 0.440 12.560 0.720 ;
        RECT  12.400 1.520 12.560 2.380 ;
        RECT  11.800 0.560 12.400 0.720 ;
        RECT  11.640 0.440 11.800 0.720 ;
        RECT  10.400 0.440 11.640 0.600 ;
        RECT  11.320 0.810 11.480 1.040 ;
        RECT  10.720 0.810 11.320 0.970 ;
        RECT  11.080 1.130 11.160 1.360 ;
        RECT  10.920 1.130 11.080 2.700 ;
        RECT  10.880 1.130 10.920 1.360 ;
        RECT  10.800 1.840 10.920 2.000 ;
        RECT  10.740 2.880 10.900 3.160 ;
        RECT  10.060 3.000 10.740 3.160 ;
        RECT  10.560 0.810 10.720 1.100 ;
        RECT  10.520 1.320 10.680 1.650 ;
        RECT  7.300 0.940 10.560 1.100 ;
        RECT  10.460 2.510 10.540 2.820 ;
        RECT  10.460 1.490 10.520 1.650 ;
        RECT  10.300 1.490 10.460 2.820 ;
        RECT  10.240 0.440 10.400 0.720 ;
        RECT  9.340 1.490 10.300 1.650 ;
        RECT  9.510 0.560 10.240 0.720 ;
        RECT  9.900 2.170 10.060 3.160 ;
        RECT  8.960 2.170 9.900 2.330 ;
        RECT  9.230 0.560 9.510 0.780 ;
        RECT  9.180 1.260 9.340 1.650 ;
        RECT  3.910 0.560 9.230 0.720 ;
        RECT  8.010 1.260 9.180 1.420 ;
        RECT  8.800 1.930 8.960 3.160 ;
        RECT  8.540 1.930 8.800 2.090 ;
        RECT  7.260 3.000 8.800 3.160 ;
        RECT  8.010 2.260 8.640 2.420 ;
        RECT  7.620 2.680 8.600 2.840 ;
        RECT  8.380 1.580 8.540 2.090 ;
        RECT  7.850 1.260 8.010 2.420 ;
        RECT  7.460 2.560 7.620 2.840 ;
        RECT  6.960 2.240 7.460 2.400 ;
        RECT  6.640 2.560 7.460 2.720 ;
        RECT  7.020 0.920 7.300 1.200 ;
        RECT  7.100 2.880 7.260 3.160 ;
        RECT  6.160 2.880 7.100 3.040 ;
        RECT  6.960 1.040 7.020 1.200 ;
        RECT  6.800 1.040 6.960 2.400 ;
        RECT  6.480 0.880 6.640 2.720 ;
        RECT  5.000 0.880 6.480 1.040 ;
        RECT  6.000 2.440 6.480 2.720 ;
        RECT  5.840 1.740 6.310 2.020 ;
        RECT  6.000 2.880 6.160 3.160 ;
        RECT  1.720 3.000 6.000 3.160 ;
        RECT  5.680 1.200 5.840 2.840 ;
        RECT  5.040 1.200 5.680 1.360 ;
        RECT  2.240 2.680 5.680 2.840 ;
        RECT  4.720 2.040 5.120 2.200 ;
        RECT  4.880 1.200 5.040 1.590 ;
        RECT  4.560 0.880 4.720 2.200 ;
        RECT  4.430 0.880 4.560 1.040 ;
        RECT  3.300 2.040 4.120 2.200 ;
        RECT  3.750 0.560 3.910 0.920 ;
        RECT  3.300 0.760 3.750 0.920 ;
        RECT  3.140 0.760 3.300 2.200 ;
        RECT  2.900 0.760 3.140 1.020 ;
        RECT  1.640 0.760 2.900 0.920 ;
        RECT  1.320 0.440 2.800 0.600 ;
        RECT  2.080 1.080 2.240 2.840 ;
        RECT  1.800 1.080 2.080 1.240 ;
        RECT  1.640 1.550 1.900 1.830 ;
        RECT  1.560 2.110 1.720 3.160 ;
        RECT  1.480 0.760 1.640 1.830 ;
        RECT  1.440 2.110 1.560 2.390 ;
        RECT  1.260 1.550 1.480 1.830 ;
        RECT  1.090 2.110 1.440 2.270 ;
        RECT  1.160 0.440 1.320 0.800 ;
        RECT  1.160 0.960 1.320 1.330 ;
        RECT  0.740 0.640 1.160 0.800 ;
        RECT  1.090 1.170 1.160 1.330 ;
        RECT  0.930 1.170 1.090 2.270 ;
        RECT  0.580 0.640 0.740 2.950 ;
        RECT  0.100 0.880 0.580 1.040 ;
        RECT  0.100 2.790 0.580 2.950 ;
    END
END SDFFSRHQX4TR

MACRO SDFFSRHQX2TR
    CLASS CORE ;
    FOREIGN SDFFSRHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 1.240 6.720 1.590 ;
        END
        ANTENNAGATEAREA 0.1968 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.290 1.560 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.640 4.320 1.960 ;
        RECT  4.000 1.640 4.160 2.510 ;
        RECT  2.360 2.350 4.000 2.510 ;
        RECT  2.200 2.230 2.360 2.510 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.720 1.790 12.030 2.190 ;
        RECT  11.610 1.790 11.720 1.970 ;
        RECT  11.280 1.640 11.610 1.970 ;
        RECT  10.650 1.640 11.280 1.800 ;
        RECT  10.490 1.520 10.650 1.800 ;
        END
        ANTENNAGATEAREA 0.216 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.720 0.440 14.800 1.310 ;
        RECT  14.590 0.440 14.720 2.790 ;
        RECT  14.480 1.150 14.590 2.790 ;
        END
        ANTENNADIFFAREA 2.804 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.240 3.520 1.620 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.770 1.640 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.340 -0.280 15.200 0.280 ;
        RECT  14.060 -0.280 14.340 0.340 ;
        RECT  12.920 -0.280 14.060 0.280 ;
        RECT  12.640 -0.280 12.920 0.340 ;
        RECT  10.570 -0.280 12.640 0.280 ;
        RECT  10.290 -0.280 10.570 0.290 ;
        RECT  6.770 -0.280 10.290 0.280 ;
        RECT  5.000 -0.280 6.770 0.290 ;
        RECT  3.320 -0.280 5.000 0.280 ;
        RECT  3.040 -0.280 3.320 0.290 ;
        RECT  0.970 -0.280 3.040 0.280 ;
        RECT  0.690 -0.280 0.970 0.340 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.100 3.320 15.200 3.880 ;
        RECT  14.820 3.260 15.100 3.880 ;
        RECT  14.180 3.320 14.820 3.880 ;
        RECT  13.500 3.260 14.180 3.880 ;
        RECT  12.240 3.320 13.500 3.880 ;
        RECT  11.960 3.260 12.240 3.880 ;
        RECT  10.190 3.320 11.960 3.880 ;
        RECT  9.910 3.260 10.190 3.880 ;
        RECT  9.210 3.320 9.910 3.880 ;
        RECT  8.930 3.260 9.210 3.880 ;
        RECT  7.880 3.320 8.930 3.880 ;
        RECT  7.600 3.260 7.880 3.880 ;
        RECT  5.580 3.320 7.600 3.880 ;
        RECT  5.300 3.260 5.580 3.880 ;
        RECT  1.390 3.320 5.300 3.880 ;
        RECT  0.870 3.160 1.390 3.880 ;
        RECT  0.560 2.650 0.870 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  14.100 0.710 14.160 1.840 ;
        RECT  14.000 0.710 14.100 2.950 ;
        RECT  13.420 0.710 14.000 0.870 ;
        RECT  13.940 1.510 14.000 2.950 ;
        RECT  12.520 2.790 13.940 2.950 ;
        RECT  13.660 2.110 13.780 2.270 ;
        RECT  13.660 1.030 13.720 1.310 ;
        RECT  13.560 1.030 13.660 2.270 ;
        RECT  13.500 1.150 13.560 2.270 ;
        RECT  13.260 1.490 13.500 1.650 ;
        RECT  13.260 0.570 13.420 0.870 ;
        RECT  11.610 0.710 13.260 0.870 ;
        RECT  13.080 1.040 13.240 1.200 ;
        RECT  12.920 1.040 13.080 2.510 ;
        RECT  11.170 2.350 12.920 2.510 ;
        RECT  12.520 1.320 12.680 2.190 ;
        RECT  11.290 1.320 12.520 1.480 ;
        RECT  12.360 2.670 12.520 2.950 ;
        RECT  11.120 2.790 12.360 2.950 ;
        RECT  11.450 0.470 11.610 1.160 ;
        RECT  11.130 0.450 11.290 1.480 ;
        RECT  11.010 2.350 11.170 2.570 ;
        RECT  3.200 0.450 11.130 0.610 ;
        RECT  11.010 1.320 11.130 1.480 ;
        RECT  8.480 2.410 11.010 2.570 ;
        RECT  10.810 0.770 10.970 1.050 ;
        RECT  10.690 1.970 10.850 2.250 ;
        RECT  10.330 0.810 10.810 0.970 ;
        RECT  10.420 2.940 10.700 3.160 ;
        RECT  10.330 2.090 10.690 2.250 ;
        RECT  8.440 2.940 10.420 3.100 ;
        RECT  10.170 0.810 10.330 2.250 ;
        RECT  9.450 0.810 10.170 0.970 ;
        RECT  8.640 2.090 10.170 2.250 ;
        RECT  9.990 1.640 10.010 1.920 ;
        RECT  9.830 1.130 9.990 1.930 ;
        RECT  9.290 1.130 9.830 1.290 ;
        RECT  8.480 1.770 9.830 1.930 ;
        RECT  8.240 1.450 9.670 1.610 ;
        RECT  9.130 0.770 9.290 1.290 ;
        RECT  6.030 0.770 9.130 0.930 ;
        RECT  8.320 1.770 8.480 2.570 ;
        RECT  8.160 2.940 8.440 3.160 ;
        RECT  8.160 1.090 8.240 1.610 ;
        RECT  8.000 1.090 8.160 2.780 ;
        RECT  6.660 2.940 8.160 3.100 ;
        RECT  7.960 1.090 8.000 1.250 ;
        RECT  6.980 2.310 8.000 2.470 ;
        RECT  7.040 1.380 7.470 1.540 ;
        RECT  6.880 1.380 7.040 1.910 ;
        RECT  6.820 2.310 6.980 2.590 ;
        RECT  6.660 1.750 6.880 1.910 ;
        RECT  6.500 1.750 6.660 3.160 ;
        RECT  5.900 3.000 6.500 3.160 ;
        RECT  6.060 2.440 6.340 2.840 ;
        RECT  5.610 2.440 6.060 2.720 ;
        RECT  5.870 0.770 6.030 1.980 ;
        RECT  5.740 2.940 5.900 3.160 ;
        RECT  4.800 2.940 5.740 3.100 ;
        RECT  5.450 0.860 5.610 2.720 ;
        RECT  4.040 0.860 5.450 1.020 ;
        RECT  4.640 2.440 5.450 2.720 ;
        RECT  4.720 1.880 5.000 2.280 ;
        RECT  4.640 2.940 4.800 3.150 ;
        RECT  4.560 1.320 4.720 2.280 ;
        RECT  1.710 2.990 4.640 3.150 ;
        RECT  4.160 1.320 4.560 1.480 ;
        RECT  4.480 2.120 4.560 2.280 ;
        RECT  4.320 2.120 4.480 2.830 ;
        RECT  2.030 2.670 4.320 2.830 ;
        RECT  4.000 1.200 4.160 1.480 ;
        RECT  3.680 0.920 3.840 2.190 ;
        RECT  3.560 0.920 3.680 1.080 ;
        RECT  3.480 2.030 3.680 2.190 ;
        RECT  3.040 0.450 3.200 0.930 ;
        RECT  2.740 0.770 3.040 0.930 ;
        RECT  1.290 0.450 2.880 0.610 ;
        RECT  2.680 1.970 2.800 2.130 ;
        RECT  2.680 0.770 2.740 1.070 ;
        RECT  2.520 0.770 2.680 2.130 ;
        RECT  1.670 0.770 2.520 0.930 ;
        RECT  2.030 1.090 2.340 1.250 ;
        RECT  1.870 1.090 2.030 2.830 ;
        RECT  1.550 1.960 1.710 3.150 ;
        RECT  1.510 0.770 1.670 1.800 ;
        RECT  1.130 1.960 1.550 2.120 ;
        RECT  1.290 1.640 1.510 1.800 ;
        RECT  1.190 1.030 1.350 1.310 ;
        RECT  1.130 0.450 1.290 0.660 ;
        RECT  1.130 1.150 1.190 1.310 ;
        RECT  0.320 0.500 1.130 0.660 ;
        RECT  0.970 1.150 1.130 2.120 ;
        RECT  0.320 1.900 0.420 2.260 ;
        RECT  0.120 0.500 0.320 2.260 ;
    END
END SDFFSRHQX2TR

MACRO SDFFSRHQX1TR
    CLASS CORE ;
    FOREIGN SDFFSRHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.320 1.240 6.500 1.520 ;
        RECT  6.080 1.240 6.320 1.560 ;
        RECT  5.980 1.240 6.080 1.520 ;
        END
        ANTENNAGATEAREA 0.1536 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.140 5.120 1.620 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.640 4.320 1.960 ;
        RECT  4.000 1.640 4.160 2.450 ;
        RECT  2.360 2.290 4.000 2.450 ;
        RECT  2.200 2.170 2.360 2.450 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 1.680 12.140 1.840 ;
        RECT  10.310 1.170 10.470 1.840 ;
        RECT  10.080 1.240 10.310 1.840 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.480 0.880 14.720 2.660 ;
        END
        ANTENNADIFFAREA 1.952 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.180 3.520 1.720 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.800 1.640 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.190 -0.280 14.800 0.280 ;
        RECT  13.910 -0.280 14.190 0.340 ;
        RECT  12.730 -0.280 13.910 0.280 ;
        RECT  12.450 -0.280 12.730 0.340 ;
        RECT  10.390 -0.280 12.450 0.280 ;
        RECT  10.110 -0.280 10.390 0.340 ;
        RECT  5.120 -0.280 10.110 0.280 ;
        RECT  4.840 -0.280 5.120 0.340 ;
        RECT  3.320 -0.280 4.840 0.280 ;
        RECT  3.040 -0.280 3.320 0.340 ;
        RECT  0.980 -0.280 3.040 0.280 ;
        RECT  0.700 -0.280 0.980 0.340 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.130 3.320 14.800 3.880 ;
        RECT  13.500 2.680 14.130 3.880 ;
        RECT  12.210 3.320 13.500 3.880 ;
        RECT  11.930 3.260 12.210 3.880 ;
        RECT  9.970 3.320 11.930 3.880 ;
        RECT  8.950 3.260 9.970 3.880 ;
        RECT  7.780 3.320 8.950 3.880 ;
        RECT  7.500 3.260 7.780 3.880 ;
        RECT  5.660 3.320 7.500 3.880 ;
        RECT  5.380 3.260 5.660 3.880 ;
        RECT  1.400 3.320 5.380 3.880 ;
        RECT  0.700 3.260 1.400 3.880 ;
        RECT  0.000 3.320 0.700 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.850 0.560 14.010 2.520 ;
        RECT  13.230 0.560 13.850 0.720 ;
        RECT  12.610 2.360 13.850 2.520 ;
        RECT  13.530 0.880 13.690 2.190 ;
        RECT  13.290 1.280 13.530 1.560 ;
        RECT  13.070 0.440 13.230 0.720 ;
        RECT  11.430 0.560 13.070 0.720 ;
        RECT  12.990 1.620 13.050 1.900 ;
        RECT  12.830 0.880 12.990 2.200 ;
        RECT  11.110 2.040 12.830 2.200 ;
        RECT  12.610 3.000 12.670 3.160 ;
        RECT  12.490 1.150 12.650 1.880 ;
        RECT  12.450 2.360 12.610 3.160 ;
        RECT  11.110 1.150 12.490 1.310 ;
        RECT  11.430 2.360 12.450 2.520 ;
        RECT  12.390 3.000 12.450 3.160 ;
        RECT  11.270 0.560 11.430 0.990 ;
        RECT  11.270 2.360 11.430 2.640 ;
        RECT  11.050 0.500 11.110 1.310 ;
        RECT  10.950 2.040 11.110 2.780 ;
        RECT  10.950 0.440 11.050 1.310 ;
        RECT  8.480 2.940 11.050 3.100 ;
        RECT  10.770 0.440 10.950 0.660 ;
        RECT  9.050 2.620 10.950 2.780 ;
        RECT  10.630 0.840 10.790 1.120 ;
        RECT  10.630 2.000 10.790 2.280 ;
        RECT  8.240 0.500 10.770 0.660 ;
        RECT  9.490 0.840 10.630 1.000 ;
        RECT  9.490 2.120 10.630 2.280 ;
        RECT  9.330 0.840 9.490 2.280 ;
        RECT  8.940 2.120 9.330 2.280 ;
        RECT  9.000 0.820 9.160 1.920 ;
        RECT  8.870 2.560 9.050 2.780 ;
        RECT  8.920 0.820 9.000 1.260 ;
        RECT  8.500 1.760 9.000 1.920 ;
        RECT  8.660 2.080 8.940 2.280 ;
        RECT  7.920 0.820 8.920 0.980 ;
        RECT  8.500 2.560 8.870 2.720 ;
        RECT  8.180 1.440 8.840 1.600 ;
        RECT  8.340 1.760 8.500 2.720 ;
        RECT  8.190 2.880 8.480 3.100 ;
        RECT  8.080 0.440 8.240 0.660 ;
        RECT  6.840 2.880 8.190 3.040 ;
        RECT  8.020 1.440 8.180 2.720 ;
        RECT  5.440 0.440 8.080 0.600 ;
        RECT  7.510 2.000 8.020 2.160 ;
        RECT  7.760 0.760 7.920 0.980 ;
        RECT  5.820 0.760 7.760 0.920 ;
        RECT  7.480 1.080 7.600 1.240 ;
        RECT  7.480 2.000 7.510 2.370 ;
        RECT  7.320 1.080 7.480 2.370 ;
        RECT  6.750 2.190 7.320 2.370 ;
        RECT  6.820 1.080 6.960 1.240 ;
        RECT  6.530 2.880 6.840 3.100 ;
        RECT  6.660 1.080 6.820 2.010 ;
        RECT  6.530 1.800 6.660 2.010 ;
        RECT  6.370 1.800 6.530 3.100 ;
        RECT  4.800 2.940 6.370 3.100 ;
        RECT  5.850 2.450 6.140 2.780 ;
        RECT  5.820 1.700 5.880 1.860 ;
        RECT  5.440 2.450 5.850 2.660 ;
        RECT  5.600 0.760 5.820 1.860 ;
        RECT  5.280 0.440 5.440 0.660 ;
        RECT  5.280 0.820 5.440 2.660 ;
        RECT  3.200 0.500 5.280 0.660 ;
        RECT  4.140 0.820 5.280 0.980 ;
        RECT  4.640 2.440 5.280 2.660 ;
        RECT  4.880 1.890 5.040 2.280 ;
        RECT  4.720 2.120 4.880 2.280 ;
        RECT  4.640 2.940 4.800 3.150 ;
        RECT  4.560 1.260 4.720 2.280 ;
        RECT  1.720 2.990 4.640 3.150 ;
        RECT  4.160 1.260 4.560 1.420 ;
        RECT  4.480 2.120 4.560 2.280 ;
        RECT  4.320 2.120 4.480 2.830 ;
        RECT  2.040 2.670 4.320 2.830 ;
        RECT  4.000 1.140 4.160 1.420 ;
        RECT  3.680 0.820 3.840 2.130 ;
        RECT  3.560 0.820 3.680 0.980 ;
        RECT  3.480 1.970 3.680 2.130 ;
        RECT  3.040 0.500 3.200 0.920 ;
        RECT  2.740 0.760 3.040 0.920 ;
        RECT  1.300 0.440 2.880 0.600 ;
        RECT  2.680 1.970 2.800 2.130 ;
        RECT  2.680 0.760 2.740 1.040 ;
        RECT  2.520 0.760 2.680 2.130 ;
        RECT  1.680 0.760 2.520 0.920 ;
        RECT  2.040 1.090 2.340 1.250 ;
        RECT  1.880 1.090 2.040 2.830 ;
        RECT  1.560 1.960 1.720 3.150 ;
        RECT  1.520 0.760 1.680 1.800 ;
        RECT  1.140 1.960 1.560 2.120 ;
        RECT  1.300 1.640 1.520 1.800 ;
        RECT  1.200 1.030 1.360 1.310 ;
        RECT  1.140 0.440 1.300 0.720 ;
        RECT  1.140 1.150 1.200 1.310 ;
        RECT  0.320 0.560 1.140 0.720 ;
        RECT  0.980 1.150 1.140 2.120 ;
        RECT  0.320 1.870 0.460 2.190 ;
        RECT  0.160 0.560 0.320 2.190 ;
    END
END SDFFSRHQX1TR

MACRO SDFFSRXLTR
    CLASS CORE ;
    FOREIGN SDFFSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 2.400 8.990 2.780 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.510 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.580 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 1.030 11.520 2.530 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.450 2.250 10.510 2.760 ;
        RECT  10.290 1.030 10.450 2.760 ;
        RECT  10.150 1.030 10.290 1.310 ;
        RECT  10.080 2.250 10.290 2.760 ;
        END
        ANTENNADIFFAREA 1.06 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.560 2.390 ;
        RECT  1.030 2.230 1.280 2.390 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.490 4.400 1.650 ;
        RECT  3.680 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.370 -0.280 11.600 0.280 ;
        RECT  9.210 -0.280 9.370 0.670 ;
        RECT  5.660 -0.280 9.210 0.280 ;
        RECT  4.570 -0.280 5.660 0.370 ;
        RECT  2.860 -0.280 4.570 0.280 ;
        RECT  2.640 -0.280 2.860 0.730 ;
        RECT  2.360 -0.280 2.640 0.280 ;
        RECT  1.220 -0.280 2.360 0.430 ;
        RECT  0.240 -0.280 1.220 0.280 ;
        RECT  0.240 1.030 0.370 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.990 3.320 11.600 3.880 ;
        RECT  10.610 3.260 10.990 3.880 ;
        RECT  9.810 3.320 10.610 3.880 ;
        RECT  9.150 2.730 9.810 3.880 ;
        RECT  7.420 3.320 9.150 3.880 ;
        RECT  7.140 3.260 7.420 3.880 ;
        RECT  5.740 3.320 7.140 3.880 ;
        RECT  4.810 3.000 5.740 3.880 ;
        RECT  3.530 3.320 4.810 3.880 ;
        RECT  3.310 2.830 3.530 3.880 ;
        RECT  1.550 3.320 3.310 3.880 ;
        RECT  1.270 3.260 1.550 3.880 ;
        RECT  0.370 3.320 1.270 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.040 1.430 11.120 1.710 ;
        RECT  10.880 0.690 11.040 3.090 ;
        RECT  10.170 0.690 10.880 0.850 ;
        RECT  10.330 2.930 10.880 3.090 ;
        RECT  10.050 2.930 10.330 3.150 ;
        RECT  10.010 0.440 10.170 0.850 ;
        RECT  9.850 1.090 9.970 1.840 ;
        RECT  9.690 1.090 9.850 2.190 ;
        RECT  9.630 1.680 9.690 2.190 ;
        RECT  9.210 1.680 9.630 1.840 ;
        RECT  9.370 1.200 9.530 1.520 ;
        RECT  7.890 1.200 9.370 1.360 ;
        RECT  9.050 1.640 9.210 1.840 ;
        RECT  8.630 1.640 9.050 1.800 ;
        RECT  8.690 0.440 8.850 0.780 ;
        RECT  8.650 1.960 8.810 2.240 ;
        RECT  6.400 0.440 8.690 0.600 ;
        RECT  8.320 2.080 8.650 2.240 ;
        RECT  8.350 1.520 8.630 1.800 ;
        RECT  8.160 2.080 8.320 3.100 ;
        RECT  8.050 0.760 8.210 1.040 ;
        RECT  8.000 1.580 8.190 1.860 ;
        RECT  6.100 2.940 8.160 3.100 ;
        RECT  7.240 0.760 8.050 0.920 ;
        RECT  7.840 1.580 8.000 2.780 ;
        RECT  7.680 1.080 7.890 1.360 ;
        RECT  4.170 2.620 7.840 2.780 ;
        RECT  7.610 1.080 7.680 2.200 ;
        RECT  7.400 1.200 7.610 2.200 ;
        RECT  7.080 0.760 7.240 2.460 ;
        RECT  6.820 1.590 7.080 1.750 ;
        RECT  6.300 2.300 7.080 2.460 ;
        RECT  6.760 0.980 6.920 1.330 ;
        RECT  6.660 1.980 6.900 2.140 ;
        RECT  6.660 1.170 6.760 1.330 ;
        RECT  6.500 1.170 6.660 2.140 ;
        RECT  6.080 1.170 6.500 1.330 ;
        RECT  6.240 0.440 6.400 1.010 ;
        RECT  6.140 1.490 6.300 2.460 ;
        RECT  5.760 1.490 6.140 1.650 ;
        RECT  5.920 0.530 6.080 1.330 ;
        RECT  5.520 1.810 5.980 1.970 ;
        RECT  4.560 0.530 5.920 0.690 ;
        RECT  5.600 0.850 5.760 1.650 ;
        RECT  4.880 0.850 5.600 1.010 ;
        RECT  5.440 1.810 5.520 2.340 ;
        RECT  5.280 1.170 5.440 2.340 ;
        RECT  5.130 1.170 5.280 1.330 ;
        RECT  5.240 2.120 5.280 2.340 ;
        RECT  4.720 0.850 4.880 1.250 ;
        RECT  4.560 1.090 4.720 2.270 ;
        RECT  3.850 3.000 4.650 3.160 ;
        RECT  4.400 0.530 4.560 0.930 ;
        RECT  4.080 1.090 4.560 1.250 ;
        RECT  4.330 1.810 4.560 2.270 ;
        RECT  3.500 0.770 4.400 0.930 ;
        RECT  3.660 1.810 4.330 1.970 ;
        RECT  3.180 0.450 4.240 0.610 ;
        RECT  4.010 2.190 4.170 2.820 ;
        RECT  2.920 2.190 4.010 2.350 ;
        RECT  3.690 2.510 3.850 3.160 ;
        RECT  2.750 2.510 3.690 2.670 ;
        RECT  3.340 0.770 3.500 2.030 ;
        RECT  3.080 1.870 3.340 2.030 ;
        RECT  3.020 0.450 3.180 1.630 ;
        RECT  2.920 1.470 3.020 1.630 ;
        RECT  2.760 1.470 2.920 2.350 ;
        RECT  2.600 0.960 2.860 1.240 ;
        RECT  2.600 2.510 2.750 2.780 ;
        RECT  2.440 0.960 2.600 2.780 ;
        RECT  2.270 0.590 2.280 2.710 ;
        RECT  2.120 0.590 2.270 2.780 ;
        RECT  0.560 0.590 2.120 0.750 ;
        RECT  1.990 2.550 2.120 2.780 ;
        RECT  0.710 2.550 1.990 2.710 ;
        RECT  1.800 0.920 1.960 1.570 ;
        RECT  0.930 0.920 1.800 1.080 ;
        RECT  0.720 0.920 0.930 1.220 ;
        RECT  0.720 2.210 0.770 2.370 ;
        RECT  0.560 0.920 0.720 2.370 ;
        RECT  0.480 2.550 0.710 3.020 ;
        RECT  0.400 0.440 0.560 0.750 ;
        RECT  0.490 2.210 0.560 2.370 ;
    END
END SDFFSRXLTR

MACRO SDFFSRX4TR
    CLASS CORE ;
    FOREIGN SDFFSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 2.440 8.720 2.870 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.510 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.580 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.610 0.630 11.920 3.160 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.570 1.090 10.850 2.380 ;
        RECT  10.480 1.440 10.570 2.380 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.560 2.390 ;
        RECT  1.030 2.230 1.280 2.390 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.490 4.400 1.650 ;
        RECT  3.680 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 -0.280 12.400 0.280 ;
        RECT  12.080 -0.280 12.310 1.270 ;
        RECT  11.350 -0.280 12.080 0.280 ;
        RECT  11.070 -0.280 11.350 0.610 ;
        RECT  10.370 -0.280 11.070 0.280 ;
        RECT  10.090 -0.280 10.370 0.610 ;
        RECT  9.330 -0.280 10.090 0.280 ;
        RECT  9.050 -0.280 9.330 0.400 ;
        RECT  5.660 -0.280 9.050 0.280 ;
        RECT  4.570 -0.280 5.660 0.370 ;
        RECT  2.860 -0.280 4.570 0.280 ;
        RECT  2.640 -0.280 2.860 0.730 ;
        RECT  2.360 -0.280 2.640 0.280 ;
        RECT  1.220 -0.280 2.360 0.430 ;
        RECT  0.240 -0.280 1.220 0.280 ;
        RECT  0.240 1.030 0.370 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 3.320 12.400 3.880 ;
        RECT  12.080 2.100 12.310 3.880 ;
        RECT  11.350 3.320 12.080 3.880 ;
        RECT  11.070 2.970 11.350 3.880 ;
        RECT  10.370 3.320 11.070 3.880 ;
        RECT  10.090 2.970 10.370 3.880 ;
        RECT  9.230 3.320 10.090 3.880 ;
        RECT  8.950 3.200 9.230 3.880 ;
        RECT  7.840 3.320 8.950 3.880 ;
        RECT  7.060 3.260 7.840 3.880 ;
        RECT  5.740 3.320 7.060 3.880 ;
        RECT  4.810 3.000 5.740 3.880 ;
        RECT  3.530 3.320 4.810 3.880 ;
        RECT  3.310 2.830 3.530 3.880 ;
        RECT  1.550 3.320 3.310 3.880 ;
        RECT  1.270 3.260 1.550 3.880 ;
        RECT  0.370 3.320 1.270 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.390 1.430 11.450 1.710 ;
        RECT  11.230 0.770 11.390 2.710 ;
        RECT  9.890 0.770 11.230 0.930 ;
        RECT  9.850 2.550 11.230 2.710 ;
        RECT  9.790 1.580 10.030 1.860 ;
        RECT  9.610 0.530 9.890 0.930 ;
        RECT  9.570 2.550 9.850 3.150 ;
        RECT  9.630 1.110 9.790 2.190 ;
        RECT  9.350 2.030 9.630 2.310 ;
        RECT  9.290 1.300 9.450 1.860 ;
        RECT  9.130 2.030 9.350 2.190 ;
        RECT  7.740 1.300 9.290 1.460 ;
        RECT  8.970 1.620 9.130 2.190 ;
        RECT  8.310 1.620 8.970 1.780 ;
        RECT  8.690 0.440 8.850 1.130 ;
        RECT  6.400 0.440 8.690 0.600 ;
        RECT  8.320 2.020 8.680 2.180 ;
        RECT  8.160 2.020 8.320 3.100 ;
        RECT  7.990 0.760 8.270 1.140 ;
        RECT  6.100 2.940 8.160 3.100 ;
        RECT  7.200 0.760 7.990 0.920 ;
        RECT  7.920 1.640 7.980 1.860 ;
        RECT  7.760 1.640 7.920 2.780 ;
        RECT  7.720 1.640 7.760 1.860 ;
        RECT  4.170 2.620 7.760 2.780 ;
        RECT  7.560 1.080 7.740 1.460 ;
        RECT  7.460 1.080 7.560 2.200 ;
        RECT  7.400 1.300 7.460 2.200 ;
        RECT  7.200 1.610 7.240 2.460 ;
        RECT  7.080 0.760 7.200 2.460 ;
        RECT  7.040 0.760 7.080 1.770 ;
        RECT  6.300 2.300 7.080 2.460 ;
        RECT  6.820 1.610 7.040 1.770 ;
        RECT  6.660 1.980 6.900 2.140 ;
        RECT  6.720 0.900 6.880 1.450 ;
        RECT  6.660 1.290 6.720 1.450 ;
        RECT  6.500 1.290 6.660 2.140 ;
        RECT  6.080 1.290 6.500 1.450 ;
        RECT  6.240 0.440 6.400 1.130 ;
        RECT  6.140 1.680 6.300 2.460 ;
        RECT  5.760 1.680 6.140 1.840 ;
        RECT  5.920 0.530 6.080 1.450 ;
        RECT  5.520 2.000 5.980 2.160 ;
        RECT  4.560 0.530 5.920 0.690 ;
        RECT  5.600 0.850 5.760 1.840 ;
        RECT  4.880 0.850 5.600 1.010 ;
        RECT  5.440 2.000 5.520 2.340 ;
        RECT  5.280 1.170 5.440 2.340 ;
        RECT  5.130 1.170 5.280 1.330 ;
        RECT  5.240 2.120 5.280 2.340 ;
        RECT  4.720 0.850 4.880 1.250 ;
        RECT  4.560 1.090 4.720 2.270 ;
        RECT  3.850 3.000 4.650 3.160 ;
        RECT  4.400 0.530 4.560 0.930 ;
        RECT  4.080 1.090 4.560 1.250 ;
        RECT  4.330 1.810 4.560 2.270 ;
        RECT  3.500 0.770 4.400 0.930 ;
        RECT  3.660 1.810 4.330 1.970 ;
        RECT  3.180 0.450 4.240 0.610 ;
        RECT  4.010 2.190 4.170 2.820 ;
        RECT  2.920 2.190 4.010 2.350 ;
        RECT  3.690 2.510 3.850 3.160 ;
        RECT  2.750 2.510 3.690 2.670 ;
        RECT  3.340 0.770 3.500 2.030 ;
        RECT  3.080 1.870 3.340 2.030 ;
        RECT  3.020 0.450 3.180 1.630 ;
        RECT  2.920 1.470 3.020 1.630 ;
        RECT  2.760 1.470 2.920 2.350 ;
        RECT  2.600 0.960 2.860 1.240 ;
        RECT  2.600 2.510 2.750 2.780 ;
        RECT  2.440 0.960 2.600 2.780 ;
        RECT  2.270 0.590 2.280 2.710 ;
        RECT  2.120 0.590 2.270 2.780 ;
        RECT  0.560 0.590 2.120 0.750 ;
        RECT  1.990 2.550 2.120 2.780 ;
        RECT  0.710 2.550 1.990 2.710 ;
        RECT  1.800 0.920 1.960 1.570 ;
        RECT  0.930 0.920 1.800 1.080 ;
        RECT  0.720 0.920 0.930 1.220 ;
        RECT  0.720 2.210 0.770 2.370 ;
        RECT  0.560 0.920 0.720 2.370 ;
        RECT  0.480 2.550 0.710 3.020 ;
        RECT  0.400 0.440 0.560 0.750 ;
        RECT  0.490 2.210 0.560 2.370 ;
    END
END SDFFSRX4TR

MACRO SDFFSRX2TR
    CLASS CORE ;
    FOREIGN SDFFSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 2.400 8.990 2.780 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.510 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.580 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 0.590 11.520 3.130 ;
        RECT  11.210 2.100 11.280 3.130 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.170 1.030 10.330 2.760 ;
        RECT  10.080 2.250 10.170 2.760 ;
        END
        ANTENNADIFFAREA 3.478 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.560 2.390 ;
        RECT  1.030 2.230 1.280 2.390 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.490 4.400 1.650 ;
        RECT  3.680 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.090 -0.280 11.600 0.280 ;
        RECT  10.810 -0.280 11.090 1.270 ;
        RECT  9.430 -0.280 10.810 0.280 ;
        RECT  9.150 -0.280 9.430 0.670 ;
        RECT  5.660 -0.280 9.150 0.280 ;
        RECT  4.570 -0.280 5.660 0.370 ;
        RECT  2.860 -0.280 4.570 0.280 ;
        RECT  2.640 -0.280 2.860 0.730 ;
        RECT  2.360 -0.280 2.640 0.280 ;
        RECT  1.220 -0.280 2.360 0.430 ;
        RECT  0.240 -0.280 1.220 0.280 ;
        RECT  0.240 1.030 0.370 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.990 3.320 11.600 3.880 ;
        RECT  10.610 3.260 10.990 3.880 ;
        RECT  9.430 3.320 10.610 3.880 ;
        RECT  9.150 2.730 9.430 3.880 ;
        RECT  7.910 3.320 9.150 3.880 ;
        RECT  7.140 3.260 7.910 3.880 ;
        RECT  5.740 3.320 7.140 3.880 ;
        RECT  4.810 3.000 5.740 3.880 ;
        RECT  3.530 3.320 4.810 3.880 ;
        RECT  3.310 2.830 3.530 3.880 ;
        RECT  1.550 3.320 3.310 3.880 ;
        RECT  1.270 3.260 1.550 3.880 ;
        RECT  0.370 3.320 1.270 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.650 1.430 11.120 1.710 ;
        RECT  10.490 0.690 10.650 3.090 ;
        RECT  10.190 0.690 10.490 0.850 ;
        RECT  9.950 2.930 10.490 3.090 ;
        RECT  9.910 0.440 10.190 0.850 ;
        RECT  9.850 1.030 9.970 1.840 ;
        RECT  9.670 2.930 9.950 3.150 ;
        RECT  9.610 1.030 9.850 2.190 ;
        RECT  9.130 2.030 9.610 2.190 ;
        RECT  9.290 1.200 9.450 1.860 ;
        RECT  7.890 1.200 9.290 1.360 ;
        RECT  8.970 1.640 9.130 2.190 ;
        RECT  8.630 1.640 8.970 1.800 ;
        RECT  8.690 0.440 8.850 0.780 ;
        RECT  8.650 1.960 8.810 2.240 ;
        RECT  6.400 0.440 8.690 0.600 ;
        RECT  8.320 2.080 8.650 2.240 ;
        RECT  8.350 1.520 8.630 1.800 ;
        RECT  8.160 2.080 8.320 3.100 ;
        RECT  8.050 0.760 8.210 1.040 ;
        RECT  8.000 1.580 8.190 1.860 ;
        RECT  6.100 2.940 8.160 3.100 ;
        RECT  7.240 0.760 8.050 0.920 ;
        RECT  7.840 1.580 8.000 2.780 ;
        RECT  7.680 1.080 7.890 1.360 ;
        RECT  4.170 2.620 7.840 2.780 ;
        RECT  7.610 1.080 7.680 2.200 ;
        RECT  7.400 1.200 7.610 2.200 ;
        RECT  7.080 0.760 7.240 2.460 ;
        RECT  6.820 1.590 7.080 1.750 ;
        RECT  6.300 2.300 7.080 2.460 ;
        RECT  6.760 0.980 6.920 1.330 ;
        RECT  6.660 1.980 6.900 2.140 ;
        RECT  6.660 1.170 6.760 1.330 ;
        RECT  6.500 1.170 6.660 2.140 ;
        RECT  6.080 1.170 6.500 1.330 ;
        RECT  6.240 0.440 6.400 1.010 ;
        RECT  6.140 1.490 6.300 2.460 ;
        RECT  5.760 1.490 6.140 1.650 ;
        RECT  5.920 0.530 6.080 1.330 ;
        RECT  5.520 1.810 5.980 1.970 ;
        RECT  4.560 0.530 5.920 0.690 ;
        RECT  5.600 0.850 5.760 1.650 ;
        RECT  4.880 0.850 5.600 1.010 ;
        RECT  5.440 1.810 5.520 2.340 ;
        RECT  5.280 1.170 5.440 2.340 ;
        RECT  5.130 1.170 5.280 1.330 ;
        RECT  5.240 2.120 5.280 2.340 ;
        RECT  4.720 0.850 4.880 1.250 ;
        RECT  4.560 1.090 4.720 2.270 ;
        RECT  3.850 3.000 4.650 3.160 ;
        RECT  4.400 0.530 4.560 0.930 ;
        RECT  4.080 1.090 4.560 1.250 ;
        RECT  4.330 1.810 4.560 2.270 ;
        RECT  3.500 0.770 4.400 0.930 ;
        RECT  3.660 1.810 4.330 1.970 ;
        RECT  3.180 0.450 4.240 0.610 ;
        RECT  4.010 2.190 4.170 2.820 ;
        RECT  2.920 2.190 4.010 2.350 ;
        RECT  3.690 2.510 3.850 3.160 ;
        RECT  2.750 2.510 3.690 2.670 ;
        RECT  3.340 0.770 3.500 2.030 ;
        RECT  3.080 1.870 3.340 2.030 ;
        RECT  3.020 0.450 3.180 1.630 ;
        RECT  2.920 1.470 3.020 1.630 ;
        RECT  2.760 1.470 2.920 2.350 ;
        RECT  2.600 0.960 2.860 1.240 ;
        RECT  2.600 2.510 2.750 2.780 ;
        RECT  2.440 0.960 2.600 2.780 ;
        RECT  2.270 0.590 2.280 2.710 ;
        RECT  2.120 0.590 2.270 2.780 ;
        RECT  0.560 0.590 2.120 0.750 ;
        RECT  1.990 2.550 2.120 2.780 ;
        RECT  0.710 2.550 1.990 2.710 ;
        RECT  1.800 0.920 1.960 1.570 ;
        RECT  0.930 0.920 1.800 1.080 ;
        RECT  0.720 0.920 0.930 1.220 ;
        RECT  0.720 2.210 0.770 2.370 ;
        RECT  0.560 0.920 0.720 2.370 ;
        RECT  0.480 2.550 0.710 3.020 ;
        RECT  0.400 0.440 0.560 0.750 ;
        RECT  0.490 2.210 0.560 2.370 ;
    END
END SDFFSRX2TR

MACRO SDFFSRX1TR
    CLASS CORE ;
    FOREIGN SDFFSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 2.400 8.990 2.780 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.510 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.580 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 1.030 11.520 2.530 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.350 1.030 10.510 2.760 ;
        RECT  10.080 2.250 10.350 2.760 ;
        END
        ANTENNADIFFAREA 1.624 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.560 2.390 ;
        RECT  1.030 2.230 1.280 2.390 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.490 4.400 1.650 ;
        RECT  3.680 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.370 -0.280 11.600 0.280 ;
        RECT  9.210 -0.280 9.370 0.670 ;
        RECT  5.660 -0.280 9.210 0.280 ;
        RECT  4.570 -0.280 5.660 0.370 ;
        RECT  2.860 -0.280 4.570 0.280 ;
        RECT  2.640 -0.280 2.860 0.730 ;
        RECT  2.360 -0.280 2.640 0.280 ;
        RECT  1.220 -0.280 2.360 0.430 ;
        RECT  0.240 -0.280 1.220 0.280 ;
        RECT  0.240 1.030 0.370 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.990 3.320 11.600 3.880 ;
        RECT  10.610 3.260 10.990 3.880 ;
        RECT  9.430 3.320 10.610 3.880 ;
        RECT  9.150 2.730 9.430 3.880 ;
        RECT  7.950 3.320 9.150 3.880 ;
        RECT  7.140 3.260 7.950 3.880 ;
        RECT  5.740 3.320 7.140 3.880 ;
        RECT  4.810 3.000 5.740 3.880 ;
        RECT  3.530 3.320 4.810 3.880 ;
        RECT  3.310 2.830 3.530 3.880 ;
        RECT  1.550 3.320 3.310 3.880 ;
        RECT  1.270 3.260 1.550 3.880 ;
        RECT  0.370 3.320 1.270 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.040 1.430 11.120 1.710 ;
        RECT  10.880 0.690 11.040 3.090 ;
        RECT  10.170 0.690 10.880 0.850 ;
        RECT  9.950 2.930 10.880 3.090 ;
        RECT  10.010 0.440 10.170 0.850 ;
        RECT  9.850 1.090 9.970 1.840 ;
        RECT  9.670 2.930 9.950 3.150 ;
        RECT  9.690 1.090 9.850 2.190 ;
        RECT  9.630 1.680 9.690 2.190 ;
        RECT  9.210 1.680 9.630 1.840 ;
        RECT  9.370 1.200 9.530 1.520 ;
        RECT  7.890 1.200 9.370 1.360 ;
        RECT  9.050 1.640 9.210 1.840 ;
        RECT  8.630 1.640 9.050 1.800 ;
        RECT  8.690 0.440 8.850 0.780 ;
        RECT  8.650 1.960 8.810 2.240 ;
        RECT  6.400 0.440 8.690 0.600 ;
        RECT  8.320 2.080 8.650 2.240 ;
        RECT  8.350 1.520 8.630 1.800 ;
        RECT  8.160 2.080 8.320 3.100 ;
        RECT  8.050 0.760 8.210 1.040 ;
        RECT  8.000 1.580 8.190 1.860 ;
        RECT  6.100 2.940 8.160 3.100 ;
        RECT  7.240 0.760 8.050 0.920 ;
        RECT  7.840 1.580 8.000 2.780 ;
        RECT  7.680 1.080 7.890 1.360 ;
        RECT  4.170 2.620 7.840 2.780 ;
        RECT  7.610 1.080 7.680 2.200 ;
        RECT  7.400 1.200 7.610 2.200 ;
        RECT  7.080 0.760 7.240 2.460 ;
        RECT  6.820 1.590 7.080 1.750 ;
        RECT  6.300 2.300 7.080 2.460 ;
        RECT  6.760 0.980 6.920 1.330 ;
        RECT  6.660 1.980 6.900 2.140 ;
        RECT  6.660 1.170 6.760 1.330 ;
        RECT  6.500 1.170 6.660 2.140 ;
        RECT  6.080 1.170 6.500 1.330 ;
        RECT  6.240 0.440 6.400 1.010 ;
        RECT  6.140 1.490 6.300 2.460 ;
        RECT  5.760 1.490 6.140 1.650 ;
        RECT  5.920 0.530 6.080 1.330 ;
        RECT  5.520 1.810 5.980 1.970 ;
        RECT  4.560 0.530 5.920 0.690 ;
        RECT  5.600 0.850 5.760 1.650 ;
        RECT  4.880 0.850 5.600 1.010 ;
        RECT  5.440 1.810 5.520 2.340 ;
        RECT  5.280 1.170 5.440 2.340 ;
        RECT  5.130 1.170 5.280 1.330 ;
        RECT  5.240 2.120 5.280 2.340 ;
        RECT  4.720 0.850 4.880 1.250 ;
        RECT  4.560 1.090 4.720 2.270 ;
        RECT  3.850 3.000 4.650 3.160 ;
        RECT  4.400 0.530 4.560 0.930 ;
        RECT  4.080 1.090 4.560 1.250 ;
        RECT  4.330 1.810 4.560 2.270 ;
        RECT  3.500 0.770 4.400 0.930 ;
        RECT  3.660 1.810 4.330 1.970 ;
        RECT  3.180 0.450 4.240 0.610 ;
        RECT  4.010 2.190 4.170 2.820 ;
        RECT  2.920 2.190 4.010 2.350 ;
        RECT  3.690 2.510 3.850 3.160 ;
        RECT  2.750 2.510 3.690 2.670 ;
        RECT  3.340 0.770 3.500 2.030 ;
        RECT  3.080 1.870 3.340 2.030 ;
        RECT  3.020 0.450 3.180 1.630 ;
        RECT  2.920 1.470 3.020 1.630 ;
        RECT  2.760 1.470 2.920 2.350 ;
        RECT  2.600 0.960 2.860 1.240 ;
        RECT  2.600 2.510 2.750 2.780 ;
        RECT  2.440 0.960 2.600 2.780 ;
        RECT  2.270 0.590 2.280 2.710 ;
        RECT  2.120 0.590 2.270 2.780 ;
        RECT  0.560 0.590 2.120 0.750 ;
        RECT  1.990 2.550 2.120 2.780 ;
        RECT  0.710 2.550 1.990 2.710 ;
        RECT  1.800 0.920 1.960 1.570 ;
        RECT  0.930 0.920 1.800 1.080 ;
        RECT  0.720 0.920 0.930 1.220 ;
        RECT  0.720 2.210 0.770 2.370 ;
        RECT  0.560 0.920 0.720 2.370 ;
        RECT  0.480 2.550 0.710 3.020 ;
        RECT  0.400 0.440 0.560 0.750 ;
        RECT  0.490 2.210 0.560 2.370 ;
    END
END SDFFSRX1TR

MACRO SDFFSHQX8TR
    CLASS CORE ;
    FOREIGN SDFFSHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.040 1.640 10.570 1.960 ;
        END
        ANTENNAGATEAREA 0.336 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.470 1.580 5.960 1.960 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.240 2.680 1.560 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.540 0.630 17.820 2.990 ;
        RECT  16.860 1.040 17.540 1.760 ;
        RECT  16.580 0.630 16.860 2.990 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.470 3.240 1.750 ;
        RECT  3.020 1.240 3.120 1.750 ;
        RECT  2.840 1.240 3.020 1.630 ;
        END
        ANTENNAGATEAREA 0.2712 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.490 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.4128 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.300 -0.280 18.400 0.280 ;
        RECT  18.020 -0.280 18.300 1.070 ;
        RECT  17.340 -0.280 18.020 0.280 ;
        RECT  17.060 -0.280 17.340 0.670 ;
        RECT  16.340 -0.280 17.060 0.280 ;
        RECT  16.060 -0.280 16.340 0.290 ;
        RECT  14.340 -0.280 16.060 0.280 ;
        RECT  14.780 1.230 15.060 1.510 ;
        RECT  14.340 1.350 14.780 1.510 ;
        RECT  14.060 -0.280 14.340 1.510 ;
        RECT  11.900 -0.280 14.060 0.280 ;
        RECT  11.620 -0.280 11.900 0.640 ;
        RECT  10.860 -0.280 11.620 0.280 ;
        RECT  10.580 -0.280 10.860 0.640 ;
        RECT  9.540 -0.280 10.580 0.280 ;
        RECT  9.260 -0.280 9.540 0.720 ;
        RECT  6.700 -0.280 9.260 0.280 ;
        RECT  6.290 -0.280 6.700 0.400 ;
        RECT  4.990 -0.280 6.290 0.280 ;
        RECT  4.710 -0.280 4.990 0.340 ;
        RECT  2.150 -0.280 4.710 0.280 ;
        RECT  1.010 -0.280 2.150 0.290 ;
        RECT  0.000 -0.280 1.010 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.300 3.320 18.400 3.880 ;
        RECT  18.020 2.130 18.300 3.880 ;
        RECT  17.340 3.320 18.020 3.880 ;
        RECT  17.060 2.130 17.340 3.880 ;
        RECT  16.180 3.320 17.060 3.880 ;
        RECT  15.900 3.200 16.180 3.880 ;
        RECT  14.020 3.320 15.900 3.880 ;
        RECT  13.740 3.200 14.020 3.880 ;
        RECT  11.690 3.320 13.740 3.880 ;
        RECT  11.410 2.890 11.690 3.880 ;
        RECT  10.690 3.320 11.410 3.880 ;
        RECT  10.410 3.200 10.690 3.880 ;
        RECT  9.300 3.260 10.410 3.880 ;
        RECT  8.620 3.200 9.300 3.880 ;
        RECT  7.050 3.320 8.620 3.880 ;
        RECT  6.770 3.200 7.050 3.880 ;
        RECT  6.050 3.320 6.770 3.880 ;
        RECT  5.770 2.930 6.050 3.880 ;
        RECT  3.830 3.260 5.770 3.880 ;
        RECT  3.550 2.930 3.830 3.880 ;
        RECT  3.190 3.320 3.550 3.880 ;
        RECT  2.830 2.930 3.190 3.880 ;
        RECT  1.290 3.320 2.830 3.880 ;
        RECT  0.610 3.200 1.290 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.260 0.450 16.420 3.040 ;
        RECT  15.490 0.450 16.260 0.610 ;
        RECT  15.660 2.880 16.260 3.040 ;
        RECT  15.940 1.580 16.100 2.720 ;
        RECT  15.820 0.890 15.940 1.860 ;
        RECT  15.200 2.560 15.940 2.720 ;
        RECT  15.780 0.770 15.820 1.860 ;
        RECT  15.540 0.770 15.780 1.050 ;
        RECT  15.620 2.110 15.780 2.390 ;
        RECT  15.380 2.880 15.660 3.160 ;
        RECT  15.460 1.230 15.620 2.390 ;
        RECT  15.400 0.440 15.490 0.610 ;
        RECT  15.340 1.230 15.460 1.830 ;
        RECT  14.900 0.440 15.400 0.600 ;
        RECT  14.880 3.000 15.380 3.160 ;
        RECT  14.220 1.670 15.340 1.830 ;
        RECT  15.050 2.560 15.200 2.830 ;
        RECT  14.880 2.600 15.050 2.830 ;
        RECT  14.740 0.440 14.900 0.890 ;
        RECT  13.880 2.670 14.880 2.830 ;
        RECT  14.580 2.110 14.860 2.440 ;
        RECT  14.620 0.610 14.740 0.890 ;
        RECT  13.780 2.110 14.580 2.270 ;
        RECT  13.940 1.670 14.220 1.950 ;
        RECT  13.720 2.430 13.880 2.830 ;
        RECT  13.560 0.450 13.780 2.270 ;
        RECT  13.400 2.430 13.720 2.590 ;
        RECT  12.220 0.450 13.560 0.610 ;
        RECT  13.280 2.750 13.560 3.030 ;
        RECT  13.240 0.800 13.400 2.590 ;
        RECT  12.700 2.750 13.280 2.910 ;
        RECT  13.180 0.800 13.240 2.220 ;
        RECT  12.540 0.800 13.180 0.960 ;
        RECT  13.080 2.060 13.180 2.220 ;
        RECT  12.860 2.060 13.080 2.340 ;
        RECT  12.700 1.120 12.980 1.720 ;
        RECT  12.540 1.560 12.700 2.910 ;
        RECT  12.380 0.800 12.540 1.400 ;
        RECT  12.320 2.060 12.540 2.340 ;
        RECT  12.220 1.120 12.380 1.400 ;
        RECT  12.100 2.570 12.380 3.160 ;
        RECT  11.810 2.060 12.320 2.280 ;
        RECT  12.060 0.450 12.220 0.960 ;
        RECT  10.610 2.570 12.100 2.730 ;
        RECT  10.060 0.800 12.060 0.960 ;
        RECT  11.650 1.170 11.810 2.280 ;
        RECT  11.100 1.170 11.650 1.450 ;
        RECT  11.210 2.120 11.650 2.280 ;
        RECT  11.210 1.680 11.490 1.960 ;
        RECT  10.890 1.680 11.210 1.840 ;
        RECT  10.930 2.120 11.210 2.410 ;
        RECT  9.740 2.120 10.930 2.280 ;
        RECT  10.730 1.200 10.890 1.840 ;
        RECT  9.300 1.200 10.730 1.480 ;
        RECT  10.450 2.570 10.610 2.980 ;
        RECT  10.050 2.820 10.450 2.980 ;
        RECT  10.010 2.440 10.290 2.660 ;
        RECT  9.780 0.760 10.060 1.040 ;
        RECT  9.770 2.820 10.050 3.100 ;
        RECT  9.300 2.440 10.010 2.600 ;
        RECT  6.530 0.880 9.780 1.040 ;
        RECT  7.540 2.820 9.770 2.980 ;
        RECT  9.460 1.810 9.740 2.280 ;
        RECT  9.140 1.200 9.300 2.600 ;
        RECT  7.700 1.200 9.140 1.480 ;
        RECT  7.980 2.440 9.140 2.600 ;
        RECT  8.700 1.920 8.980 2.200 ;
        RECT  7.540 1.920 8.700 2.080 ;
        RECT  7.890 0.440 8.170 0.720 ;
        RECT  7.700 2.320 7.980 2.600 ;
        RECT  5.670 0.560 7.890 0.720 ;
        RECT  7.380 1.640 7.540 2.980 ;
        RECT  7.080 1.640 7.380 1.920 ;
        RECT  2.510 2.610 7.380 2.770 ;
        RECT  6.940 2.140 7.220 2.450 ;
        RECT  6.530 2.290 6.940 2.450 ;
        RECT  6.370 0.880 6.530 2.450 ;
        RECT  6.050 0.880 6.370 1.040 ;
        RECT  2.830 2.290 6.370 2.450 ;
        RECT  5.830 0.880 6.050 1.160 ;
        RECT  5.510 0.560 5.670 1.160 ;
        RECT  5.310 1.000 5.510 1.160 ;
        RECT  5.130 0.440 5.350 0.720 ;
        RECT  5.150 1.000 5.310 2.130 ;
        RECT  4.320 1.000 5.150 1.160 ;
        RECT  4.590 1.910 5.150 2.130 ;
        RECT  4.260 0.560 5.130 0.720 ;
        RECT  3.940 1.470 4.990 1.750 ;
        RECT  3.560 1.910 4.390 2.130 ;
        RECT  4.100 0.880 4.320 1.160 ;
        RECT  4.100 0.450 4.260 0.720 ;
        RECT  0.930 0.450 4.100 0.610 ;
        RECT  3.720 0.770 3.940 1.750 ;
        RECT  2.480 0.770 3.720 0.930 ;
        RECT  3.400 1.090 3.560 2.130 ;
        RECT  3.280 1.090 3.400 1.310 ;
        RECT  2.990 1.910 3.400 2.130 ;
        RECT  2.670 1.840 2.830 2.450 ;
        RECT  2.500 1.840 2.670 2.000 ;
        RECT  2.070 2.930 2.630 3.150 ;
        RECT  2.230 2.160 2.510 2.770 ;
        RECT  2.220 1.720 2.500 2.000 ;
        RECT  2.200 0.770 2.480 1.050 ;
        RECT  1.810 2.160 2.230 2.320 ;
        RECT  1.370 0.770 2.200 0.930 ;
        RECT  1.910 2.480 2.070 3.150 ;
        RECT  1.370 2.480 1.910 2.640 ;
        RECT  1.530 1.090 1.810 2.320 ;
        RECT  1.530 2.800 1.750 3.080 ;
        RECT  0.370 2.800 1.530 2.960 ;
        RECT  1.210 0.770 1.370 2.640 ;
        RECT  0.770 0.450 0.930 2.190 ;
        RECT  0.650 0.770 0.770 2.190 ;
        RECT  0.490 0.770 0.650 1.050 ;
        RECT  0.090 2.680 0.370 2.960 ;
    END
END SDFFSHQX8TR

MACRO SDFFSHQX4TR
    CLASS CORE ;
    FOREIGN SDFFSHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.210 1.630 10.720 1.960 ;
        END
        ANTENNAGATEAREA 0.336 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.870 1.640 6.320 1.970 ;
        RECT  5.650 1.590 5.870 1.970 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.210 2.700 1.560 ;
        RECT  2.080 1.240 2.480 1.560 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.010 1.000 17.120 1.800 ;
        RECT  17.000 1.000 17.010 2.860 ;
        RECT  16.790 0.540 17.000 2.860 ;
        RECT  16.720 0.540 16.790 1.480 ;
        RECT  16.680 0.540 16.720 0.840 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.220 1.470 3.340 1.750 ;
        RECT  3.090 1.240 3.220 1.750 ;
        RECT  2.880 1.240 3.090 1.580 ;
        END
        ANTENNAGATEAREA 0.2712 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.420 2.130 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.4128 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.460 -0.280 17.600 0.280 ;
        RECT  17.180 -0.280 17.460 0.780 ;
        RECT  16.460 -0.280 17.180 0.280 ;
        RECT  16.180 -0.280 16.460 0.340 ;
        RECT  14.470 -0.280 16.180 0.280 ;
        RECT  14.750 1.180 15.030 1.460 ;
        RECT  14.470 1.300 14.750 1.460 ;
        RECT  14.190 -0.280 14.470 1.460 ;
        RECT  12.090 -0.280 14.190 0.280 ;
        RECT  11.810 -0.280 12.090 0.570 ;
        RECT  11.050 -0.280 11.810 0.290 ;
        RECT  10.770 -0.280 11.050 0.570 ;
        RECT  9.690 -0.280 10.770 0.290 ;
        RECT  9.410 -0.280 9.690 0.730 ;
        RECT  6.730 -0.280 9.410 0.290 ;
        RECT  6.450 -0.280 6.730 0.340 ;
        RECT  5.130 -0.280 6.450 0.290 ;
        RECT  4.840 -0.280 5.130 0.370 ;
        RECT  2.100 -0.280 4.840 0.280 ;
        RECT  1.420 -0.280 2.100 0.290 ;
        RECT  0.000 -0.280 1.420 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.510 3.320 17.600 3.880 ;
        RECT  17.230 2.060 17.510 3.880 ;
        RECT  16.450 3.320 17.230 3.880 ;
        RECT  16.170 3.190 16.450 3.880 ;
        RECT  14.220 3.320 16.170 3.880 ;
        RECT  13.940 3.190 14.220 3.880 ;
        RECT  11.830 3.320 13.940 3.880 ;
        RECT  11.550 2.890 11.830 3.880 ;
        RECT  10.830 3.270 11.550 3.880 ;
        RECT  10.550 3.210 10.830 3.880 ;
        RECT  9.470 3.270 10.550 3.880 ;
        RECT  8.770 3.210 9.470 3.880 ;
        RECT  7.210 3.320 8.770 3.880 ;
        RECT  6.930 3.210 7.210 3.880 ;
        RECT  6.210 3.320 6.930 3.880 ;
        RECT  5.930 3.000 6.210 3.880 ;
        RECT  4.010 3.270 5.930 3.880 ;
        RECT  3.730 3.000 4.010 3.880 ;
        RECT  3.260 3.320 3.730 3.880 ;
        RECT  2.980 2.940 3.260 3.880 ;
        RECT  1.290 3.320 2.980 3.880 ;
        RECT  0.630 3.190 1.290 3.880 ;
        RECT  0.000 3.320 0.630 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.350 0.530 16.510 2.980 ;
        RECT  16.020 0.530 16.350 0.690 ;
        RECT  15.830 2.820 16.350 2.980 ;
        RECT  16.060 1.530 16.190 2.660 ;
        RECT  16.030 0.850 16.060 2.660 ;
        RECT  15.900 0.850 16.030 1.810 ;
        RECT  15.410 2.500 16.030 2.660 ;
        RECT  15.860 0.450 16.020 0.690 ;
        RECT  15.700 0.850 15.900 1.010 ;
        RECT  15.580 2.060 15.870 2.340 ;
        RECT  15.030 0.450 15.860 0.610 ;
        RECT  15.610 2.820 15.830 3.160 ;
        RECT  15.420 0.780 15.700 1.010 ;
        RECT  15.150 3.000 15.610 3.160 ;
        RECT  15.420 1.240 15.580 2.340 ;
        RECT  15.310 1.240 15.420 1.780 ;
        RECT  15.250 2.500 15.410 2.760 ;
        RECT  14.330 1.620 15.310 1.780 ;
        RECT  14.140 2.600 15.250 2.760 ;
        RECT  14.830 2.060 15.110 2.390 ;
        RECT  14.870 0.450 15.030 1.000 ;
        RECT  14.750 0.720 14.870 1.000 ;
        RECT  14.010 2.060 14.830 2.220 ;
        RECT  14.170 1.620 14.330 1.900 ;
        RECT  13.980 2.380 14.140 2.760 ;
        RECT  13.850 0.440 14.010 2.220 ;
        RECT  13.630 2.380 13.980 2.540 ;
        RECT  12.410 0.440 13.850 0.600 ;
        RECT  13.480 2.700 13.760 2.980 ;
        RECT  13.470 0.760 13.630 2.540 ;
        RECT  12.840 2.700 13.480 2.860 ;
        RECT  13.410 0.760 13.470 2.460 ;
        RECT  12.830 0.760 13.410 0.920 ;
        RECT  13.000 2.180 13.410 2.460 ;
        RECT  12.990 1.080 13.150 1.860 ;
        RECT  12.840 1.700 12.990 1.860 ;
        RECT  12.680 1.700 12.840 2.860 ;
        RECT  12.670 0.760 12.830 1.360 ;
        RECT  12.520 2.090 12.680 2.350 ;
        RECT  12.450 1.080 12.670 1.360 ;
        RECT  11.950 2.090 12.520 2.290 ;
        RECT  12.240 2.570 12.520 3.030 ;
        RECT  12.250 0.440 12.410 0.920 ;
        RECT  10.210 0.760 12.250 0.920 ;
        RECT  11.210 2.570 12.240 2.730 ;
        RECT  11.790 1.090 11.950 2.290 ;
        RECT  11.290 1.090 11.790 1.370 ;
        RECT  11.350 2.130 11.790 2.290 ;
        RECT  11.350 1.570 11.630 1.850 ;
        RECT  11.050 1.570 11.350 1.730 ;
        RECT  11.070 2.130 11.350 2.410 ;
        RECT  11.050 2.570 11.210 3.010 ;
        RECT  9.890 2.130 11.070 2.290 ;
        RECT  10.890 1.210 11.050 1.730 ;
        RECT  10.190 2.850 11.050 3.010 ;
        RECT  9.450 1.210 10.890 1.450 ;
        RECT  10.150 2.450 10.430 2.690 ;
        RECT  9.930 0.710 10.210 1.050 ;
        RECT  9.910 2.850 10.190 3.110 ;
        RECT  9.450 2.450 10.150 2.610 ;
        RECT  6.750 0.890 9.930 1.050 ;
        RECT  7.690 2.850 9.910 3.010 ;
        RECT  9.610 1.780 9.890 2.290 ;
        RECT  9.290 1.210 9.450 2.610 ;
        RECT  8.250 1.210 9.290 1.490 ;
        RECT  8.130 2.450 9.290 2.610 ;
        RECT  8.850 1.950 9.130 2.230 ;
        RECT  7.750 1.950 8.850 2.110 ;
        RECT  7.850 2.330 8.130 2.610 ;
        RECT  6.890 0.450 7.840 0.730 ;
        RECT  7.690 1.670 7.750 2.110 ;
        RECT  7.530 1.670 7.690 3.010 ;
        RECT  7.130 1.670 7.530 1.830 ;
        RECT  2.610 2.620 7.530 2.780 ;
        RECT  7.150 2.060 7.370 2.460 ;
        RECT  6.750 2.300 7.150 2.460 ;
        RECT  5.770 0.570 6.890 0.730 ;
        RECT  6.590 0.890 6.750 2.460 ;
        RECT  6.210 0.890 6.590 1.050 ;
        RECT  2.930 2.300 6.590 2.460 ;
        RECT  5.930 0.890 6.210 1.170 ;
        RECT  5.610 0.570 5.770 1.170 ;
        RECT  5.490 1.010 5.610 1.170 ;
        RECT  5.330 1.010 5.490 2.140 ;
        RECT  5.290 0.450 5.450 0.730 ;
        RECT  4.420 1.010 5.330 1.170 ;
        RECT  4.770 1.920 5.330 2.140 ;
        RECT  4.300 0.570 5.290 0.730 ;
        RECT  3.980 1.480 5.170 1.760 ;
        RECT  3.660 1.920 4.570 2.140 ;
        RECT  4.140 0.890 4.420 1.170 ;
        RECT  4.140 0.450 4.300 0.730 ;
        RECT  0.830 0.450 4.140 0.610 ;
        RECT  3.820 0.770 3.980 1.760 ;
        RECT  3.220 0.770 3.820 0.930 ;
        RECT  3.500 1.090 3.660 2.140 ;
        RECT  3.380 1.090 3.500 1.310 ;
        RECT  3.120 1.920 3.500 2.140 ;
        RECT  2.120 0.770 3.220 0.990 ;
        RECT  2.770 1.830 2.930 2.460 ;
        RECT  2.170 2.940 2.780 3.100 ;
        RECT  2.610 1.830 2.770 1.990 ;
        RECT  2.310 1.730 2.610 1.990 ;
        RECT  2.330 2.150 2.610 2.780 ;
        RECT  1.770 2.150 2.330 2.310 ;
        RECT  2.010 2.470 2.170 3.100 ;
        RECT  1.200 0.770 2.120 0.930 ;
        RECT  1.310 2.470 2.010 2.630 ;
        RECT  1.630 2.820 1.850 3.130 ;
        RECT  1.640 1.160 1.770 2.310 ;
        RECT  1.610 1.090 1.640 2.310 ;
        RECT  0.370 2.820 1.630 2.980 ;
        RECT  1.360 1.090 1.610 1.320 ;
        RECT  1.200 1.530 1.310 2.630 ;
        RECT  1.150 0.770 1.200 2.630 ;
        RECT  1.040 0.770 1.150 1.690 ;
        RECT  0.830 1.920 0.890 2.200 ;
        RECT  0.670 0.450 0.830 2.200 ;
        RECT  0.260 0.840 0.670 1.060 ;
        RECT  0.090 2.700 0.370 2.980 ;
    END
END SDFFSHQX4TR

MACRO SDFFSHQX2TR
    CLASS CORE ;
    FOREIGN SDFFSHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.260 1.240 8.400 1.560 ;
        RECT  8.040 1.200 8.260 1.560 ;
        END
        ANTENNAGATEAREA 0.2016 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.560 4.760 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.480 1.230 13.520 2.370 ;
        RECT  13.200 0.440 13.480 3.100 ;
        END
        ANTENNADIFFAREA 3.424 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.480 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.24 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.760 -0.280 13.600 0.280 ;
        RECT  10.480 -0.280 10.760 0.980 ;
        RECT  8.600 -0.280 10.480 0.280 ;
        RECT  8.320 -0.280 8.600 0.360 ;
        RECT  8.020 -0.280 8.320 0.280 ;
        RECT  7.740 -0.280 8.020 0.720 ;
        RECT  5.680 -0.280 7.740 0.280 ;
        RECT  5.400 -0.280 5.680 0.360 ;
        RECT  4.620 -0.280 5.400 0.280 ;
        RECT  4.340 -0.280 4.620 0.290 ;
        RECT  0.380 -0.280 4.340 0.280 ;
        RECT  0.100 -0.280 0.380 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.960 3.320 13.600 3.880 ;
        RECT  12.680 3.200 12.960 3.880 ;
        RECT  10.880 3.320 12.680 3.880 ;
        RECT  10.600 2.560 10.880 3.880 ;
        RECT  8.860 3.320 10.600 3.880 ;
        RECT  8.580 2.940 8.860 3.880 ;
        RECT  7.360 3.320 8.580 3.880 ;
        RECT  7.080 3.200 7.360 3.880 ;
        RECT  5.600 3.320 7.080 3.880 ;
        RECT  5.320 2.930 5.600 3.880 ;
        RECT  4.780 3.320 5.320 3.880 ;
        RECT  4.500 3.200 4.780 3.880 ;
        RECT  2.340 3.260 4.500 3.880 ;
        RECT  2.060 2.880 2.340 3.880 ;
        RECT  0.830 3.320 2.060 3.880 ;
        RECT  0.820 3.200 0.830 3.880 ;
        RECT  0.540 2.800 0.820 3.880 ;
        RECT  0.000 3.320 0.540 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.880 0.440 13.040 3.040 ;
        RECT  11.320 0.440 12.880 0.600 ;
        RECT  12.300 2.880 12.880 3.040 ;
        RECT  12.600 1.310 12.720 2.650 ;
        RECT  12.560 0.760 12.600 2.650 ;
        RECT  12.440 0.760 12.560 1.590 ;
        RECT  11.840 2.490 12.560 2.650 ;
        RECT  11.500 0.760 12.440 0.920 ;
        RECT  12.240 1.900 12.400 2.190 ;
        RECT  12.020 2.880 12.300 3.160 ;
        RECT  12.070 1.080 12.240 2.190 ;
        RECT  11.960 1.080 12.070 1.500 ;
        RECT  11.320 3.000 12.020 3.160 ;
        RECT  10.400 1.220 11.960 1.500 ;
        RECT  11.720 2.490 11.840 2.840 ;
        RECT  11.440 1.660 11.720 1.940 ;
        RECT  11.560 2.100 11.720 2.840 ;
        RECT  11.200 2.100 11.560 2.260 ;
        RECT  10.200 1.660 11.440 1.820 ;
        RECT  11.160 0.440 11.320 1.060 ;
        RECT  11.040 2.640 11.320 3.160 ;
        RECT  9.880 1.980 11.200 2.260 ;
        RECT  11.040 0.780 11.160 1.060 ;
        RECT  9.500 2.420 10.420 2.700 ;
        RECT  10.040 0.630 10.200 1.820 ;
        RECT  9.870 2.860 10.150 3.140 ;
        RECT  9.500 0.630 10.040 0.790 ;
        RECT  9.660 0.950 9.880 2.260 ;
        RECT  9.180 2.860 9.870 3.020 ;
        RECT  9.280 0.630 9.500 1.560 ;
        RECT  9.340 2.180 9.500 2.700 ;
        RECT  9.120 2.180 9.340 2.460 ;
        RECT  8.340 0.630 9.280 0.790 ;
        RECT  9.020 2.620 9.180 3.020 ;
        RECT  8.840 0.950 9.120 2.460 ;
        RECT  8.200 2.620 9.020 2.780 ;
        RECT  8.340 2.300 8.840 2.460 ;
        RECT  8.400 1.720 8.680 2.000 ;
        RECT  7.560 1.720 8.400 1.880 ;
        RECT  8.180 0.630 8.340 1.040 ;
        RECT  8.060 2.180 8.340 2.460 ;
        RECT  8.040 2.620 8.200 3.040 ;
        RECT  7.380 0.880 8.180 1.040 ;
        RECT  7.240 2.180 8.060 2.340 ;
        RECT  6.790 2.880 8.040 3.040 ;
        RECT  6.800 2.500 7.880 2.720 ;
        RECT  7.400 1.530 7.560 1.880 ;
        RECT  7.000 1.530 7.400 1.690 ;
        RECT  7.160 0.880 7.380 1.160 ;
        RECT  6.960 1.850 7.240 2.340 ;
        RECT  6.930 0.440 7.210 0.720 ;
        RECT  5.880 0.880 7.160 1.040 ;
        RECT  6.800 1.300 7.000 1.690 ;
        RECT  5.560 0.560 6.930 0.720 ;
        RECT  6.720 1.300 6.800 2.720 ;
        RECT  6.510 2.880 6.790 3.160 ;
        RECT  6.640 1.530 6.720 2.720 ;
        RECT  6.280 2.440 6.640 2.720 ;
        RECT  6.120 2.880 6.510 3.040 ;
        RECT  6.120 1.630 6.320 1.910 ;
        RECT  5.960 1.630 6.120 3.040 ;
        RECT  4.920 2.610 5.960 2.770 ;
        RECT  5.800 0.880 5.880 1.250 ;
        RECT  5.720 0.880 5.800 2.420 ;
        RECT  5.520 1.090 5.720 2.420 ;
        RECT  5.400 0.560 5.560 0.930 ;
        RECT  4.800 1.090 5.520 1.310 ;
        RECT  4.600 2.140 5.520 2.420 ;
        RECT  4.280 0.770 5.400 0.930 ;
        RECT  0.700 0.450 5.240 0.610 ;
        RECT  4.760 2.610 4.920 3.040 ;
        RECT  2.660 2.880 4.760 3.040 ;
        RECT  4.440 2.140 4.600 2.720 ;
        RECT  2.980 2.560 4.440 2.720 ;
        RECT  4.120 0.770 4.280 2.400 ;
        RECT  3.860 1.070 4.120 1.230 ;
        RECT  3.560 2.120 4.120 2.400 ;
        RECT  3.680 1.470 3.960 1.960 ;
        RECT  3.640 0.950 3.860 1.230 ;
        RECT  3.480 1.470 3.680 1.630 ;
        RECT  3.200 0.770 3.480 1.630 ;
        RECT  3.140 1.790 3.360 2.400 ;
        RECT  1.060 0.770 3.200 0.930 ;
        RECT  3.040 1.790 3.140 1.950 ;
        RECT  2.880 1.090 3.040 1.950 ;
        RECT  2.820 2.120 2.980 2.720 ;
        RECT  2.760 1.090 2.880 1.310 ;
        RECT  2.070 2.120 2.820 2.280 ;
        RECT  2.500 2.540 2.660 3.040 ;
        RECT  1.750 2.540 2.500 2.700 ;
        RECT  1.910 1.720 2.070 2.280 ;
        RECT  1.700 1.720 1.910 1.880 ;
        RECT  1.150 2.880 1.840 3.160 ;
        RECT  1.470 2.040 1.750 2.700 ;
        RECT  1.540 1.580 1.700 1.880 ;
        RECT  1.380 2.040 1.470 2.200 ;
        RECT  1.380 1.090 1.460 1.310 ;
        RECT  1.220 1.090 1.380 2.200 ;
        RECT  1.060 2.360 1.150 3.160 ;
        RECT  0.990 0.770 1.060 3.160 ;
        RECT  0.900 0.770 0.990 2.520 ;
        RECT  0.540 0.450 0.700 1.210 ;
        RECT  0.280 0.990 0.540 1.210 ;
        RECT  0.410 2.120 0.500 2.280 ;
        RECT  0.280 2.120 0.410 2.400 ;
        RECT  0.120 0.990 0.280 2.400 ;
        RECT  0.090 0.990 0.120 1.210 ;
    END
END SDFFSHQX2TR

MACRO SDFFSHQX1TR
    CLASS CORE ;
    FOREIGN SDFFSHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.950 8.010 2.360 ;
        RECT  7.540 1.950 7.680 2.170 ;
        END
        ANTENNAGATEAREA 0.1536 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.640 4.810 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.210 2.320 1.570 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.160 2.030 11.280 2.210 ;
        RECT  10.840 0.840 11.160 2.210 ;
        RECT  10.730 0.840 10.840 1.270 ;
        END
        ANTENNADIFFAREA 1.528 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.640 2.810 2.020 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.630 1.970 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.910 -0.280 12.000 0.280 ;
        RECT  10.630 -0.280 10.910 0.610 ;
        RECT  9.850 -0.280 10.630 0.280 ;
        RECT  9.570 -0.280 9.850 0.350 ;
        RECT  8.230 -0.280 9.570 0.280 ;
        RECT  7.960 -0.280 8.230 0.340 ;
        RECT  7.610 -0.280 7.960 0.310 ;
        RECT  7.450 -0.280 7.610 0.670 ;
        RECT  5.350 -0.280 7.450 0.280 ;
        RECT  5.070 -0.280 5.350 0.340 ;
        RECT  4.600 -0.280 5.070 0.310 ;
        RECT  2.700 -0.280 4.600 0.340 ;
        RECT  2.420 -0.280 2.700 0.350 ;
        RECT  0.630 -0.280 2.420 0.290 ;
        RECT  0.350 -0.280 0.630 0.360 ;
        RECT  0.000 -0.280 0.350 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.760 3.320 12.000 3.880 ;
        RECT  10.480 2.970 10.760 3.880 ;
        RECT  7.800 3.320 10.480 3.880 ;
        RECT  7.520 3.010 7.800 3.880 ;
        RECT  7.000 3.320 7.520 3.880 ;
        RECT  6.720 3.210 7.000 3.880 ;
        RECT  5.510 3.320 6.720 3.880 ;
        RECT  5.180 3.270 5.510 3.880 ;
        RECT  4.490 3.320 5.180 3.880 ;
        RECT  4.210 3.210 4.490 3.880 ;
        RECT  2.170 3.270 4.210 3.880 ;
        RECT  1.890 2.830 2.170 3.880 ;
        RECT  0.830 3.320 1.890 3.880 ;
        RECT  0.550 3.060 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.790 0.950 11.850 1.270 ;
        RECT  11.630 0.460 11.790 2.750 ;
        RECT  11.420 0.460 11.630 0.620 ;
        RECT  11.390 2.470 11.630 2.750 ;
        RECT  10.280 2.470 11.390 2.630 ;
        RECT  10.350 0.960 10.510 2.080 ;
        RECT  10.070 0.450 10.350 0.690 ;
        RECT  10.210 0.960 10.350 1.180 ;
        RECT  9.960 1.870 10.350 2.080 ;
        RECT  10.120 2.470 10.280 3.100 ;
        RECT  9.520 1.370 10.190 1.530 ;
        RECT  10.000 2.890 10.120 3.100 ;
        RECT  9.520 0.530 10.070 0.690 ;
        RECT  9.680 1.870 9.960 2.150 ;
        RECT  9.390 0.530 9.520 2.590 ;
        RECT  9.360 0.450 9.390 2.590 ;
        RECT  9.110 0.450 9.360 0.690 ;
        RECT  8.990 2.430 9.360 2.590 ;
        RECT  8.950 1.990 9.200 2.270 ;
        RECT  8.710 2.430 8.990 2.710 ;
        RECT  8.840 0.530 8.950 2.270 ;
        RECT  8.790 0.460 8.840 2.270 ;
        RECT  8.560 0.460 8.790 0.690 ;
        RECT  8.120 2.940 8.790 3.100 ;
        RECT  8.470 0.850 8.630 1.790 ;
        RECT  8.000 0.530 8.560 0.690 ;
        RECT  8.350 0.850 8.470 1.070 ;
        RECT  8.450 1.630 8.470 1.790 ;
        RECT  8.290 1.630 8.450 2.710 ;
        RECT  6.450 1.230 8.310 1.450 ;
        RECT  6.890 1.630 8.290 1.790 ;
        RECT  7.960 2.690 8.120 3.100 ;
        RECT  7.840 0.530 8.000 1.050 ;
        RECT  6.530 2.690 7.960 2.850 ;
        RECT  7.150 0.890 7.840 1.050 ;
        RECT  6.450 2.330 7.520 2.490 ;
        RECT  6.870 0.510 7.150 1.050 ;
        RECT  6.610 1.630 6.890 1.910 ;
        RECT  5.760 0.890 6.870 1.050 ;
        RECT  6.430 0.480 6.710 0.730 ;
        RECT  6.370 2.690 6.530 3.160 ;
        RECT  6.290 1.230 6.450 2.490 ;
        RECT  5.380 0.570 6.430 0.730 ;
        RECT  6.190 2.890 6.370 3.160 ;
        RECT  6.200 2.330 6.290 2.490 ;
        RECT  6.020 2.330 6.200 2.670 ;
        RECT  5.860 2.890 6.190 3.050 ;
        RECT  5.860 1.650 5.990 1.930 ;
        RECT  5.700 1.650 5.860 3.050 ;
        RECT  5.600 0.890 5.760 1.380 ;
        RECT  2.490 2.890 5.700 3.050 ;
        RECT  5.490 1.210 5.600 1.380 ;
        RECT  5.330 1.210 5.490 2.610 ;
        RECT  5.220 0.570 5.380 1.050 ;
        RECT  4.540 1.210 5.330 1.430 ;
        RECT  4.950 2.450 5.330 2.610 ;
        RECT  4.240 0.890 5.220 1.050 ;
        RECT  4.760 0.510 5.040 0.730 ;
        RECT  4.670 2.450 4.950 2.730 ;
        RECT  2.260 0.570 4.760 0.730 ;
        RECT  2.810 2.570 4.670 2.730 ;
        RECT  4.080 0.890 4.240 2.400 ;
        RECT  3.660 0.950 4.080 1.110 ;
        RECT  3.450 2.240 4.080 2.400 ;
        RECT  3.640 1.390 3.920 2.030 ;
        RECT  3.480 1.390 3.640 1.550 ;
        RECT  3.320 0.890 3.480 1.550 ;
        RECT  1.940 0.890 3.320 1.050 ;
        RECT  3.150 1.810 3.250 2.400 ;
        RECT  2.970 1.210 3.150 2.400 ;
        RECT  2.860 1.210 2.970 1.430 ;
        RECT  2.650 2.190 2.810 2.730 ;
        RECT  2.070 2.190 2.650 2.350 ;
        RECT  2.330 2.510 2.490 3.050 ;
        RECT  1.750 2.510 2.330 2.670 ;
        RECT  2.100 0.450 2.260 0.730 ;
        RECT  0.950 0.450 2.100 0.610 ;
        RECT  1.970 1.790 2.070 2.350 ;
        RECT  1.910 1.730 1.970 2.350 ;
        RECT  1.780 0.770 1.940 1.050 ;
        RECT  1.810 1.730 1.910 2.010 ;
        RECT  1.270 0.770 1.780 0.930 ;
        RECT  1.590 2.180 1.750 2.670 ;
        RECT  1.270 2.830 1.610 3.110 ;
        RECT  1.470 1.090 1.590 2.670 ;
        RECT  1.430 1.090 1.470 2.340 ;
        RECT  1.110 0.770 1.270 3.110 ;
        RECT  0.790 0.450 0.950 2.680 ;
        RECT  0.110 0.920 0.790 1.080 ;
        RECT  0.110 2.520 0.790 2.680 ;
    END
END SDFFSHQX1TR

MACRO SDFFSXLTR
    CLASS CORE ;
    FOREIGN SDFFSXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.240 8.080 1.640 ;
        RECT  7.680 1.240 7.740 3.160 ;
        RECT  7.580 1.480 7.680 3.160 ;
        RECT  6.820 2.940 7.580 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.580 1.330 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.580 0.400 1.860 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.080 1.030 10.320 2.360 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.110 1.030 9.270 2.760 ;
        RECT  9.030 1.030 9.110 1.310 ;
        RECT  9.100 2.060 9.110 2.760 ;
        RECT  8.880 2.440 9.100 2.760 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.040 1.920 2.360 ;
        RECT  1.550 1.330 1.710 2.360 ;
        RECT  1.370 2.170 1.550 2.360 ;
        RECT  1.090 2.170 1.370 2.450 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.640 4.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.840 -0.280 10.400 0.280 ;
        RECT  9.560 -0.280 9.840 0.420 ;
        RECT  8.470 -0.280 9.560 0.280 ;
        RECT  8.190 -0.280 8.470 0.760 ;
        RECT  3.950 -0.280 8.190 0.280 ;
        RECT  3.670 -0.280 3.950 0.390 ;
        RECT  1.610 -0.280 3.670 0.340 ;
        RECT  1.330 -0.280 1.610 0.400 ;
        RECT  0.350 -0.280 1.330 0.280 ;
        RECT  0.350 1.030 0.400 1.310 ;
        RECT  0.080 -0.280 0.350 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.890 3.320 10.400 3.880 ;
        RECT  9.570 3.240 9.890 3.880 ;
        RECT  8.220 3.320 9.570 3.880 ;
        RECT  7.940 2.460 8.220 3.880 ;
        RECT  6.660 3.320 7.940 3.880 ;
        RECT  6.440 2.850 6.660 3.880 ;
        RECT  5.000 3.320 6.440 3.880 ;
        RECT  4.720 2.990 5.000 3.880 ;
        RECT  3.950 3.320 4.720 3.880 ;
        RECT  3.670 2.990 3.950 3.880 ;
        RECT  1.610 3.260 3.670 3.880 ;
        RECT  1.330 3.200 1.610 3.880 ;
        RECT  0.090 3.260 1.330 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.670 1.700 9.920 1.980 ;
        RECT  9.510 0.710 9.670 3.080 ;
        RECT  9.140 0.710 9.510 0.870 ;
        RECT  9.320 2.920 9.510 3.080 ;
        RECT  9.040 2.920 9.320 3.160 ;
        RECT  8.860 0.440 9.140 0.870 ;
        RECT  8.870 1.450 8.950 1.730 ;
        RECT  8.710 1.030 8.870 2.190 ;
        RECT  8.560 1.030 8.710 1.310 ;
        RECT  7.900 1.910 8.710 2.190 ;
        RECT  8.400 1.470 8.520 1.750 ;
        RECT  8.240 0.920 8.400 1.750 ;
        RECT  7.420 0.920 8.240 1.080 ;
        RECT  7.580 0.440 7.860 0.760 ;
        RECT  5.080 0.440 7.580 0.600 ;
        RECT  7.260 0.760 7.420 2.780 ;
        RECT  6.720 0.760 7.260 0.920 ;
        RECT  6.940 2.380 7.260 2.780 ;
        RECT  6.880 1.200 7.100 2.220 ;
        RECT  6.720 2.380 6.940 2.540 ;
        RECT  6.680 1.200 6.880 1.360 ;
        RECT  6.440 1.910 6.720 2.540 ;
        RECT  6.280 1.080 6.680 1.360 ;
        RECT  5.540 0.760 6.440 0.920 ;
        RECT  6.120 1.080 6.280 3.160 ;
        RECT  5.700 1.080 6.120 1.300 ;
        RECT  5.560 3.000 6.120 3.160 ;
        RECT  5.740 1.460 5.960 2.590 ;
        RECT  5.540 1.460 5.740 1.620 ;
        RECT  5.280 2.220 5.560 3.160 ;
        RECT  5.380 0.760 5.540 1.620 ;
        RECT  4.600 1.450 5.380 1.610 ;
        RECT  5.110 1.780 5.330 2.060 ;
        RECT  5.160 2.990 5.280 3.160 ;
        RECT  4.950 1.780 5.110 2.830 ;
        RECT  4.920 0.440 5.080 1.290 ;
        RECT  4.510 2.670 4.950 2.830 ;
        RECT  4.800 1.010 4.920 1.290 ;
        RECT  3.190 2.330 4.790 2.490 ;
        RECT  4.440 1.030 4.600 1.610 ;
        RECT  4.440 1.910 4.560 2.130 ;
        RECT  2.750 0.550 4.510 0.830 ;
        RECT  4.230 2.670 4.510 2.890 ;
        RECT  4.280 1.030 4.440 2.130 ;
        RECT  3.830 1.320 4.280 1.480 ;
        RECT  3.430 2.670 4.230 2.830 ;
        RECT  3.550 1.200 3.830 1.480 ;
        RECT  3.150 2.670 3.430 2.900 ;
        RECT  2.910 0.990 3.190 2.490 ;
        RECT  2.750 2.670 3.150 2.830 ;
        RECT  2.590 0.550 2.750 2.830 ;
        RECT  2.270 0.690 2.430 2.780 ;
        RECT  0.730 0.690 2.270 0.850 ;
        RECT  0.730 2.620 2.270 2.780 ;
        RECT  1.890 1.010 2.110 1.500 ;
        RECT  0.990 1.010 1.890 1.170 ;
        RECT  0.720 1.010 0.990 1.310 ;
        RECT  0.720 2.120 0.930 2.400 ;
        RECT  0.510 0.470 0.730 0.850 ;
        RECT  0.480 2.620 0.730 2.990 ;
        RECT  0.560 1.010 0.720 2.400 ;
    END
END SDFFSXLTR

MACRO SDFFSX4TR
    CLASS CORE ;
    FOREIGN SDFFSX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.240 7.920 1.640 ;
        RECT  7.620 1.480 7.680 1.640 ;
        RECT  7.460 1.480 7.620 3.160 ;
        RECT  6.800 2.940 7.460 3.160 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.310 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.880 1.090 11.120 2.210 ;
        RECT  10.750 1.090 10.880 1.250 ;
        RECT  10.750 1.930 10.880 2.210 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 0.770 11.440 2.560 ;
        RECT  9.790 0.770 11.280 0.930 ;
        RECT  10.320 2.400 11.280 2.560 ;
        RECT  10.080 1.840 10.320 2.560 ;
        RECT  10.070 1.930 10.080 2.560 ;
        RECT  9.790 1.930 10.070 3.010 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.040 1.920 2.360 ;
        RECT  1.610 1.300 1.770 2.360 ;
        RECT  1.470 1.300 1.610 1.460 ;
        RECT  1.350 2.170 1.610 2.360 ;
        RECT  1.070 2.170 1.350 2.450 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.640 4.070 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.510 -0.280 11.600 0.280 ;
        RECT  11.230 -0.280 11.510 0.610 ;
        RECT  10.550 -0.280 11.230 0.280 ;
        RECT  10.270 -0.280 10.550 0.610 ;
        RECT  9.820 -0.280 10.270 0.290 ;
        RECT  9.590 -0.280 9.820 0.280 ;
        RECT  9.320 -0.280 9.590 1.220 ;
        RECT  8.270 -0.280 9.320 0.280 ;
        RECT  7.990 -0.280 8.270 0.760 ;
        RECT  3.870 -0.280 7.990 0.280 ;
        RECT  3.590 -0.280 3.870 0.390 ;
        RECT  1.590 -0.280 3.590 0.340 ;
        RECT  1.310 -0.280 1.590 0.400 ;
        RECT  0.330 -0.280 1.310 0.280 ;
        RECT  0.330 1.030 0.390 1.310 ;
        RECT  0.170 -0.280 0.330 1.310 ;
        RECT  0.000 -0.280 0.170 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.510 3.320 11.600 3.880 ;
        RECT  11.230 2.880 11.510 3.880 ;
        RECT  10.550 3.320 11.230 3.880 ;
        RECT  10.270 2.930 10.550 3.880 ;
        RECT  9.590 3.320 10.270 3.880 ;
        RECT  9.310 2.970 9.590 3.880 ;
        RECT  8.080 3.320 9.310 3.880 ;
        RECT  7.800 3.200 8.080 3.880 ;
        RECT  6.640 3.320 7.800 3.880 ;
        RECT  6.420 2.850 6.640 3.880 ;
        RECT  4.980 3.320 6.420 3.880 ;
        RECT  4.700 2.990 4.980 3.880 ;
        RECT  3.930 3.320 4.700 3.880 ;
        RECT  3.650 2.990 3.930 3.880 ;
        RECT  1.470 3.260 3.650 3.880 ;
        RECT  1.190 3.200 1.470 3.880 ;
        RECT  0.370 3.260 1.190 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.250 1.410 10.670 1.660 ;
        RECT  9.110 1.380 9.250 2.780 ;
        RECT  9.090 1.030 9.110 2.780 ;
        RECT  8.830 1.030 9.090 1.660 ;
        RECT  9.030 2.620 9.090 2.780 ;
        RECT  8.750 2.620 9.030 3.130 ;
        RECT  8.670 0.540 8.750 0.820 ;
        RECT  8.510 0.540 8.670 2.460 ;
        RECT  8.470 0.540 8.510 0.820 ;
        RECT  8.030 2.300 8.510 2.460 ;
        RECT  8.240 1.360 8.350 1.640 ;
        RECT  8.080 0.920 8.240 1.640 ;
        RECT  7.300 0.920 8.080 1.080 ;
        RECT  7.780 1.910 8.030 2.460 ;
        RECT  7.460 0.440 7.740 0.760 ;
        RECT  4.910 0.440 7.460 0.600 ;
        RECT  7.140 0.760 7.300 2.780 ;
        RECT  6.700 0.760 7.140 0.920 ;
        RECT  6.920 2.380 7.140 2.780 ;
        RECT  6.820 1.200 6.980 2.220 ;
        RECT  6.580 2.380 6.920 2.540 ;
        RECT  6.660 1.200 6.820 1.360 ;
        RECT  6.260 1.080 6.660 1.360 ;
        RECT  6.420 1.910 6.580 2.540 ;
        RECT  5.290 0.760 6.420 0.920 ;
        RECT  6.100 1.080 6.260 3.160 ;
        RECT  5.590 1.080 6.100 1.300 ;
        RECT  5.540 3.000 6.100 3.160 ;
        RECT  5.720 1.460 5.940 2.590 ;
        RECT  5.290 1.460 5.720 1.620 ;
        RECT  5.320 2.220 5.540 3.160 ;
        RECT  5.140 2.990 5.320 3.160 ;
        RECT  5.160 1.780 5.310 2.060 ;
        RECT  5.130 0.760 5.290 1.620 ;
        RECT  5.000 1.780 5.160 2.830 ;
        RECT  4.390 1.460 5.130 1.620 ;
        RECT  4.510 2.670 5.000 2.830 ;
        RECT  4.750 0.440 4.910 1.290 ;
        RECT  4.450 2.300 4.770 2.490 ;
        RECT  4.630 1.010 4.750 1.290 ;
        RECT  4.390 1.910 4.540 2.130 ;
        RECT  4.230 2.670 4.510 2.910 ;
        RECT  3.170 2.300 4.450 2.460 ;
        RECT  4.110 0.450 4.390 0.830 ;
        RECT  4.230 1.030 4.390 2.130 ;
        RECT  4.150 1.030 4.230 1.480 ;
        RECT  3.410 2.670 4.230 2.830 ;
        RECT  3.750 1.320 4.150 1.480 ;
        RECT  2.730 0.550 4.110 0.830 ;
        RECT  3.470 1.200 3.750 1.480 ;
        RECT  3.130 2.670 3.410 2.900 ;
        RECT  3.050 2.180 3.170 2.460 ;
        RECT  2.730 2.670 3.130 2.830 ;
        RECT  2.890 0.990 3.050 2.460 ;
        RECT  2.570 0.550 2.730 2.830 ;
        RECT  2.250 0.640 2.410 2.780 ;
        RECT  0.710 0.640 2.250 0.800 ;
        RECT  0.710 2.620 2.250 2.780 ;
        RECT  1.930 0.960 2.090 1.500 ;
        RECT  0.970 0.960 1.930 1.120 ;
        RECT  0.810 0.960 0.970 1.310 ;
        RECT  0.710 1.030 0.810 1.310 ;
        RECT  0.490 0.470 0.710 0.800 ;
        RECT  0.550 1.030 0.710 2.190 ;
        RECT  0.480 2.500 0.710 2.780 ;
    END
END SDFFSX4TR

MACRO SDFFSX2TR
    CLASS CORE ;
    FOREIGN SDFFSX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.240 8.080 1.640 ;
        RECT  7.680 1.240 7.740 3.160 ;
        RECT  7.580 1.480 7.680 3.160 ;
        RECT  6.820 2.940 7.580 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.580 1.330 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.580 0.400 1.860 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.480 0.600 10.720 3.090 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.760 1.030 9.920 2.760 ;
        RECT  9.390 1.030 9.760 1.310 ;
        RECT  9.390 2.000 9.760 2.760 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.040 1.920 2.360 ;
        RECT  1.550 1.330 1.710 2.360 ;
        RECT  1.370 2.170 1.550 2.360 ;
        RECT  1.090 2.170 1.370 2.450 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.640 4.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.190 -0.280 10.800 0.280 ;
        RECT  9.910 -0.280 10.190 0.420 ;
        RECT  8.440 -0.280 9.910 0.280 ;
        RECT  8.160 -0.280 8.440 0.740 ;
        RECT  3.950 -0.280 8.160 0.280 ;
        RECT  3.670 -0.280 3.950 0.390 ;
        RECT  1.610 -0.280 3.670 0.340 ;
        RECT  1.330 -0.280 1.610 0.400 ;
        RECT  0.350 -0.280 1.330 0.280 ;
        RECT  0.350 1.030 0.400 1.310 ;
        RECT  0.080 -0.280 0.350 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.190 3.320 10.800 3.880 ;
        RECT  9.910 3.240 10.190 3.880 ;
        RECT  8.220 3.320 9.910 3.880 ;
        RECT  7.940 2.400 8.220 3.880 ;
        RECT  6.660 3.320 7.940 3.880 ;
        RECT  6.440 2.850 6.660 3.880 ;
        RECT  5.000 3.320 6.440 3.880 ;
        RECT  4.720 2.990 5.000 3.880 ;
        RECT  3.950 3.320 4.720 3.880 ;
        RECT  3.670 2.990 3.950 3.880 ;
        RECT  1.610 3.260 3.670 3.880 ;
        RECT  1.330 3.200 1.610 3.880 ;
        RECT  0.090 3.260 1.330 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.260 1.520 10.320 1.800 ;
        RECT  10.100 0.710 10.260 3.080 ;
        RECT  9.140 0.710 10.100 0.870 ;
        RECT  8.890 2.920 10.100 3.080 ;
        RECT  9.210 1.480 9.600 1.760 ;
        RECT  9.050 1.030 9.210 2.190 ;
        RECT  8.860 0.440 9.140 0.870 ;
        RECT  8.650 1.030 9.050 1.310 ;
        RECT  7.900 1.910 9.050 2.190 ;
        RECT  8.610 2.920 8.890 3.160 ;
        RECT  8.490 1.470 8.520 1.750 ;
        RECT  8.330 0.920 8.490 1.750 ;
        RECT  7.420 0.920 8.330 1.080 ;
        RECT  7.580 0.440 7.860 0.760 ;
        RECT  5.080 0.440 7.580 0.600 ;
        RECT  7.260 0.760 7.420 2.780 ;
        RECT  6.720 0.760 7.260 0.920 ;
        RECT  6.940 2.380 7.260 2.780 ;
        RECT  6.880 1.200 7.100 2.220 ;
        RECT  6.720 2.380 6.940 2.540 ;
        RECT  6.680 1.200 6.880 1.360 ;
        RECT  6.440 1.910 6.720 2.540 ;
        RECT  6.280 1.080 6.680 1.360 ;
        RECT  5.540 0.760 6.440 0.920 ;
        RECT  6.120 1.080 6.280 3.160 ;
        RECT  5.700 1.080 6.120 1.300 ;
        RECT  5.560 3.000 6.120 3.160 ;
        RECT  5.740 1.460 5.960 2.590 ;
        RECT  5.540 1.460 5.740 1.620 ;
        RECT  5.280 2.220 5.560 3.160 ;
        RECT  5.380 0.760 5.540 1.620 ;
        RECT  4.600 1.450 5.380 1.610 ;
        RECT  5.110 1.780 5.330 2.060 ;
        RECT  5.160 2.990 5.280 3.160 ;
        RECT  4.950 1.780 5.110 2.830 ;
        RECT  4.920 0.440 5.080 1.290 ;
        RECT  4.510 2.670 4.950 2.830 ;
        RECT  4.800 1.010 4.920 1.290 ;
        RECT  3.190 2.330 4.790 2.490 ;
        RECT  4.440 1.030 4.600 1.610 ;
        RECT  4.440 1.910 4.560 2.130 ;
        RECT  2.750 0.550 4.510 0.830 ;
        RECT  4.230 2.670 4.510 2.890 ;
        RECT  4.280 1.030 4.440 2.130 ;
        RECT  3.830 1.320 4.280 1.480 ;
        RECT  3.430 2.670 4.230 2.830 ;
        RECT  3.550 1.200 3.830 1.480 ;
        RECT  3.150 2.670 3.430 2.900 ;
        RECT  2.910 0.990 3.190 2.490 ;
        RECT  2.750 2.670 3.150 2.830 ;
        RECT  2.590 0.550 2.750 2.830 ;
        RECT  2.270 0.690 2.430 2.780 ;
        RECT  0.730 0.690 2.270 0.850 ;
        RECT  0.730 2.620 2.270 2.780 ;
        RECT  1.890 1.010 2.110 1.500 ;
        RECT  0.990 1.010 1.890 1.170 ;
        RECT  0.720 1.010 0.990 1.310 ;
        RECT  0.720 2.120 0.930 2.400 ;
        RECT  0.510 0.470 0.730 0.850 ;
        RECT  0.480 2.620 0.730 2.990 ;
        RECT  0.560 1.010 0.720 2.400 ;
    END
END SDFFSX2TR

MACRO SDFFSX1TR
    CLASS CORE ;
    FOREIGN SDFFSX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.240 8.080 1.640 ;
        RECT  7.580 1.240 7.740 3.160 ;
        RECT  6.820 2.940 7.580 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.580 1.330 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.580 0.400 1.860 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.080 1.030 10.320 2.450 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.270 1.030 9.350 1.310 ;
        RECT  9.110 1.030 9.270 2.760 ;
        RECT  8.880 2.440 9.110 2.760 ;
        END
        ANTENNADIFFAREA 1.604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 2.040 1.920 2.360 ;
        RECT  1.550 1.330 1.710 2.360 ;
        RECT  1.370 2.170 1.550 2.360 ;
        RECT  1.090 2.170 1.370 2.450 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.640 4.120 2.040 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.910 -0.280 10.400 0.280 ;
        RECT  9.630 -0.280 9.910 0.420 ;
        RECT  8.470 -0.280 9.630 0.280 ;
        RECT  8.180 -0.280 8.470 0.760 ;
        RECT  3.950 -0.280 8.180 0.280 ;
        RECT  3.670 -0.280 3.950 0.390 ;
        RECT  1.610 -0.280 3.670 0.340 ;
        RECT  1.330 -0.280 1.610 0.400 ;
        RECT  0.350 -0.280 1.330 0.280 ;
        RECT  0.350 1.030 0.400 1.310 ;
        RECT  0.080 -0.280 0.350 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.790 3.320 10.400 3.880 ;
        RECT  9.430 3.240 9.790 3.880 ;
        RECT  8.220 3.320 9.430 3.880 ;
        RECT  7.940 2.460 8.220 3.880 ;
        RECT  6.660 3.320 7.940 3.880 ;
        RECT  6.440 2.850 6.660 3.880 ;
        RECT  5.000 3.320 6.440 3.880 ;
        RECT  4.720 2.990 5.000 3.880 ;
        RECT  3.950 3.320 4.720 3.880 ;
        RECT  3.670 2.990 3.950 3.880 ;
        RECT  1.610 3.260 3.670 3.880 ;
        RECT  1.330 3.200 1.610 3.880 ;
        RECT  0.090 3.260 1.330 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.670 1.700 9.790 1.980 ;
        RECT  9.510 0.710 9.670 3.080 ;
        RECT  9.140 0.710 9.510 0.870 ;
        RECT  8.850 2.920 9.510 3.080 ;
        RECT  8.860 0.440 9.140 0.870 ;
        RECT  8.870 1.030 8.950 1.730 ;
        RECT  8.710 1.030 8.870 2.190 ;
        RECT  8.570 2.920 8.850 3.160 ;
        RECT  8.650 1.030 8.710 1.310 ;
        RECT  7.900 1.910 8.710 2.190 ;
        RECT  8.490 1.470 8.520 1.750 ;
        RECT  8.330 0.920 8.490 1.750 ;
        RECT  7.420 0.920 8.330 1.080 ;
        RECT  7.580 0.440 7.860 0.760 ;
        RECT  5.080 0.440 7.580 0.600 ;
        RECT  7.260 0.760 7.420 2.780 ;
        RECT  6.720 0.760 7.260 0.920 ;
        RECT  6.940 2.380 7.260 2.780 ;
        RECT  6.880 1.200 7.100 2.220 ;
        RECT  6.720 2.380 6.940 2.540 ;
        RECT  6.680 1.200 6.880 1.360 ;
        RECT  6.440 1.910 6.720 2.540 ;
        RECT  6.280 1.080 6.680 1.360 ;
        RECT  5.540 0.760 6.440 0.920 ;
        RECT  6.120 1.080 6.280 3.160 ;
        RECT  5.700 1.080 6.120 1.300 ;
        RECT  5.560 3.000 6.120 3.160 ;
        RECT  5.740 1.460 5.960 2.590 ;
        RECT  5.540 1.460 5.740 1.620 ;
        RECT  5.280 2.220 5.560 3.160 ;
        RECT  5.380 0.760 5.540 1.620 ;
        RECT  4.600 1.450 5.380 1.610 ;
        RECT  5.110 1.780 5.330 2.060 ;
        RECT  5.160 2.990 5.280 3.160 ;
        RECT  4.950 1.780 5.110 2.830 ;
        RECT  4.920 0.440 5.080 1.290 ;
        RECT  4.510 2.670 4.950 2.830 ;
        RECT  4.800 1.010 4.920 1.290 ;
        RECT  3.190 2.330 4.790 2.490 ;
        RECT  4.440 1.030 4.600 1.610 ;
        RECT  4.440 1.910 4.560 2.130 ;
        RECT  2.750 0.550 4.510 0.830 ;
        RECT  4.230 2.670 4.510 2.890 ;
        RECT  4.280 1.030 4.440 2.130 ;
        RECT  3.830 1.320 4.280 1.480 ;
        RECT  3.430 2.670 4.230 2.830 ;
        RECT  3.550 1.200 3.830 1.480 ;
        RECT  3.150 2.670 3.430 2.900 ;
        RECT  2.910 0.990 3.190 2.490 ;
        RECT  2.750 2.670 3.150 2.830 ;
        RECT  2.590 0.550 2.750 2.830 ;
        RECT  2.270 0.690 2.430 2.780 ;
        RECT  0.730 0.690 2.270 0.850 ;
        RECT  0.730 2.620 2.270 2.780 ;
        RECT  1.890 1.010 2.110 1.500 ;
        RECT  0.990 1.010 1.890 1.170 ;
        RECT  0.720 1.010 0.990 1.310 ;
        RECT  0.720 2.120 0.930 2.400 ;
        RECT  0.510 0.470 0.730 0.850 ;
        RECT  0.480 2.620 0.730 2.990 ;
        RECT  0.560 1.010 0.720 2.400 ;
    END
END SDFFSX1TR

MACRO SDFFRHQX8TR
    CLASS CORE ;
    FOREIGN SDFFRHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.240 5.920 1.560 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.160 2.770 1.640 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.320 1.670 13.480 1.950 ;
        RECT  11.240 1.790 13.320 1.950 ;
        RECT  11.080 1.240 11.240 1.950 ;
        RECT  10.880 1.240 11.080 1.560 ;
        RECT  10.170 1.240 10.880 1.400 ;
        RECT  10.010 1.240 10.170 1.520 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.660 0.580 16.940 3.160 ;
        RECT  16.020 1.040 16.660 1.760 ;
        RECT  15.700 0.630 16.020 2.990 ;
        END
        ANTENNADIFFAREA 7.668 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.500 3.660 1.780 ;
        RECT  3.280 1.240 3.520 1.780 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.100 0.720 1.560 ;
        END
        ANTENNAGATEAREA 0.3936 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.420 -0.280 17.600 0.280 ;
        RECT  17.150 -0.280 17.420 1.210 ;
        RECT  16.460 -0.280 17.150 0.280 ;
        RECT  16.200 -0.280 16.460 0.870 ;
        RECT  15.490 -0.280 16.200 0.280 ;
        RECT  15.210 -0.280 15.490 1.280 ;
        RECT  14.390 -0.280 15.210 0.280 ;
        RECT  14.110 -0.280 14.390 0.290 ;
        RECT  11.670 -0.280 14.110 0.280 ;
        RECT  11.390 -0.280 11.670 0.290 ;
        RECT  9.990 -0.280 11.390 0.280 ;
        RECT  9.710 -0.280 9.990 0.290 ;
        RECT  8.820 -0.280 9.710 0.280 ;
        RECT  8.540 -0.280 8.820 0.340 ;
        RECT  7.180 -0.280 8.540 0.280 ;
        RECT  6.900 -0.280 7.180 0.940 ;
        RECT  5.520 -0.280 6.900 0.280 ;
        RECT  5.240 -0.280 5.520 0.340 ;
        RECT  3.440 -0.280 5.240 0.280 ;
        RECT  3.160 -0.280 3.440 0.290 ;
        RECT  0.790 -0.280 3.160 0.280 ;
        RECT  0.510 -0.280 0.790 0.290 ;
        RECT  0.000 -0.280 0.510 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.400 3.320 17.600 3.880 ;
        RECT  17.150 2.010 17.400 3.880 ;
        RECT  16.450 3.320 17.150 3.880 ;
        RECT  16.180 2.010 16.450 3.880 ;
        RECT  15.260 3.320 16.180 3.880 ;
        RECT  14.940 2.870 15.260 3.880 ;
        RECT  13.880 3.320 14.940 3.880 ;
        RECT  13.610 2.920 13.880 3.880 ;
        RECT  10.980 3.320 13.610 3.880 ;
        RECT  10.700 3.230 10.980 3.880 ;
        RECT  9.940 3.320 10.700 3.880 ;
        RECT  9.660 3.230 9.940 3.880 ;
        RECT  8.440 3.320 9.660 3.880 ;
        RECT  8.160 3.260 8.440 3.880 ;
        RECT  6.760 3.320 8.160 3.880 ;
        RECT  6.480 3.260 6.760 3.880 ;
        RECT  5.840 3.320 6.480 3.880 ;
        RECT  5.560 3.260 5.840 3.880 ;
        RECT  3.650 3.320 5.560 3.880 ;
        RECT  3.370 2.930 3.650 3.880 ;
        RECT  2.690 3.320 3.370 3.880 ;
        RECT  2.400 2.990 2.690 3.880 ;
        RECT  0.560 3.260 2.400 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.230 1.540 15.500 1.700 ;
        RECT  15.070 1.540 15.230 2.710 ;
        RECT  14.630 2.550 15.070 2.710 ;
        RECT  14.690 1.030 14.890 2.190 ;
        RECT  14.600 1.430 14.690 1.710 ;
        RECT  14.350 2.550 14.630 3.160 ;
        RECT  14.280 0.450 14.440 2.280 ;
        RECT  14.120 2.550 14.350 2.710 ;
        RECT  13.300 0.450 14.280 0.610 ;
        RECT  13.960 0.770 14.120 2.710 ;
        RECT  11.950 0.770 13.960 0.930 ;
        RECT  11.920 2.550 13.960 2.710 ;
        RECT  13.640 1.210 13.800 2.390 ;
        RECT  12.490 1.210 13.640 1.370 ;
        RECT  12.400 2.230 13.640 2.390 ;
        RECT  13.020 0.440 13.300 0.610 ;
        RECT  9.340 0.450 13.020 0.610 ;
        RECT  12.210 1.090 12.490 1.370 ;
        RECT  12.240 2.110 12.400 2.390 ;
        RECT  11.440 2.110 12.240 2.270 ;
        RECT  11.560 1.210 12.210 1.370 ;
        RECT  11.790 0.770 11.950 1.050 ;
        RECT  11.760 2.430 11.920 2.710 ;
        RECT  9.210 2.880 11.780 3.040 ;
        RECT  11.400 0.920 11.560 1.370 ;
        RECT  11.280 2.110 11.440 2.390 ;
        RECT  10.550 0.920 11.400 1.080 ;
        RECT  10.460 2.110 11.280 2.270 ;
        RECT  10.410 1.560 10.570 1.840 ;
        RECT  10.180 2.110 10.460 2.670 ;
        RECT  9.850 1.680 10.410 1.840 ;
        RECT  9.530 2.110 10.180 2.270 ;
        RECT  9.690 1.040 9.850 1.840 ;
        RECT  8.890 1.040 9.690 1.250 ;
        RECT  9.370 1.580 9.530 2.270 ;
        RECT  9.180 0.450 9.340 0.860 ;
        RECT  9.050 2.240 9.210 3.040 ;
        RECT  7.540 0.700 9.180 0.860 ;
        RECT  7.220 2.880 9.050 3.040 ;
        RECT  8.730 1.040 8.890 2.720 ;
        RECT  7.700 1.040 8.730 1.200 ;
        RECT  7.540 2.560 8.730 2.720 ;
        RECT  8.360 1.360 8.520 2.280 ;
        RECT  7.220 2.120 8.360 2.280 ;
        RECT  7.540 1.800 8.200 1.960 ;
        RECT  7.380 0.700 7.540 1.960 ;
        RECT  7.380 2.440 7.540 2.720 ;
        RECT  6.680 1.100 7.380 1.260 ;
        RECT  7.060 1.420 7.220 3.040 ;
        RECT  6.940 1.420 7.060 1.580 ;
        RECT  3.970 2.880 7.060 3.040 ;
        RECT  6.560 1.760 6.900 2.040 ;
        RECT  6.580 0.440 6.740 0.720 ;
        RECT  6.560 0.990 6.680 1.260 ;
        RECT  6.240 0.560 6.580 0.720 ;
        RECT  6.400 0.990 6.560 2.570 ;
        RECT  4.290 2.410 6.400 2.570 ;
        RECT  6.080 0.560 6.240 2.040 ;
        RECT  4.620 0.890 6.080 1.050 ;
        RECT  5.100 1.880 6.080 2.040 ;
        RECT  5.680 0.440 5.840 0.720 ;
        RECT  4.940 0.560 5.680 0.720 ;
        RECT  4.300 1.560 5.360 1.720 ;
        RECT  4.940 1.880 5.100 2.160 ;
        RECT  4.780 0.450 4.940 0.720 ;
        RECT  1.040 0.450 4.780 0.610 ;
        RECT  4.460 0.770 4.620 1.050 ;
        RECT  4.460 1.970 4.620 2.250 ;
        RECT  3.980 1.970 4.460 2.130 ;
        RECT  4.140 0.770 4.300 1.720 ;
        RECT  4.130 2.290 4.290 2.570 ;
        RECT  3.120 0.770 4.140 0.930 ;
        RECT  2.210 2.290 4.130 2.450 ;
        RECT  3.820 1.090 3.980 2.130 ;
        RECT  3.810 2.610 3.970 3.040 ;
        RECT  3.680 1.090 3.820 1.250 ;
        RECT  3.440 1.970 3.820 2.130 ;
        RECT  1.700 2.610 3.810 2.770 ;
        RECT  2.960 0.770 3.120 2.130 ;
        RECT  2.780 0.770 2.960 0.930 ;
        RECT  2.690 1.970 2.960 2.130 ;
        RECT  2.470 0.770 2.780 1.000 ;
        RECT  2.200 1.590 2.210 2.450 ;
        RECT  2.050 1.560 2.200 2.450 ;
        RECT  1.380 0.980 2.080 1.160 ;
        RECT  1.730 1.560 2.050 1.870 ;
        RECT  1.540 2.250 1.700 2.770 ;
        RECT  1.380 2.250 1.540 2.420 ;
        RECT  1.200 0.980 1.380 2.420 ;
        RECT  0.880 0.450 1.040 1.880 ;
        RECT  0.710 0.700 0.880 0.860 ;
        RECT  0.310 1.720 0.880 1.880 ;
        RECT  0.150 1.720 0.310 2.200 ;
    END
END SDFFRHQX8TR

MACRO SDFFRHQX4TR
    CLASS CORE ;
    FOREIGN SDFFRHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.240 5.920 1.560 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.160 2.770 1.640 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.320 1.670 13.480 1.950 ;
        RECT  11.240 1.790 13.320 1.950 ;
        RECT  11.080 1.240 11.240 1.950 ;
        RECT  10.880 1.240 11.080 1.560 ;
        RECT  10.170 1.240 10.880 1.400 ;
        RECT  10.010 1.240 10.170 1.520 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.610 0.630 15.920 2.990 ;
        END
        ANTENNADIFFAREA 3.834 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.500 3.660 1.780 ;
        RECT  3.280 1.240 3.520 1.780 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.100 0.720 1.560 ;
        END
        ANTENNAGATEAREA 0.3936 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.250 -0.280 16.400 0.280 ;
        RECT  16.090 -0.280 16.250 1.210 ;
        RECT  15.310 -0.280 16.090 0.280 ;
        RECT  15.030 -0.280 15.310 0.340 ;
        RECT  14.390 -0.280 15.030 0.280 ;
        RECT  14.110 -0.280 14.390 0.290 ;
        RECT  11.670 -0.280 14.110 0.280 ;
        RECT  11.390 -0.280 11.670 0.290 ;
        RECT  9.990 -0.280 11.390 0.280 ;
        RECT  9.710 -0.280 9.990 0.290 ;
        RECT  8.820 -0.280 9.710 0.280 ;
        RECT  8.540 -0.280 8.820 0.340 ;
        RECT  7.180 -0.280 8.540 0.280 ;
        RECT  6.900 -0.280 7.180 0.940 ;
        RECT  5.520 -0.280 6.900 0.280 ;
        RECT  5.240 -0.280 5.520 0.340 ;
        RECT  3.440 -0.280 5.240 0.280 ;
        RECT  3.160 -0.280 3.440 0.290 ;
        RECT  0.790 -0.280 3.160 0.280 ;
        RECT  0.510 -0.280 0.790 0.290 ;
        RECT  0.000 -0.280 0.510 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.250 3.320 16.400 3.880 ;
        RECT  16.090 2.010 16.250 3.880 ;
        RECT  15.260 3.320 16.090 3.880 ;
        RECT  14.940 2.870 15.260 3.880 ;
        RECT  13.880 3.320 14.940 3.880 ;
        RECT  13.610 2.920 13.880 3.880 ;
        RECT  10.980 3.320 13.610 3.880 ;
        RECT  10.700 3.230 10.980 3.880 ;
        RECT  9.940 3.320 10.700 3.880 ;
        RECT  9.660 3.230 9.940 3.880 ;
        RECT  8.440 3.320 9.660 3.880 ;
        RECT  8.160 3.260 8.440 3.880 ;
        RECT  6.760 3.320 8.160 3.880 ;
        RECT  6.480 3.260 6.760 3.880 ;
        RECT  5.840 3.320 6.480 3.880 ;
        RECT  5.560 3.260 5.840 3.880 ;
        RECT  3.650 3.320 5.560 3.880 ;
        RECT  3.370 2.930 3.650 3.880 ;
        RECT  2.690 3.320 3.370 3.880 ;
        RECT  2.400 2.990 2.690 3.880 ;
        RECT  0.560 3.260 2.400 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.230 1.540 15.350 1.700 ;
        RECT  15.070 1.540 15.230 2.710 ;
        RECT  14.630 2.550 15.070 2.710 ;
        RECT  14.690 1.030 14.890 2.190 ;
        RECT  14.600 1.430 14.690 1.710 ;
        RECT  14.350 2.550 14.630 3.160 ;
        RECT  14.280 0.450 14.440 2.280 ;
        RECT  14.120 2.550 14.350 2.710 ;
        RECT  13.300 0.450 14.280 0.610 ;
        RECT  13.960 0.770 14.120 2.710 ;
        RECT  11.950 0.770 13.960 0.930 ;
        RECT  11.920 2.550 13.960 2.710 ;
        RECT  13.640 1.210 13.800 2.390 ;
        RECT  12.490 1.210 13.640 1.370 ;
        RECT  12.400 2.230 13.640 2.390 ;
        RECT  13.020 0.440 13.300 0.610 ;
        RECT  9.340 0.450 13.020 0.610 ;
        RECT  12.210 1.090 12.490 1.370 ;
        RECT  12.240 2.110 12.400 2.390 ;
        RECT  11.440 2.110 12.240 2.270 ;
        RECT  11.560 1.210 12.210 1.370 ;
        RECT  11.790 0.770 11.950 1.050 ;
        RECT  11.760 2.430 11.920 2.710 ;
        RECT  9.210 2.880 11.780 3.040 ;
        RECT  11.400 0.920 11.560 1.370 ;
        RECT  11.280 2.110 11.440 2.390 ;
        RECT  10.550 0.920 11.400 1.080 ;
        RECT  10.460 2.110 11.280 2.270 ;
        RECT  10.410 1.560 10.570 1.840 ;
        RECT  10.180 2.110 10.460 2.670 ;
        RECT  9.850 1.680 10.410 1.840 ;
        RECT  9.530 2.110 10.180 2.270 ;
        RECT  9.690 1.040 9.850 1.840 ;
        RECT  8.890 1.040 9.690 1.250 ;
        RECT  9.370 1.580 9.530 2.270 ;
        RECT  9.180 0.450 9.340 0.860 ;
        RECT  9.050 2.240 9.210 3.040 ;
        RECT  7.540 0.700 9.180 0.860 ;
        RECT  7.220 2.880 9.050 3.040 ;
        RECT  8.730 1.040 8.890 2.720 ;
        RECT  7.700 1.040 8.730 1.200 ;
        RECT  7.540 2.560 8.730 2.720 ;
        RECT  8.360 1.360 8.520 2.280 ;
        RECT  7.220 2.120 8.360 2.280 ;
        RECT  7.540 1.800 8.200 1.960 ;
        RECT  7.380 0.700 7.540 1.960 ;
        RECT  7.380 2.440 7.540 2.720 ;
        RECT  6.680 1.100 7.380 1.260 ;
        RECT  7.060 1.420 7.220 3.040 ;
        RECT  6.940 1.420 7.060 1.580 ;
        RECT  3.970 2.880 7.060 3.040 ;
        RECT  6.560 1.760 6.900 2.040 ;
        RECT  6.580 0.440 6.740 0.720 ;
        RECT  6.560 0.990 6.680 1.260 ;
        RECT  6.240 0.560 6.580 0.720 ;
        RECT  6.400 0.990 6.560 2.570 ;
        RECT  4.290 2.410 6.400 2.570 ;
        RECT  6.080 0.560 6.240 2.040 ;
        RECT  4.620 0.890 6.080 1.050 ;
        RECT  5.100 1.880 6.080 2.040 ;
        RECT  5.680 0.440 5.840 0.720 ;
        RECT  4.940 0.560 5.680 0.720 ;
        RECT  4.300 1.560 5.360 1.720 ;
        RECT  4.940 1.880 5.100 2.160 ;
        RECT  4.780 0.450 4.940 0.720 ;
        RECT  1.040 0.450 4.780 0.610 ;
        RECT  4.460 0.770 4.620 1.050 ;
        RECT  4.460 1.970 4.620 2.250 ;
        RECT  3.980 1.970 4.460 2.130 ;
        RECT  4.140 0.770 4.300 1.720 ;
        RECT  4.130 2.290 4.290 2.570 ;
        RECT  3.120 0.770 4.140 0.930 ;
        RECT  2.210 2.290 4.130 2.450 ;
        RECT  3.820 1.090 3.980 2.130 ;
        RECT  3.810 2.610 3.970 3.040 ;
        RECT  3.680 1.090 3.820 1.250 ;
        RECT  3.440 1.970 3.820 2.130 ;
        RECT  1.700 2.610 3.810 2.770 ;
        RECT  2.960 0.770 3.120 2.130 ;
        RECT  2.780 0.770 2.960 0.930 ;
        RECT  2.690 1.970 2.960 2.130 ;
        RECT  2.470 0.770 2.780 1.000 ;
        RECT  2.200 1.590 2.210 2.450 ;
        RECT  2.050 1.560 2.200 2.450 ;
        RECT  1.380 0.980 2.080 1.160 ;
        RECT  1.730 1.560 2.050 1.870 ;
        RECT  1.540 2.250 1.700 2.770 ;
        RECT  1.380 2.250 1.540 2.420 ;
        RECT  1.200 0.980 1.380 2.420 ;
        RECT  0.880 0.450 1.040 1.880 ;
        RECT  0.710 0.700 0.880 0.860 ;
        RECT  0.310 1.720 0.880 1.880 ;
        RECT  0.150 1.720 0.310 2.200 ;
    END
END SDFFRHQX4TR

MACRO SDFFRHQX2TR
    CLASS CORE ;
    FOREIGN SDFFRHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.320 4.360 1.960 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.160 1.440 9.280 1.600 ;
        RECT  9.000 1.440 9.160 2.010 ;
        RECT  8.340 1.850 9.000 2.010 ;
        RECT  8.220 1.850 8.340 2.060 ;
        RECT  8.060 1.850 8.220 2.340 ;
        RECT  7.520 2.180 8.060 2.340 ;
        RECT  7.360 1.560 7.520 2.340 ;
        RECT  7.280 1.560 7.360 1.960 ;
        RECT  7.220 1.560 7.280 1.720 ;
        END
        ANTENNAGATEAREA 0.2376 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.080 0.440 12.320 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.380 2.360 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.790 -0.280 12.400 0.280 ;
        RECT  11.510 -0.280 11.790 1.270 ;
        RECT  7.260 -0.280 11.510 0.280 ;
        RECT  6.980 -0.280 7.260 0.340 ;
        RECT  5.360 -0.280 6.980 0.280 ;
        RECT  5.080 -0.280 5.360 0.340 ;
        RECT  4.420 -0.280 5.080 0.280 ;
        RECT  4.140 -0.280 4.420 0.340 ;
        RECT  2.540 -0.280 4.140 0.280 ;
        RECT  2.260 -0.280 2.540 0.340 ;
        RECT  0.940 -0.280 2.260 0.280 ;
        RECT  0.660 -0.280 0.940 0.340 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.830 3.320 12.400 3.880 ;
        RECT  11.530 2.930 11.830 3.880 ;
        RECT  10.230 3.320 11.530 3.880 ;
        RECT  9.950 2.930 10.230 3.880 ;
        RECT  8.100 3.320 9.950 3.880 ;
        RECT  7.820 3.260 8.100 3.880 ;
        RECT  7.180 3.320 7.820 3.880 ;
        RECT  6.900 3.260 7.180 3.880 ;
        RECT  5.540 3.320 6.900 3.880 ;
        RECT  5.260 3.260 5.540 3.880 ;
        RECT  4.540 3.320 5.260 3.880 ;
        RECT  4.260 3.260 4.540 3.880 ;
        RECT  2.360 3.320 4.260 3.880 ;
        RECT  2.200 2.940 2.360 3.880 ;
        RECT  0.880 3.320 2.200 3.880 ;
        RECT  0.580 3.180 0.880 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.490 1.540 11.650 2.770 ;
        RECT  11.050 2.610 11.490 2.770 ;
        RECT  11.170 1.580 11.330 2.190 ;
        RECT  11.010 1.030 11.170 1.740 ;
        RECT  10.890 2.610 11.050 2.890 ;
        RECT  10.400 1.580 11.010 1.740 ;
        RECT  9.920 2.610 10.890 2.770 ;
        RECT  10.240 2.230 10.870 2.390 ;
        RECT  10.080 0.440 10.240 2.390 ;
        RECT  7.580 0.440 10.080 0.600 ;
        RECT  9.760 0.760 9.920 2.770 ;
        RECT  6.780 2.940 9.790 3.100 ;
        RECT  8.520 0.760 9.760 0.920 ;
        RECT  9.040 2.610 9.760 2.770 ;
        RECT  9.440 1.080 9.600 2.450 ;
        RECT  8.840 1.080 9.440 1.240 ;
        RECT  9.360 2.170 9.440 2.450 ;
        RECT  8.660 2.170 9.360 2.330 ;
        RECT  8.880 2.490 9.040 2.770 ;
        RECT  8.680 1.080 8.840 1.370 ;
        RECT  8.160 1.210 8.680 1.370 ;
        RECT  8.500 2.170 8.660 2.660 ;
        RECT  8.360 0.760 8.520 1.050 ;
        RECT  8.400 2.290 8.500 2.660 ;
        RECT  7.640 2.500 8.400 2.660 ;
        RECT  8.000 0.910 8.160 1.370 ;
        RECT  7.820 0.910 8.000 1.070 ;
        RECT  7.680 1.230 7.840 2.020 ;
        RECT  6.320 1.230 7.680 1.390 ;
        RECT  7.480 2.500 7.640 2.780 ;
        RECT  7.420 0.440 7.580 0.920 ;
        RECT  7.040 2.500 7.480 2.660 ;
        RECT  6.710 0.760 7.420 0.920 ;
        RECT  6.880 1.840 7.040 2.660 ;
        RECT  6.500 2.900 6.780 3.100 ;
        RECT  6.550 0.580 6.710 0.920 ;
        RECT  6.000 0.760 6.550 0.920 ;
        RECT  5.780 2.940 6.500 3.100 ;
        RECT  6.160 1.230 6.320 2.680 ;
        RECT  5.680 0.440 6.180 0.600 ;
        RECT  6.080 2.310 6.160 2.680 ;
        RECT  5.840 0.760 6.000 1.300 ;
        RECT  5.320 1.140 5.840 1.300 ;
        RECT  5.620 1.560 5.780 3.100 ;
        RECT  5.520 0.440 5.680 0.980 ;
        RECT  5.500 1.560 5.620 1.720 ;
        RECT  2.680 2.940 5.620 3.100 ;
        RECT  4.680 0.820 5.520 0.980 ;
        RECT  5.160 1.140 5.320 2.780 ;
        RECT  4.880 1.140 5.160 1.420 ;
        RECT  3.000 2.620 5.160 2.780 ;
        RECT  0.700 0.500 4.870 0.660 ;
        RECT  4.520 0.820 4.680 2.340 ;
        RECT  4.500 0.820 4.520 1.160 ;
        RECT  3.580 2.180 4.520 2.340 ;
        RECT  3.520 1.000 4.500 1.160 ;
        RECT  3.760 1.320 3.920 2.000 ;
        RECT  3.360 1.320 3.760 1.480 ;
        RECT  3.200 0.820 3.360 1.480 ;
        RECT  3.160 1.640 3.320 2.460 ;
        RECT  1.020 0.820 3.200 0.980 ;
        RECT  3.040 1.640 3.160 1.800 ;
        RECT  2.880 1.140 3.040 1.800 ;
        RECT  2.840 2.120 3.000 2.780 ;
        RECT  2.720 1.140 2.880 1.300 ;
        RECT  2.120 2.120 2.840 2.280 ;
        RECT  2.520 2.590 2.680 3.100 ;
        RECT  1.800 2.590 2.520 2.750 ;
        RECT  1.960 1.720 2.120 2.280 ;
        RECT  1.660 1.720 1.960 1.880 ;
        RECT  1.200 3.000 1.900 3.160 ;
        RECT  1.640 2.040 1.800 2.750 ;
        RECT  1.500 1.600 1.660 1.880 ;
        RECT  1.340 2.040 1.640 2.200 ;
        RECT  1.340 1.140 1.500 1.360 ;
        RECT  1.180 1.140 1.340 2.200 ;
        RECT  1.040 2.360 1.200 3.160 ;
        RECT  1.020 2.360 1.040 2.520 ;
        RECT  0.860 0.820 1.020 2.520 ;
        RECT  0.540 0.500 0.700 2.680 ;
        RECT  0.370 0.500 0.540 0.660 ;
        RECT  0.230 2.520 0.540 2.680 ;
        RECT  0.090 0.440 0.370 0.660 ;
    END
END SDFFRHQX2TR

MACRO SDFFRHQX1TR
    CLASS CORE ;
    FOREIGN SDFFRHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.360 1.580 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.240 2.320 1.640 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.060 1.580 9.220 2.030 ;
        RECT  8.160 1.640 9.060 2.030 ;
        RECT  7.460 1.870 8.160 2.030 ;
        RECT  7.300 1.380 7.460 2.030 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.520 0.840 11.760 2.650 ;
        RECT  11.280 0.840 11.520 1.960 ;
        END
        ANTENNADIFFAREA 1.92 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.270 -0.280 12.000 0.280 ;
        RECT  10.920 -0.280 11.270 0.670 ;
        RECT  9.970 -0.280 10.920 0.280 ;
        RECT  9.690 -0.280 9.970 0.340 ;
        RECT  7.250 -0.280 9.690 0.280 ;
        RECT  6.970 -0.280 7.250 0.340 ;
        RECT  5.730 -0.280 6.970 0.280 ;
        RECT  5.450 -0.280 5.730 0.290 ;
        RECT  4.700 -0.280 5.450 0.280 ;
        RECT  4.420 -0.280 4.700 0.290 ;
        RECT  2.480 -0.280 4.420 0.280 ;
        RECT  2.200 -0.280 2.480 0.290 ;
        RECT  0.840 -0.280 2.200 0.280 ;
        RECT  0.560 -0.280 0.840 0.290 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.300 3.320 12.000 3.880 ;
        RECT  11.060 2.320 11.300 3.880 ;
        RECT  9.600 3.320 11.060 3.880 ;
        RECT  9.320 2.930 9.600 3.880 ;
        RECT  8.120 3.320 9.320 3.880 ;
        RECT  7.840 3.260 8.120 3.880 ;
        RECT  7.320 3.320 7.840 3.880 ;
        RECT  7.040 3.260 7.320 3.880 ;
        RECT  5.550 3.320 7.040 3.880 ;
        RECT  5.270 3.260 5.550 3.880 ;
        RECT  4.460 3.320 5.270 3.880 ;
        RECT  4.180 3.260 4.460 3.880 ;
        RECT  2.200 3.320 4.180 3.880 ;
        RECT  2.040 2.760 2.200 3.880 ;
        RECT  0.840 3.320 2.040 3.880 ;
        RECT  0.560 3.260 0.840 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.900 1.580 11.030 1.860 ;
        RECT  10.740 1.580 10.900 2.540 ;
        RECT  10.500 2.370 10.740 2.540 ;
        RECT  10.420 1.020 10.580 2.190 ;
        RECT  10.200 2.370 10.500 2.670 ;
        RECT  10.340 1.430 10.420 1.710 ;
        RECT  9.860 2.510 10.200 2.670 ;
        RECT  10.020 0.620 10.180 2.210 ;
        RECT  8.510 0.620 10.020 0.780 ;
        RECT  9.700 0.940 9.860 2.670 ;
        RECT  8.360 0.940 9.700 1.100 ;
        RECT  9.160 2.510 9.700 2.670 ;
        RECT  9.380 1.260 9.540 2.350 ;
        RECT  8.180 1.260 9.380 1.420 ;
        RECT  8.620 2.190 9.380 2.350 ;
        RECT  8.880 2.510 9.160 2.730 ;
        RECT  6.050 2.940 8.810 3.100 ;
        RECT  8.460 2.190 8.620 2.470 ;
        RECT  8.230 0.480 8.510 0.780 ;
        RECT  7.660 2.310 8.460 2.470 ;
        RECT  6.670 0.620 8.230 0.780 ;
        RECT  8.020 0.950 8.180 1.420 ;
        RECT  7.940 0.950 8.020 1.230 ;
        RECT  7.780 1.430 7.860 1.710 ;
        RECT  7.620 1.020 7.780 1.710 ;
        RECT  7.500 2.190 7.660 2.470 ;
        RECT  6.990 1.020 7.620 1.180 ;
        RECT  6.960 2.310 7.500 2.470 ;
        RECT  6.960 1.690 7.080 1.980 ;
        RECT  6.830 1.020 6.990 1.250 ;
        RECT  6.800 1.690 6.960 2.470 ;
        RECT  6.430 1.090 6.830 1.250 ;
        RECT  6.510 0.480 6.670 0.930 ;
        RECT  6.040 0.770 6.510 0.930 ;
        RECT  6.210 1.090 6.430 2.370 ;
        RECT  5.720 0.450 6.250 0.610 ;
        RECT  5.890 1.420 6.050 3.100 ;
        RECT  5.880 0.770 6.040 1.250 ;
        RECT  5.550 1.420 5.890 1.580 ;
        RECT  2.520 2.940 5.890 3.100 ;
        RECT  5.040 1.090 5.880 1.250 ;
        RECT  5.570 1.760 5.730 2.040 ;
        RECT  5.560 0.450 5.720 0.930 ;
        RECT  5.100 1.880 5.570 2.040 ;
        RECT  4.200 0.770 5.560 0.930 ;
        RECT  0.640 0.450 5.290 0.610 ;
        RECT  5.040 1.880 5.100 2.690 ;
        RECT  4.880 1.090 5.040 2.690 ;
        RECT  2.840 2.530 4.880 2.690 ;
        RECT  4.040 0.770 4.200 2.360 ;
        RECT  3.690 0.770 4.040 0.930 ;
        RECT  3.420 2.200 4.040 2.360 ;
        RECT  3.660 1.210 3.820 2.040 ;
        RECT  3.530 0.770 3.690 1.050 ;
        RECT  3.360 1.210 3.660 1.370 ;
        RECT  3.600 1.760 3.660 2.040 ;
        RECT  3.200 0.770 3.360 1.370 ;
        RECT  0.960 0.770 3.200 0.930 ;
        RECT  3.040 1.530 3.160 2.370 ;
        RECT  3.000 1.090 3.040 2.370 ;
        RECT  2.880 1.090 3.000 1.690 ;
        RECT  2.740 1.090 2.880 1.310 ;
        RECT  2.680 2.120 2.840 2.690 ;
        RECT  2.120 2.120 2.680 2.280 ;
        RECT  2.360 2.440 2.520 3.100 ;
        RECT  1.800 2.440 2.360 2.600 ;
        RECT  1.960 1.800 2.120 2.280 ;
        RECT  1.600 1.800 1.960 1.960 ;
        RECT  1.640 2.120 1.800 2.600 ;
        RECT  1.460 2.810 1.740 3.090 ;
        RECT  1.280 2.120 1.640 2.280 ;
        RECT  1.440 1.540 1.600 1.960 ;
        RECT  0.960 2.870 1.460 3.030 ;
        RECT  1.280 1.090 1.400 1.310 ;
        RECT  1.120 1.090 1.280 2.280 ;
        RECT  0.800 0.770 0.960 3.030 ;
        RECT  0.480 0.450 0.640 2.830 ;
        RECT  0.120 0.860 0.480 1.080 ;
        RECT  0.090 2.610 0.480 2.830 ;
    END
END SDFFRHQX1TR

MACRO SDFFRXLTR
    CLASS CORE ;
    FOREIGN SDFFRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 2.840 2.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.640 1.470 1.960 ;
        RECT  0.760 1.800 1.190 1.960 ;
        RECT  0.400 1.640 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.430 1.360 8.690 1.640 ;
        RECT  8.050 1.360 8.430 1.520 ;
        RECT  7.890 0.470 8.050 1.520 ;
        RECT  6.810 0.470 7.890 0.630 ;
        RECT  6.650 0.470 6.810 1.010 ;
        RECT  6.490 0.850 6.650 1.010 ;
        RECT  6.210 0.850 6.490 1.510 ;
        RECT  6.170 0.850 6.210 1.010 ;
        RECT  6.010 0.440 6.170 1.010 ;
        RECT  4.150 0.440 6.010 0.600 ;
        RECT  3.990 0.440 4.150 0.700 ;
        RECT  2.720 0.540 3.990 0.700 ;
        RECT  2.560 0.540 2.720 1.640 ;
        RECT  2.480 0.840 2.560 1.640 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.270 1.640 10.320 2.390 ;
        RECT  10.110 1.030 10.270 2.390 ;
        RECT  9.810 1.030 10.110 1.310 ;
        RECT  10.080 1.640 10.110 2.390 ;
        RECT  9.850 2.110 10.080 2.390 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.830 0.840 11.120 2.390 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.770 1.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.290 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.550 -0.280 11.200 0.280 ;
        RECT  10.270 -0.280 10.550 0.400 ;
        RECT  8.490 -0.280 10.270 0.280 ;
        RECT  8.210 -0.280 8.490 0.740 ;
        RECT  6.490 -0.280 8.210 0.280 ;
        RECT  6.330 -0.280 6.490 0.690 ;
        RECT  3.830 -0.280 6.330 0.280 ;
        RECT  2.930 -0.280 3.830 0.340 ;
        RECT  2.650 -0.280 2.930 0.380 ;
        RECT  0.370 -0.280 2.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.590 3.320 11.200 3.880 ;
        RECT  9.290 3.200 10.590 3.880 ;
        RECT  8.080 3.320 9.290 3.880 ;
        RECT  7.800 3.200 8.080 3.880 ;
        RECT  5.670 3.320 7.800 3.880 ;
        RECT  5.390 2.450 5.670 3.880 ;
        RECT  3.630 3.320 5.390 3.880 ;
        RECT  3.350 3.200 3.630 3.880 ;
        RECT  2.600 3.260 3.350 3.880 ;
        RECT  2.320 2.740 2.600 3.880 ;
        RECT  0.680 3.320 2.320 3.880 ;
        RECT  0.400 2.800 0.680 3.880 ;
        RECT  0.000 3.320 0.400 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.640 2.600 10.920 2.880 ;
        RECT  9.010 2.680 10.640 2.880 ;
        RECT  9.650 1.670 9.730 1.950 ;
        RECT  9.650 0.450 9.710 0.670 ;
        RECT  9.490 0.450 9.650 2.520 ;
        RECT  9.430 0.450 9.490 0.670 ;
        RECT  9.370 2.240 9.490 2.520 ;
        RECT  9.010 1.030 9.330 1.310 ;
        RECT  8.850 1.030 9.010 3.160 ;
        RECT  8.290 1.900 8.850 2.060 ;
        RECT  8.260 2.940 8.850 3.160 ;
        RECT  8.470 2.500 8.690 2.780 ;
        RECT  7.730 2.500 8.470 2.660 ;
        RECT  8.010 1.780 8.290 2.060 ;
        RECT  7.570 0.790 7.730 2.880 ;
        RECT  7.450 0.790 7.570 1.070 ;
        RECT  7.190 2.720 7.570 2.880 ;
        RECT  7.130 2.310 7.410 2.560 ;
        RECT  6.970 0.790 7.190 1.830 ;
        RECT  6.910 2.720 7.190 2.990 ;
        RECT  6.750 2.310 7.130 2.470 ;
        RECT  6.370 1.670 6.970 1.830 ;
        RECT  6.590 2.310 6.750 2.940 ;
        RECT  5.990 2.780 6.590 2.940 ;
        RECT  6.370 2.340 6.430 2.620 ;
        RECT  6.150 1.670 6.370 2.620 ;
        RECT  5.850 1.170 5.990 2.940 ;
        RECT  5.830 0.760 5.850 2.940 ;
        RECT  5.690 0.760 5.830 1.330 ;
        RECT  4.470 0.760 5.690 0.920 ;
        RECT  5.510 2.010 5.670 2.290 ;
        RECT  5.290 1.080 5.530 1.300 ;
        RECT  5.230 2.010 5.510 2.170 ;
        RECT  5.230 1.080 5.290 1.620 ;
        RECT  5.130 1.080 5.230 3.020 ;
        RECT  5.070 1.460 5.130 3.020 ;
        RECT  4.710 2.860 5.070 3.020 ;
        RECT  4.850 1.080 4.970 1.300 ;
        RECT  4.690 1.080 4.850 2.510 ;
        RECT  4.430 2.860 4.710 3.160 ;
        RECT  4.190 2.350 4.690 2.510 ;
        RECT  4.470 1.380 4.530 1.660 ;
        RECT  4.410 0.760 4.470 1.660 ;
        RECT  3.170 2.860 4.430 3.020 ;
        RECT  4.310 0.760 4.410 2.130 ;
        RECT  4.250 0.980 4.310 2.130 ;
        RECT  4.110 0.980 4.250 1.260 ;
        RECT  3.870 1.910 4.250 2.130 ;
        RECT  3.910 2.350 4.190 2.650 ;
        RECT  2.230 2.350 3.910 2.580 ;
        RECT  3.550 0.860 3.710 2.070 ;
        RECT  3.110 0.860 3.550 1.080 ;
        RECT  3.170 1.910 3.550 2.070 ;
        RECT  2.890 1.910 3.170 2.190 ;
        RECT  2.890 2.740 3.170 3.020 ;
        RECT  0.830 0.500 2.400 0.660 ;
        RECT  2.070 0.820 2.230 2.580 ;
        RECT  1.430 0.820 2.070 0.980 ;
        RECT  1.430 2.360 2.070 2.580 ;
        RECT  1.630 1.220 1.910 2.160 ;
        RECT  0.830 1.220 1.630 1.380 ;
        RECT  0.550 0.500 0.830 0.800 ;
        RECT  0.550 1.030 0.830 1.380 ;
        RECT  0.240 1.220 0.550 1.380 ;
        RECT  0.240 2.120 0.370 2.400 ;
        RECT  0.080 1.220 0.240 2.400 ;
    END
END SDFFRXLTR

MACRO SDFFRX4TR
    CLASS CORE ;
    FOREIGN SDFFRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 2.840 2.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.640 1.470 1.960 ;
        RECT  0.760 1.800 1.190 1.960 ;
        RECT  0.400 1.640 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.430 1.360 8.690 1.640 ;
        RECT  8.050 1.360 8.430 1.520 ;
        RECT  7.890 0.470 8.050 1.520 ;
        RECT  6.790 0.470 7.890 0.630 ;
        RECT  6.630 0.470 6.790 1.010 ;
        RECT  6.490 0.850 6.630 1.010 ;
        RECT  6.210 0.850 6.490 1.510 ;
        RECT  6.150 0.850 6.210 1.010 ;
        RECT  5.990 0.440 6.150 1.010 ;
        RECT  4.150 0.440 5.990 0.600 ;
        RECT  3.990 0.440 4.150 0.700 ;
        RECT  2.720 0.540 3.990 0.700 ;
        RECT  2.560 0.540 2.720 1.640 ;
        RECT  2.480 0.840 2.560 1.640 ;
        END
        ANTENNAGATEAREA 0.3024 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.890 1.030 11.120 1.760 ;
        RECT  10.590 0.600 10.890 2.390 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.860 0.840 11.920 1.760 ;
        RECT  11.680 0.840 11.860 3.060 ;
        RECT  11.550 0.840 11.680 1.170 ;
        RECT  11.600 1.930 11.680 3.060 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.770 1.200 3.160 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.290 1.620 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 -0.280 12.400 0.280 ;
        RECT  12.080 -0.280 12.310 1.150 ;
        RECT  11.350 -0.280 12.080 0.280 ;
        RECT  11.070 -0.280 11.350 0.860 ;
        RECT  10.300 -0.280 11.070 0.280 ;
        RECT  10.020 -0.280 10.300 1.170 ;
        RECT  8.490 -0.280 10.020 0.280 ;
        RECT  8.210 -0.280 8.490 0.740 ;
        RECT  6.470 -0.280 8.210 0.280 ;
        RECT  6.310 -0.280 6.470 0.690 ;
        RECT  3.830 -0.280 6.310 0.280 ;
        RECT  2.930 -0.280 3.830 0.340 ;
        RECT  2.650 -0.280 2.930 0.380 ;
        RECT  0.370 -0.280 2.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 3.320 12.400 3.880 ;
        RECT  12.070 2.080 12.310 3.880 ;
        RECT  11.350 3.320 12.070 3.880 ;
        RECT  11.070 2.990 11.350 3.880 ;
        RECT  10.390 3.320 11.070 3.880 ;
        RECT  10.110 2.990 10.390 3.880 ;
        RECT  9.270 3.320 10.110 3.880 ;
        RECT  8.990 3.260 9.270 3.880 ;
        RECT  8.160 3.320 8.990 3.880 ;
        RECT  7.870 2.730 8.160 3.880 ;
        RECT  5.670 3.320 7.870 3.880 ;
        RECT  5.390 2.450 5.670 3.880 ;
        RECT  3.630 3.320 5.390 3.880 ;
        RECT  3.350 3.200 3.630 3.880 ;
        RECT  2.600 3.260 3.350 3.880 ;
        RECT  2.320 2.740 2.600 3.880 ;
        RECT  0.720 3.320 2.320 3.880 ;
        RECT  0.440 2.800 0.720 3.880 ;
        RECT  0.000 3.320 0.440 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.280 1.530 11.440 2.830 ;
        RECT  9.600 2.670 11.280 2.830 ;
        RECT  9.790 1.530 10.430 1.750 ;
        RECT  9.630 0.450 9.790 2.510 ;
        RECT  9.400 0.450 9.630 0.670 ;
        RECT  9.510 2.230 9.630 2.510 ;
        RECT  9.270 2.670 9.600 3.100 ;
        RECT  9.270 1.030 9.350 1.320 ;
        RECT  9.110 1.030 9.270 3.100 ;
        RECT  9.070 1.030 9.110 1.960 ;
        RECT  8.450 2.940 9.110 3.100 ;
        RECT  8.050 1.800 9.070 1.960 ;
        RECT  8.760 2.200 8.950 2.480 ;
        RECT  8.730 2.220 8.760 2.480 ;
        RECT  7.670 2.220 8.730 2.380 ;
        RECT  7.830 1.780 8.050 2.060 ;
        RECT  7.510 0.790 7.670 2.930 ;
        RECT  7.450 0.790 7.510 1.070 ;
        RECT  6.910 2.770 7.510 2.930 ;
        RECT  7.120 2.310 7.350 2.610 ;
        RECT  6.950 0.790 7.170 1.830 ;
        RECT  6.750 2.450 7.120 2.610 ;
        RECT  6.370 1.670 6.950 1.830 ;
        RECT  6.590 2.450 6.750 2.940 ;
        RECT  5.990 2.780 6.590 2.940 ;
        RECT  6.370 2.340 6.430 2.620 ;
        RECT  6.150 1.670 6.370 2.620 ;
        RECT  5.830 1.170 5.990 2.940 ;
        RECT  5.670 0.760 5.830 1.330 ;
        RECT  4.530 0.760 5.670 0.920 ;
        RECT  5.510 2.010 5.670 2.290 ;
        RECT  5.230 2.010 5.510 2.170 ;
        RECT  5.290 1.080 5.470 1.360 ;
        RECT  5.230 1.080 5.290 1.620 ;
        RECT  5.130 1.080 5.230 3.020 ;
        RECT  5.070 1.460 5.130 3.020 ;
        RECT  4.710 2.860 5.070 3.020 ;
        RECT  4.850 1.080 4.970 1.300 ;
        RECT  4.690 1.080 4.850 2.510 ;
        RECT  4.430 2.860 4.710 3.160 ;
        RECT  4.190 2.350 4.690 2.510 ;
        RECT  4.410 0.760 4.530 1.660 ;
        RECT  3.170 2.860 4.430 3.020 ;
        RECT  4.310 0.760 4.410 2.130 ;
        RECT  4.250 0.980 4.310 2.130 ;
        RECT  4.110 0.980 4.250 1.260 ;
        RECT  3.870 1.910 4.250 2.130 ;
        RECT  3.910 2.350 4.190 2.650 ;
        RECT  2.230 2.350 3.910 2.580 ;
        RECT  3.550 0.860 3.710 2.070 ;
        RECT  3.110 0.860 3.550 1.080 ;
        RECT  3.170 1.910 3.550 2.070 ;
        RECT  2.890 1.910 3.170 2.190 ;
        RECT  2.890 2.740 3.170 3.020 ;
        RECT  0.830 0.500 2.400 0.660 ;
        RECT  2.070 0.820 2.230 2.580 ;
        RECT  1.430 0.820 2.070 0.980 ;
        RECT  1.430 2.360 2.070 2.580 ;
        RECT  1.630 1.220 1.910 2.160 ;
        RECT  0.830 1.220 1.630 1.380 ;
        RECT  0.550 0.500 0.830 0.800 ;
        RECT  0.550 1.030 0.830 1.380 ;
        RECT  0.240 1.220 0.550 1.380 ;
        RECT  0.240 2.120 0.370 2.400 ;
        RECT  0.080 1.220 0.240 2.400 ;
    END
END SDFFRX4TR

MACRO SDFFRX2TR
    CLASS CORE ;
    FOREIGN SDFFRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 2.840 2.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.640 1.470 1.960 ;
        RECT  0.760 1.800 1.190 1.960 ;
        RECT  0.400 1.640 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.430 1.360 8.690 1.640 ;
        RECT  8.050 1.360 8.430 1.520 ;
        RECT  7.890 0.470 8.050 1.520 ;
        RECT  6.790 0.470 7.890 0.630 ;
        RECT  6.630 0.470 6.790 1.010 ;
        RECT  6.490 0.850 6.630 1.010 ;
        RECT  6.210 0.850 6.490 1.510 ;
        RECT  6.150 0.850 6.210 1.010 ;
        RECT  5.990 0.440 6.150 1.010 ;
        RECT  4.150 0.440 5.990 0.600 ;
        RECT  3.990 0.440 4.150 0.700 ;
        RECT  2.720 0.540 3.990 0.700 ;
        RECT  2.560 0.540 2.720 1.640 ;
        RECT  2.480 0.840 2.560 1.640 ;
        END
        ANTENNAGATEAREA 0.2184 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.270 1.640 10.320 2.390 ;
        RECT  10.110 1.030 10.270 2.390 ;
        RECT  9.870 1.030 10.110 1.310 ;
        RECT  10.080 1.640 10.110 2.390 ;
        RECT  9.870 2.110 10.080 2.390 ;
        END
        ANTENNADIFFAREA 3.25 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.880 0.840 11.120 3.010 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.770 1.200 3.160 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.290 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.630 -0.280 11.200 0.280 ;
        RECT  10.350 -0.280 10.630 0.860 ;
        RECT  8.490 -0.280 10.350 0.280 ;
        RECT  8.210 -0.280 8.490 0.740 ;
        RECT  6.470 -0.280 8.210 0.280 ;
        RECT  6.310 -0.280 6.470 0.690 ;
        RECT  3.830 -0.280 6.310 0.280 ;
        RECT  2.930 -0.280 3.830 0.340 ;
        RECT  2.650 -0.280 2.930 0.380 ;
        RECT  0.370 -0.280 2.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.630 3.320 11.200 3.880 ;
        RECT  10.350 2.990 10.630 3.880 ;
        RECT  9.270 3.320 10.350 3.880 ;
        RECT  8.990 3.260 9.270 3.880 ;
        RECT  8.170 3.320 8.990 3.880 ;
        RECT  7.890 2.800 8.170 3.880 ;
        RECT  5.670 3.320 7.890 3.880 ;
        RECT  5.390 2.450 5.670 3.880 ;
        RECT  3.630 3.320 5.390 3.880 ;
        RECT  3.350 3.200 3.630 3.880 ;
        RECT  2.600 3.260 3.350 3.880 ;
        RECT  2.320 2.740 2.600 3.880 ;
        RECT  0.720 3.320 2.320 3.880 ;
        RECT  0.440 2.800 0.720 3.880 ;
        RECT  0.000 3.320 0.440 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.560 1.530 10.720 2.830 ;
        RECT  9.480 2.670 10.560 2.830 ;
        RECT  9.670 0.450 9.810 0.670 ;
        RECT  9.670 1.670 9.730 1.950 ;
        RECT  9.650 2.230 9.690 2.510 ;
        RECT  9.650 0.450 9.670 1.950 ;
        RECT  9.510 0.450 9.650 2.510 ;
        RECT  9.490 1.410 9.510 2.510 ;
        RECT  9.410 2.230 9.490 2.510 ;
        RECT  9.230 2.670 9.480 2.890 ;
        RECT  9.230 1.030 9.350 1.250 ;
        RECT  9.070 1.030 9.230 3.100 ;
        RECT  8.290 1.900 9.070 2.060 ;
        RECT  8.470 2.940 9.070 3.100 ;
        RECT  8.660 2.220 8.880 2.780 ;
        RECT  7.730 2.220 8.660 2.380 ;
        RECT  8.010 1.780 8.290 2.060 ;
        RECT  7.570 0.790 7.730 2.880 ;
        RECT  7.450 0.790 7.570 1.070 ;
        RECT  7.190 2.720 7.570 2.880 ;
        RECT  7.130 2.310 7.410 2.560 ;
        RECT  6.910 2.720 7.190 2.990 ;
        RECT  6.950 0.790 7.170 1.830 ;
        RECT  6.750 2.310 7.130 2.470 ;
        RECT  6.370 1.670 6.950 1.830 ;
        RECT  6.590 2.310 6.750 2.940 ;
        RECT  5.990 2.780 6.590 2.940 ;
        RECT  6.370 2.340 6.430 2.620 ;
        RECT  6.150 1.670 6.370 2.620 ;
        RECT  5.830 1.170 5.990 2.940 ;
        RECT  5.670 0.760 5.830 1.330 ;
        RECT  4.470 0.760 5.670 0.920 ;
        RECT  5.510 2.010 5.670 2.290 ;
        RECT  5.230 2.010 5.510 2.170 ;
        RECT  5.290 1.080 5.470 1.360 ;
        RECT  5.230 1.080 5.290 1.620 ;
        RECT  5.130 1.080 5.230 3.020 ;
        RECT  5.070 1.460 5.130 3.020 ;
        RECT  4.710 2.860 5.070 3.020 ;
        RECT  4.850 1.080 4.970 1.300 ;
        RECT  4.690 1.080 4.850 2.510 ;
        RECT  4.430 2.860 4.710 3.160 ;
        RECT  4.190 2.350 4.690 2.510 ;
        RECT  4.470 1.380 4.530 1.660 ;
        RECT  4.410 0.760 4.470 1.660 ;
        RECT  3.170 2.860 4.430 3.020 ;
        RECT  4.310 0.760 4.410 2.130 ;
        RECT  4.250 0.980 4.310 2.130 ;
        RECT  4.110 0.980 4.250 1.260 ;
        RECT  3.870 1.910 4.250 2.130 ;
        RECT  3.910 2.350 4.190 2.650 ;
        RECT  2.230 2.350 3.910 2.580 ;
        RECT  3.550 0.860 3.710 2.070 ;
        RECT  3.110 0.860 3.550 1.080 ;
        RECT  3.170 1.910 3.550 2.070 ;
        RECT  2.890 1.910 3.170 2.190 ;
        RECT  2.890 2.740 3.170 3.020 ;
        RECT  0.830 0.500 2.400 0.660 ;
        RECT  2.070 0.820 2.230 2.580 ;
        RECT  1.430 0.820 2.070 0.980 ;
        RECT  1.430 2.360 2.070 2.580 ;
        RECT  1.630 1.220 1.910 2.160 ;
        RECT  0.830 1.220 1.630 1.380 ;
        RECT  0.550 0.500 0.830 0.800 ;
        RECT  0.550 1.030 0.830 1.380 ;
        RECT  0.240 1.220 0.550 1.380 ;
        RECT  0.240 2.120 0.370 2.400 ;
        RECT  0.080 1.220 0.240 2.400 ;
    END
END SDFFRX2TR

MACRO SDFFRX1TR
    CLASS CORE ;
    FOREIGN SDFFRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 2.840 2.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.640 1.470 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.430 1.360 8.690 1.720 ;
        RECT  8.050 1.360 8.430 1.520 ;
        RECT  7.890 0.470 8.050 1.520 ;
        RECT  6.810 0.470 7.890 0.630 ;
        RECT  6.650 0.470 6.810 1.010 ;
        RECT  6.490 0.850 6.650 1.010 ;
        RECT  6.210 0.850 6.490 1.510 ;
        RECT  6.170 0.850 6.210 1.010 ;
        RECT  6.010 0.440 6.170 1.010 ;
        RECT  4.150 0.440 6.010 0.600 ;
        RECT  3.990 0.440 4.150 0.700 ;
        RECT  2.720 0.540 3.990 0.700 ;
        RECT  2.560 0.540 2.720 1.640 ;
        RECT  2.480 0.840 2.560 1.640 ;
        END
        ANTENNAGATEAREA 0.1824 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.080 1.030 10.320 2.390 ;
        RECT  9.870 1.030 10.080 1.310 ;
        RECT  9.850 2.120 10.080 2.390 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.830 0.840 11.120 2.190 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.770 1.220 3.160 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.360 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.670 -0.280 11.200 0.280 ;
        RECT  10.390 -0.280 10.670 0.400 ;
        RECT  8.490 -0.280 10.390 0.280 ;
        RECT  8.210 -0.280 8.490 0.740 ;
        RECT  6.490 -0.280 8.210 0.280 ;
        RECT  6.330 -0.280 6.490 0.690 ;
        RECT  3.830 -0.280 6.330 0.280 ;
        RECT  2.930 -0.280 3.830 0.340 ;
        RECT  2.650 -0.280 2.930 0.380 ;
        RECT  0.370 -0.280 2.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.580 3.320 11.200 3.880 ;
        RECT  9.290 3.200 10.580 3.880 ;
        RECT  8.080 3.320 9.290 3.880 ;
        RECT  7.800 3.200 8.080 3.880 ;
        RECT  5.670 3.320 7.800 3.880 ;
        RECT  5.390 2.450 5.670 3.880 ;
        RECT  3.630 3.320 5.390 3.880 ;
        RECT  3.350 3.200 3.630 3.880 ;
        RECT  2.600 3.260 3.350 3.880 ;
        RECT  2.320 2.740 2.600 3.880 ;
        RECT  0.680 3.320 2.320 3.880 ;
        RECT  0.400 2.800 0.680 3.880 ;
        RECT  0.000 3.320 0.400 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.630 2.680 10.920 2.940 ;
        RECT  9.070 2.680 10.630 2.880 ;
        RECT  9.670 1.670 9.850 1.950 ;
        RECT  9.670 0.450 9.710 0.670 ;
        RECT  9.650 0.450 9.670 1.950 ;
        RECT  9.510 0.450 9.650 2.500 ;
        RECT  9.430 0.450 9.510 0.670 ;
        RECT  9.490 1.410 9.510 2.500 ;
        RECT  9.370 2.220 9.490 2.500 ;
        RECT  9.070 1.030 9.350 1.310 ;
        RECT  8.910 1.030 9.070 3.160 ;
        RECT  8.240 1.900 8.910 2.060 ;
        RECT  8.260 2.940 8.910 3.160 ;
        RECT  8.470 2.500 8.750 2.780 ;
        RECT  7.730 2.500 8.470 2.660 ;
        RECT  7.950 1.780 8.240 2.060 ;
        RECT  7.570 0.790 7.730 2.880 ;
        RECT  7.450 0.790 7.570 1.070 ;
        RECT  7.200 2.720 7.570 2.880 ;
        RECT  7.130 2.310 7.410 2.560 ;
        RECT  6.920 2.720 7.200 2.990 ;
        RECT  6.970 0.790 7.190 1.830 ;
        RECT  6.750 2.310 7.130 2.470 ;
        RECT  6.430 1.670 6.970 1.830 ;
        RECT  6.590 2.310 6.750 2.940 ;
        RECT  5.990 2.780 6.590 2.940 ;
        RECT  6.150 1.670 6.430 2.620 ;
        RECT  5.850 1.170 5.990 2.940 ;
        RECT  5.830 0.760 5.850 2.940 ;
        RECT  5.690 0.760 5.830 1.330 ;
        RECT  4.470 0.760 5.690 0.920 ;
        RECT  5.510 2.010 5.670 2.290 ;
        RECT  5.290 1.080 5.530 1.300 ;
        RECT  5.290 2.010 5.510 2.170 ;
        RECT  5.230 1.080 5.290 2.170 ;
        RECT  5.130 1.080 5.230 3.020 ;
        RECT  5.070 1.460 5.130 3.020 ;
        RECT  4.710 2.860 5.070 3.020 ;
        RECT  4.850 1.080 4.970 1.300 ;
        RECT  4.690 1.080 4.850 2.510 ;
        RECT  4.430 2.860 4.710 3.160 ;
        RECT  4.190 2.350 4.690 2.510 ;
        RECT  4.470 1.530 4.530 1.810 ;
        RECT  4.410 0.760 4.470 1.810 ;
        RECT  3.170 2.860 4.430 3.020 ;
        RECT  4.310 0.760 4.410 2.130 ;
        RECT  4.250 0.980 4.310 2.130 ;
        RECT  4.110 0.980 4.250 1.260 ;
        RECT  3.870 1.970 4.250 2.130 ;
        RECT  3.910 2.350 4.190 2.650 ;
        RECT  3.710 1.510 4.030 1.770 ;
        RECT  2.230 2.350 3.910 2.580 ;
        RECT  3.550 0.860 3.710 2.070 ;
        RECT  3.110 0.860 3.550 1.080 ;
        RECT  3.170 1.910 3.550 2.070 ;
        RECT  2.890 1.910 3.170 2.190 ;
        RECT  2.890 2.740 3.170 3.020 ;
        RECT  0.830 0.500 2.400 0.660 ;
        RECT  2.070 0.820 2.230 2.580 ;
        RECT  1.380 0.820 2.070 0.980 ;
        RECT  1.430 2.360 2.070 2.580 ;
        RECT  1.630 1.220 1.910 2.160 ;
        RECT  0.830 1.220 1.630 1.380 ;
        RECT  0.550 0.500 0.830 0.800 ;
        RECT  0.550 1.030 0.830 1.380 ;
        RECT  0.240 1.220 0.550 1.380 ;
        RECT  0.240 2.120 0.370 2.400 ;
        RECT  0.080 1.220 0.240 2.400 ;
    END
END SDFFRX1TR

MACRO SDFFQXLTR
    CLASS CORE ;
    FOREIGN SDFFQXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.640 1.520 2.080 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.920 1.960 2.360 ;
        RECT  1.680 1.920 1.840 2.720 ;
        RECT  0.420 2.560 1.680 2.720 ;
        RECT  0.260 1.550 0.420 2.720 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.640 0.770 8.720 2.910 ;
        RECT  8.560 0.440 8.640 2.910 ;
        RECT  8.480 0.440 8.560 0.930 ;
        RECT  8.470 2.440 8.560 2.910 ;
        RECT  8.080 2.440 8.470 2.760 ;
        END
        ANTENNADIFFAREA 1.102 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.100 2.320 1.560 ;
        RECT  2.060 1.280 2.080 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.040 2.040 4.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.100 -0.280 8.800 0.280 ;
        RECT  7.820 -0.280 8.100 0.610 ;
        RECT  5.960 -0.280 7.820 0.280 ;
        RECT  5.800 -0.280 5.960 0.700 ;
        RECT  4.530 -0.280 5.800 0.280 ;
        RECT  3.760 -0.280 4.530 0.640 ;
        RECT  1.760 -0.280 3.760 0.280 ;
        RECT  1.480 -0.280 1.760 0.340 ;
        RECT  0.310 -0.280 1.480 0.280 ;
        RECT  0.150 -0.280 0.310 1.310 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.920 3.320 8.800 3.880 ;
        RECT  7.620 2.630 7.920 3.880 ;
        RECT  6.120 3.320 7.620 3.880 ;
        RECT  5.840 3.260 6.120 3.880 ;
        RECT  4.920 3.320 5.840 3.880 ;
        RECT  4.640 3.260 4.920 3.880 ;
        RECT  3.940 3.320 4.640 3.880 ;
        RECT  3.660 3.260 3.940 3.880 ;
        RECT  1.840 3.320 3.660 3.880 ;
        RECT  1.560 3.260 1.840 3.880 ;
        RECT  0.370 3.320 1.560 3.880 ;
        RECT  0.090 3.050 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.240 1.090 8.400 2.230 ;
        RECT  8.120 1.090 8.240 1.250 ;
        RECT  8.120 1.800 8.240 2.230 ;
        RECT  7.640 1.800 8.120 1.960 ;
        RECT  7.820 1.350 7.980 1.640 ;
        RECT  7.180 1.350 7.820 1.510 ;
        RECT  7.380 1.680 7.640 1.960 ;
        RECT  7.020 1.090 7.180 3.160 ;
        RECT  6.780 1.090 7.020 1.250 ;
        RECT  6.780 0.550 6.940 0.890 ;
        RECT  6.700 1.500 6.860 2.990 ;
        RECT  6.620 0.730 6.780 0.890 ;
        RECT  6.620 1.500 6.700 1.780 ;
        RECT  4.340 2.830 6.700 2.990 ;
        RECT  6.460 0.730 6.620 1.780 ;
        RECT  6.380 2.110 6.540 2.670 ;
        RECT  6.060 1.500 6.460 1.780 ;
        RECT  5.900 2.110 6.380 2.270 ;
        RECT  5.200 2.510 6.380 2.670 ;
        RECT  6.140 1.000 6.300 1.310 ;
        RECT  5.900 1.150 6.140 1.310 ;
        RECT  5.740 1.150 5.900 2.270 ;
        RECT  5.420 0.690 5.580 2.270 ;
        RECT  5.330 0.690 5.420 0.850 ;
        RECT  5.150 0.440 5.330 0.850 ;
        RECT  5.200 1.110 5.260 1.880 ;
        RECT  5.100 1.110 5.200 2.670 ;
        RECT  4.810 0.440 5.150 0.600 ;
        RECT  5.040 1.720 5.100 2.670 ;
        RECT  3.680 1.720 5.040 1.880 ;
        RECT  3.120 1.400 4.940 1.560 ;
        RECT  3.430 1.020 4.420 1.180 ;
        RECT  4.180 2.520 4.340 2.990 ;
        RECT  3.360 2.830 4.180 2.990 ;
        RECT  3.520 1.720 3.680 2.000 ;
        RECT  3.270 0.610 3.430 1.180 ;
        RECT  3.200 2.830 3.360 3.110 ;
        RECT  2.670 0.610 3.270 0.770 ;
        RECT  2.800 2.830 3.200 2.990 ;
        RECT  3.110 1.400 3.120 2.670 ;
        RECT  2.960 0.930 3.110 2.670 ;
        RECT  2.950 0.930 2.960 1.560 ;
        RECT  2.830 0.930 2.950 1.210 ;
        RECT  2.670 1.720 2.800 2.990 ;
        RECT  2.670 1.370 2.790 1.530 ;
        RECT  2.640 0.610 2.670 2.990 ;
        RECT  2.510 0.610 2.640 1.880 ;
        RECT  2.200 2.880 2.480 3.140 ;
        RECT  2.070 0.480 2.350 0.720 ;
        RECT  0.900 2.880 2.200 3.040 ;
        RECT  0.800 0.560 2.070 0.720 ;
        RECT  0.870 1.320 1.880 1.480 ;
        RECT  0.870 2.240 1.200 2.400 ;
        RECT  0.740 2.880 0.900 3.160 ;
        RECT  0.710 1.030 0.870 2.400 ;
        RECT  0.640 0.440 0.800 0.720 ;
        RECT  0.590 1.910 0.710 2.190 ;
    END
END SDFFQXLTR

MACRO SDFFQX4TR
    CLASS CORE ;
    FOREIGN SDFFQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.640 1.520 2.080 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.920 1.960 2.360 ;
        RECT  1.680 1.920 1.840 2.720 ;
        RECT  0.420 2.560 1.680 2.720 ;
        RECT  0.260 1.550 0.420 2.720 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.980 0.620 9.260 3.020 ;
        RECT  8.880 1.240 8.980 2.360 ;
        END
        ANTENNADIFFAREA 4.07 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.100 2.320 1.560 ;
        RECT  2.060 1.280 2.080 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.040 2.040 4.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.750 -0.280 10.000 0.280 ;
        RECT  9.470 -0.280 9.750 1.170 ;
        RECT  8.780 -0.280 9.470 0.280 ;
        RECT  8.480 -0.280 8.780 1.070 ;
        RECT  7.740 -0.280 8.480 0.280 ;
        RECT  7.460 -0.280 7.740 0.610 ;
        RECT  5.960 -0.280 7.460 0.280 ;
        RECT  5.800 -0.280 5.960 0.700 ;
        RECT  4.530 -0.280 5.800 0.280 ;
        RECT  3.760 -0.280 4.530 0.640 ;
        RECT  1.760 -0.280 3.760 0.280 ;
        RECT  1.480 -0.280 1.760 0.340 ;
        RECT  0.310 -0.280 1.480 0.280 ;
        RECT  0.150 -0.280 0.310 1.310 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.750 3.320 10.000 3.880 ;
        RECT  9.450 2.040 9.750 3.880 ;
        RECT  8.780 3.320 9.450 3.880 ;
        RECT  8.480 2.530 8.780 3.880 ;
        RECT  7.910 3.320 8.480 3.880 ;
        RECT  7.620 2.820 7.910 3.880 ;
        RECT  6.120 3.320 7.620 3.880 ;
        RECT  5.840 3.260 6.120 3.880 ;
        RECT  4.920 3.320 5.840 3.880 ;
        RECT  4.640 3.260 4.920 3.880 ;
        RECT  3.940 3.320 4.640 3.880 ;
        RECT  3.660 3.260 3.940 3.880 ;
        RECT  1.840 3.320 3.660 3.880 ;
        RECT  1.560 3.260 1.840 3.880 ;
        RECT  0.370 3.320 1.560 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.320 1.480 8.600 1.740 ;
        RECT  8.160 0.980 8.320 2.230 ;
        RECT  8.040 0.980 8.160 1.140 ;
        RECT  8.020 1.800 8.160 2.230 ;
        RECT  7.640 1.800 8.020 1.960 ;
        RECT  7.820 1.350 7.980 1.640 ;
        RECT  7.180 1.350 7.820 1.510 ;
        RECT  7.380 1.680 7.640 1.960 ;
        RECT  6.620 0.630 7.240 0.790 ;
        RECT  7.020 1.010 7.180 3.160 ;
        RECT  6.780 1.010 7.020 1.310 ;
        RECT  6.700 1.630 6.860 2.990 ;
        RECT  6.620 1.630 6.700 1.790 ;
        RECT  4.340 2.830 6.700 2.990 ;
        RECT  6.460 0.630 6.620 1.790 ;
        RECT  6.380 2.110 6.540 2.670 ;
        RECT  6.060 1.500 6.460 1.790 ;
        RECT  5.900 2.110 6.380 2.270 ;
        RECT  5.200 2.510 6.380 2.670 ;
        RECT  6.140 1.000 6.300 1.310 ;
        RECT  5.900 1.150 6.140 1.310 ;
        RECT  5.740 1.150 5.900 2.270 ;
        RECT  5.420 0.690 5.580 2.270 ;
        RECT  5.330 0.690 5.420 0.850 ;
        RECT  5.150 0.440 5.330 0.850 ;
        RECT  5.200 1.110 5.260 1.880 ;
        RECT  5.100 1.110 5.200 2.670 ;
        RECT  4.810 0.440 5.150 0.600 ;
        RECT  5.040 1.720 5.100 2.670 ;
        RECT  3.680 1.720 5.040 1.880 ;
        RECT  3.120 1.400 4.940 1.560 ;
        RECT  3.430 1.020 4.420 1.180 ;
        RECT  4.180 2.520 4.340 2.990 ;
        RECT  3.360 2.830 4.180 2.990 ;
        RECT  3.520 1.720 3.680 2.000 ;
        RECT  3.270 0.610 3.430 1.180 ;
        RECT  3.200 2.830 3.360 3.110 ;
        RECT  2.670 0.610 3.270 0.770 ;
        RECT  2.800 2.830 3.200 2.990 ;
        RECT  3.110 1.400 3.120 2.670 ;
        RECT  2.960 0.930 3.110 2.670 ;
        RECT  2.950 0.930 2.960 1.560 ;
        RECT  2.830 0.930 2.950 1.210 ;
        RECT  2.670 1.720 2.800 2.990 ;
        RECT  2.670 1.370 2.790 1.530 ;
        RECT  2.640 0.610 2.670 2.990 ;
        RECT  2.510 0.610 2.640 1.880 ;
        RECT  2.200 2.880 2.480 3.140 ;
        RECT  2.070 0.480 2.350 0.720 ;
        RECT  0.900 2.880 2.200 3.040 ;
        RECT  0.800 0.560 2.070 0.720 ;
        RECT  0.870 1.320 1.880 1.480 ;
        RECT  0.870 2.240 1.200 2.400 ;
        RECT  0.740 2.880 0.900 3.160 ;
        RECT  0.710 1.030 0.870 2.400 ;
        RECT  0.640 0.440 0.800 0.720 ;
        RECT  0.590 1.910 0.710 2.190 ;
    END
END SDFFQX4TR

MACRO SDFFQX2TR
    CLASS CORE ;
    FOREIGN SDFFQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.640 1.520 1.990 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.890 1.960 2.360 ;
        RECT  1.680 1.890 1.840 2.720 ;
        RECT  0.370 2.560 1.680 2.720 ;
        RECT  0.090 1.580 0.370 2.720 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.350 0.630 8.720 3.000 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.240 2.320 1.640 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 2.040 4.400 2.370 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 -0.280 9.200 0.280 ;
        RECT  8.890 -0.280 9.110 1.070 ;
        RECT  7.610 -0.280 8.890 0.280 ;
        RECT  7.330 -0.280 7.610 0.720 ;
        RECT  5.930 -0.280 7.330 0.280 ;
        RECT  5.650 -0.280 5.930 0.850 ;
        RECT  4.300 -0.280 5.650 0.280 ;
        RECT  3.620 -0.280 4.300 0.650 ;
        RECT  0.370 -0.280 3.620 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 3.320 9.200 3.880 ;
        RECT  8.890 2.110 9.110 3.880 ;
        RECT  7.730 3.320 8.890 3.880 ;
        RECT  7.450 2.630 7.730 3.880 ;
        RECT  5.920 3.320 7.450 3.880 ;
        RECT  5.640 3.260 5.920 3.880 ;
        RECT  4.900 3.320 5.640 3.880 ;
        RECT  3.640 3.260 4.900 3.880 ;
        RECT  1.840 3.320 3.640 3.880 ;
        RECT  1.560 3.200 1.840 3.880 ;
        RECT  0.410 3.320 1.560 3.880 ;
        RECT  0.130 3.200 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.030 0.950 8.190 2.520 ;
        RECT  7.950 0.950 8.030 1.230 ;
        RECT  7.850 1.830 8.030 2.520 ;
        RECT  7.490 1.830 7.850 2.070 ;
        RECT  7.020 1.270 7.750 1.550 ;
        RECT  7.210 1.790 7.490 2.070 ;
        RECT  6.470 0.590 7.090 0.870 ;
        RECT  6.960 1.270 7.020 3.110 ;
        RECT  6.800 1.030 6.960 3.110 ;
        RECT  6.630 1.030 6.800 1.310 ;
        RECT  6.480 1.590 6.640 3.050 ;
        RECT  6.470 1.590 6.480 1.750 ;
        RECT  4.380 2.830 6.480 3.050 ;
        RECT  6.310 0.590 6.470 1.750 ;
        RECT  6.100 1.910 6.320 2.670 ;
        RECT  5.940 1.470 6.310 1.750 ;
        RECT  5.930 1.030 6.150 1.310 ;
        RECT  5.780 1.910 6.100 2.070 ;
        RECT  5.140 2.450 6.100 2.670 ;
        RECT  5.780 1.150 5.930 1.310 ;
        RECT  5.620 1.150 5.780 2.070 ;
        RECT  5.300 0.610 5.460 2.270 ;
        RECT  4.970 0.610 5.300 0.890 ;
        RECT  4.980 1.110 5.140 2.670 ;
        RECT  4.920 1.110 4.980 1.880 ;
        RECT  4.690 0.440 4.970 0.890 ;
        RECT  3.720 1.720 4.920 1.880 ;
        RECT  3.200 1.340 4.760 1.560 ;
        RECT  4.100 2.550 4.380 3.050 ;
        RECT  3.410 0.960 4.300 1.180 ;
        RECT  3.400 2.830 4.100 3.050 ;
        RECT  3.440 1.720 3.720 2.000 ;
        RECT  3.250 0.610 3.410 1.180 ;
        RECT  3.120 2.830 3.400 3.110 ;
        RECT  2.640 0.610 3.250 0.770 ;
        RECT  3.090 1.340 3.200 2.670 ;
        RECT  2.770 2.830 3.120 2.990 ;
        RECT  2.930 0.930 3.090 2.670 ;
        RECT  2.800 0.930 2.930 1.210 ;
        RECT  2.640 1.370 2.770 2.990 ;
        RECT  2.600 0.610 2.640 2.990 ;
        RECT  2.480 0.610 2.600 1.650 ;
        RECT  2.160 2.880 2.440 3.160 ;
        RECT  2.040 0.440 2.320 0.720 ;
        RECT  0.960 2.880 2.160 3.040 ;
        RECT  0.810 0.560 2.040 0.720 ;
        RECT  0.930 1.260 1.840 1.480 ;
        RECT  0.810 2.180 1.200 2.400 ;
        RECT  0.680 2.880 0.960 3.160 ;
        RECT  0.810 1.030 0.930 1.480 ;
        RECT  0.530 0.440 0.810 0.720 ;
        RECT  0.650 1.030 0.810 2.400 ;
        RECT  0.530 1.910 0.650 2.190 ;
    END
END SDFFQX2TR

MACRO SDFFQX1TR
    CLASS CORE ;
    FOREIGN SDFFQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.640 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.920 1.960 2.360 ;
        RECT  1.680 1.920 1.840 2.720 ;
        RECT  0.420 2.560 1.680 2.720 ;
        RECT  0.260 1.550 0.420 2.720 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.560 0.440 8.720 3.010 ;
        RECT  8.480 0.440 8.560 0.930 ;
        RECT  8.470 2.440 8.560 3.010 ;
        RECT  7.610 0.770 8.480 0.930 ;
        RECT  8.080 2.440 8.470 2.760 ;
        RECT  7.450 0.450 7.610 0.930 ;
        RECT  7.140 0.450 7.450 0.610 ;
        END
        ANTENNADIFFAREA 2.014 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.170 2.320 1.620 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 2.040 4.390 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.100 -0.280 8.800 0.280 ;
        RECT  7.820 -0.280 8.100 0.610 ;
        RECT  6.020 -0.280 7.820 0.280 ;
        RECT  5.740 -0.280 6.020 0.700 ;
        RECT  4.530 -0.280 5.740 0.280 ;
        RECT  3.760 -0.280 4.530 0.640 ;
        RECT  1.760 -0.280 3.760 0.280 ;
        RECT  1.480 -0.280 1.760 0.340 ;
        RECT  0.310 -0.280 1.480 0.280 ;
        RECT  0.150 -0.280 0.310 1.310 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.250 3.320 8.800 3.880 ;
        RECT  7.940 2.920 8.250 3.880 ;
        RECT  6.120 3.320 7.940 3.880 ;
        RECT  5.840 3.260 6.120 3.880 ;
        RECT  4.920 3.320 5.840 3.880 ;
        RECT  4.640 3.260 4.920 3.880 ;
        RECT  3.940 3.320 4.640 3.880 ;
        RECT  3.660 3.260 3.940 3.880 ;
        RECT  1.840 3.320 3.660 3.880 ;
        RECT  1.560 3.260 1.840 3.880 ;
        RECT  0.370 3.320 1.560 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.240 1.090 8.400 2.230 ;
        RECT  8.120 1.090 8.240 1.250 ;
        RECT  8.120 1.860 8.240 2.230 ;
        RECT  7.640 1.860 8.120 2.020 ;
        RECT  7.960 1.380 8.000 1.700 ;
        RECT  7.800 1.350 7.960 1.700 ;
        RECT  7.180 1.350 7.800 1.510 ;
        RECT  7.380 1.680 7.640 2.020 ;
        RECT  7.180 2.880 7.240 3.160 ;
        RECT  7.020 1.090 7.180 3.160 ;
        RECT  6.780 1.090 7.020 1.250 ;
        RECT  6.780 0.550 6.940 0.890 ;
        RECT  6.700 1.500 6.860 2.990 ;
        RECT  6.620 0.730 6.780 0.890 ;
        RECT  6.620 1.500 6.700 1.780 ;
        RECT  4.400 2.830 6.700 2.990 ;
        RECT  6.460 0.730 6.620 1.780 ;
        RECT  6.380 2.110 6.540 2.570 ;
        RECT  6.060 1.500 6.460 1.780 ;
        RECT  5.900 2.110 6.380 2.270 ;
        RECT  6.140 1.000 6.300 1.310 ;
        RECT  5.900 1.150 6.140 1.310 ;
        RECT  5.740 1.150 5.900 2.670 ;
        RECT  5.200 2.510 5.740 2.670 ;
        RECT  5.420 0.690 5.580 2.270 ;
        RECT  5.330 0.690 5.420 0.910 ;
        RECT  5.150 0.440 5.330 0.910 ;
        RECT  5.200 1.110 5.260 1.880 ;
        RECT  5.100 1.110 5.200 2.670 ;
        RECT  4.810 0.440 5.150 0.660 ;
        RECT  5.040 1.720 5.100 2.670 ;
        RECT  3.740 1.720 5.040 1.880 ;
        RECT  3.120 1.400 4.930 1.560 ;
        RECT  3.430 1.020 4.420 1.180 ;
        RECT  4.120 2.520 4.400 2.990 ;
        RECT  3.350 2.830 4.120 2.990 ;
        RECT  3.460 1.720 3.740 1.940 ;
        RECT  3.270 0.610 3.430 1.180 ;
        RECT  3.070 2.830 3.350 3.110 ;
        RECT  2.670 0.610 3.270 0.770 ;
        RECT  3.120 2.390 3.180 2.670 ;
        RECT  3.110 1.400 3.120 2.670 ;
        RECT  2.960 0.930 3.110 2.670 ;
        RECT  2.800 2.830 3.070 2.990 ;
        RECT  2.950 0.930 2.960 1.560 ;
        RECT  2.830 0.930 2.950 1.210 ;
        RECT  2.790 1.720 2.800 2.990 ;
        RECT  2.670 1.380 2.790 2.990 ;
        RECT  2.640 0.610 2.670 2.990 ;
        RECT  2.510 0.610 2.640 1.880 ;
        RECT  2.200 2.880 2.480 3.140 ;
        RECT  2.070 0.480 2.350 0.720 ;
        RECT  0.900 2.880 2.200 3.040 ;
        RECT  0.800 0.560 2.070 0.720 ;
        RECT  0.930 1.260 1.880 1.480 ;
        RECT  0.870 2.230 1.200 2.390 ;
        RECT  0.870 1.030 0.930 1.480 ;
        RECT  0.680 2.880 0.900 3.160 ;
        RECT  0.710 1.030 0.870 2.390 ;
        RECT  0.640 0.440 0.800 0.720 ;
        RECT  0.590 1.910 0.710 2.190 ;
    END
END SDFFQX1TR

MACRO SDFFNSRXLTR
    CLASS CORE ;
    FOREIGN SDFFNSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 2.440 9.520 2.800 ;
        RECT  8.860 2.520 9.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.540 2.320 1.960 ;
        RECT  1.460 1.540 2.080 1.820 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.410 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 1.030 11.520 2.360 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 2.040 10.720 2.360 ;
        RECT  10.260 1.030 10.420 2.360 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.140 1.680 1.300 ;
        RECT  1.300 2.040 1.520 2.480 ;
        RECT  1.140 1.140 1.300 2.480 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.470 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.040 -0.280 11.600 0.280 ;
        RECT  10.760 -0.280 11.040 0.520 ;
        RECT  9.470 -0.280 10.760 0.280 ;
        RECT  9.190 -0.280 9.470 1.140 ;
        RECT  5.580 -0.280 9.190 0.280 ;
        RECT  4.740 -0.280 5.580 0.290 ;
        RECT  3.780 -0.280 4.740 0.280 ;
        RECT  3.500 -0.280 3.780 0.290 ;
        RECT  1.540 -0.280 3.500 0.280 ;
        RECT  1.380 -0.280 1.540 0.340 ;
        RECT  0.340 -0.280 1.380 0.280 ;
        RECT  0.180 -0.280 0.340 1.310 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.000 3.320 11.600 3.880 ;
        RECT  10.720 3.260 11.000 3.880 ;
        RECT  9.460 3.320 10.720 3.880 ;
        RECT  9.180 3.200 9.460 3.880 ;
        RECT  7.420 3.320 9.180 3.880 ;
        RECT  7.140 2.930 7.420 3.880 ;
        RECT  5.900 3.320 7.140 3.880 ;
        RECT  4.870 2.890 5.900 3.880 ;
        RECT  3.780 3.320 4.870 3.880 ;
        RECT  3.500 3.150 3.780 3.880 ;
        RECT  1.620 3.320 3.500 3.880 ;
        RECT  1.340 3.200 1.620 3.880 ;
        RECT  0.440 3.320 1.340 3.880 ;
        RECT  0.160 3.200 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.960 0.680 11.120 2.930 ;
        RECT  10.440 0.680 10.960 0.840 ;
        RECT  10.140 2.770 10.960 2.930 ;
        RECT  10.160 0.510 10.440 0.840 ;
        RECT  9.940 1.000 10.100 1.920 ;
        RECT  9.740 1.000 9.940 1.160 ;
        RECT  9.920 1.760 9.940 1.920 ;
        RECT  9.760 1.760 9.920 2.190 ;
        RECT  8.560 1.760 9.760 1.920 ;
        RECT  9.480 1.320 9.640 1.600 ;
        RECT  8.560 1.320 9.480 1.480 ;
        RECT  8.820 0.470 8.880 0.750 ;
        RECT  8.580 2.080 8.860 2.360 ;
        RECT  8.720 0.450 8.820 0.750 ;
        RECT  6.400 0.450 8.720 0.610 ;
        RECT  8.560 2.200 8.580 2.360 ;
        RECT  8.400 1.210 8.560 1.480 ;
        RECT  8.400 1.640 8.560 1.920 ;
        RECT  8.400 2.200 8.560 2.770 ;
        RECT  7.920 1.210 8.400 1.370 ;
        RECT  6.140 2.610 8.400 2.770 ;
        RECT  8.080 0.770 8.240 1.050 ;
        RECT  8.080 1.530 8.240 2.450 ;
        RECT  7.480 0.770 8.080 0.930 ;
        RECT  7.960 1.530 8.080 1.810 ;
        RECT  5.760 2.290 8.080 2.450 ;
        RECT  7.800 1.090 7.920 1.370 ;
        RECT  7.800 1.970 7.920 2.130 ;
        RECT  7.640 1.090 7.800 2.130 ;
        RECT  7.320 0.770 7.480 2.130 ;
        RECT  6.720 0.770 7.320 0.930 ;
        RECT  7.200 1.850 7.320 2.130 ;
        RECT  7.040 1.090 7.160 1.310 ;
        RECT  6.880 1.090 7.040 2.130 ;
        RECT  6.660 1.620 6.880 2.130 ;
        RECT  6.560 0.770 6.720 1.460 ;
        RECT  5.760 1.620 6.660 1.780 ;
        RECT  6.080 1.300 6.560 1.460 ;
        RECT  6.240 0.450 6.400 1.140 ;
        RECT  5.440 1.940 6.230 2.100 ;
        RECT  5.920 0.450 6.080 1.460 ;
        RECT  2.640 0.450 5.920 0.610 ;
        RECT  5.600 0.770 5.760 1.780 ;
        RECT  5.600 2.290 5.760 2.540 ;
        RECT  3.600 0.770 5.600 0.930 ;
        RECT  5.090 2.380 5.600 2.540 ;
        RECT  5.280 1.090 5.440 2.220 ;
        RECT  5.080 1.090 5.280 1.250 ;
        RECT  4.930 2.120 5.090 2.540 ;
        RECT  3.920 2.120 4.930 2.280 ;
        RECT  4.470 2.450 4.710 3.160 ;
        RECT  2.960 2.450 4.470 2.610 ;
        RECT  3.920 1.090 4.460 1.310 ;
        RECT  4.020 2.770 4.300 3.050 ;
        RECT  3.260 2.770 4.020 2.930 ;
        RECT  3.760 1.090 3.920 2.280 ;
        RECT  3.340 2.120 3.760 2.280 ;
        RECT  3.440 0.770 3.600 1.310 ;
        RECT  3.120 1.550 3.340 2.280 ;
        RECT  2.980 2.770 3.260 3.050 ;
        RECT  2.640 2.770 2.980 2.930 ;
        RECT  2.800 0.780 2.960 2.610 ;
        RECT  2.480 0.450 2.640 2.930 ;
        RECT  2.160 0.500 2.320 0.930 ;
        RECT  2.100 2.370 2.320 2.810 ;
        RECT  0.660 0.500 2.160 0.660 ;
        RECT  2.000 1.090 2.140 1.250 ;
        RECT  0.760 2.650 2.100 2.810 ;
        RECT  1.840 0.820 2.000 1.250 ;
        RECT  0.980 0.820 1.840 0.980 ;
        RECT  0.820 0.820 0.980 2.190 ;
        RECT  0.660 2.530 0.760 2.810 ;
        RECT  0.500 0.440 0.660 2.810 ;
    END
END SDFFNSRXLTR

MACRO SDFFNSRX4TR
    CLASS CORE ;
    FOREIGN SDFFNSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.760 2.440 9.120 2.760 ;
        RECT  8.600 2.440 8.760 3.160 ;
        RECT  8.460 3.000 8.600 3.160 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.540 2.320 1.960 ;
        RECT  1.460 1.540 2.080 1.820 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.410 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.840 1.040 11.920 1.760 ;
        RECT  11.600 0.600 11.840 3.130 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.650 1.090 10.870 2.360 ;
        RECT  10.590 1.090 10.650 2.160 ;
        RECT  10.480 1.440 10.590 2.160 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.140 1.680 1.300 ;
        RECT  1.300 2.040 1.520 2.480 ;
        RECT  1.140 1.140 1.300 2.480 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.470 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 -0.280 12.400 0.280 ;
        RECT  12.080 -0.280 12.310 1.110 ;
        RECT  12.030 -0.280 12.080 0.710 ;
        RECT  11.350 -0.280 12.030 0.280 ;
        RECT  11.070 -0.280 11.350 0.610 ;
        RECT  10.390 -0.280 11.070 0.280 ;
        RECT  10.110 -0.280 10.390 0.610 ;
        RECT  9.450 -0.280 10.110 0.280 ;
        RECT  9.170 -0.280 9.450 0.400 ;
        RECT  5.420 -0.280 9.170 0.280 ;
        RECT  4.740 -0.280 5.420 0.290 ;
        RECT  3.780 -0.280 4.740 0.280 ;
        RECT  3.500 -0.280 3.780 0.290 ;
        RECT  1.540 -0.280 3.500 0.280 ;
        RECT  1.380 -0.280 1.540 0.340 ;
        RECT  0.340 -0.280 1.380 0.280 ;
        RECT  0.180 -0.280 0.340 1.310 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.310 3.320 12.400 3.880 ;
        RECT  12.030 2.430 12.310 3.880 ;
        RECT  11.350 3.320 12.030 3.880 ;
        RECT  11.070 2.840 11.350 3.880 ;
        RECT  10.390 3.320 11.070 3.880 ;
        RECT  10.110 2.840 10.390 3.880 ;
        RECT  9.260 3.320 10.110 3.880 ;
        RECT  8.980 3.200 9.260 3.880 ;
        RECT  7.420 3.320 8.980 3.880 ;
        RECT  7.140 2.990 7.420 3.880 ;
        RECT  5.900 3.320 7.140 3.880 ;
        RECT  4.870 2.890 5.900 3.880 ;
        RECT  3.780 3.320 4.870 3.880 ;
        RECT  3.500 3.150 3.780 3.880 ;
        RECT  1.620 3.320 3.500 3.880 ;
        RECT  1.340 3.200 1.620 3.880 ;
        RECT  0.440 3.320 1.340 3.880 ;
        RECT  0.160 3.200 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.190 1.350 11.440 1.640 ;
        RECT  11.030 0.770 11.190 2.680 ;
        RECT  9.910 0.770 11.030 0.930 ;
        RECT  9.910 2.520 11.030 2.680 ;
        RECT  10.160 1.090 10.320 2.170 ;
        RECT  9.570 1.090 10.160 1.370 ;
        RECT  9.710 2.010 10.160 2.170 ;
        RECT  9.630 0.450 9.910 0.930 ;
        RECT  9.630 2.520 9.910 3.150 ;
        RECT  9.430 2.010 9.710 2.290 ;
        RECT  9.050 1.560 9.570 1.850 ;
        RECT  8.620 2.010 9.430 2.170 ;
        RECT  8.880 1.210 9.050 1.850 ;
        RECT  8.630 0.450 8.910 0.750 ;
        RECT  7.860 1.210 8.880 1.370 ;
        RECT  6.400 0.450 8.630 0.610 ;
        RECT  8.400 1.640 8.620 2.170 ;
        RECT  6.420 2.670 8.400 2.830 ;
        RECT  8.080 1.530 8.240 2.510 ;
        RECT  8.050 0.770 8.210 1.050 ;
        RECT  7.960 1.530 8.080 1.810 ;
        RECT  6.740 2.350 8.080 2.510 ;
        RECT  7.480 0.770 8.050 0.930 ;
        RECT  7.800 1.970 7.920 2.190 ;
        RECT  7.800 1.090 7.860 1.370 ;
        RECT  7.640 1.090 7.800 2.190 ;
        RECT  7.320 0.770 7.480 2.170 ;
        RECT  6.720 0.770 7.320 0.930 ;
        RECT  7.200 1.890 7.320 2.170 ;
        RECT  7.040 1.090 7.160 1.310 ;
        RECT  6.880 1.090 7.040 2.130 ;
        RECT  6.660 1.620 6.880 2.130 ;
        RECT  6.580 2.290 6.740 2.510 ;
        RECT  6.560 0.770 6.720 1.460 ;
        RECT  5.760 1.620 6.660 1.780 ;
        RECT  5.760 2.290 6.580 2.450 ;
        RECT  6.080 1.300 6.560 1.460 ;
        RECT  6.140 2.610 6.420 2.830 ;
        RECT  6.240 0.450 6.400 1.140 ;
        RECT  5.440 1.940 6.230 2.100 ;
        RECT  5.920 0.450 6.080 1.460 ;
        RECT  2.640 0.450 5.920 0.610 ;
        RECT  5.600 0.770 5.760 1.780 ;
        RECT  5.600 2.290 5.760 2.540 ;
        RECT  3.600 0.770 5.600 0.930 ;
        RECT  5.090 2.380 5.600 2.540 ;
        RECT  5.280 1.090 5.440 2.220 ;
        RECT  5.080 1.090 5.280 1.250 ;
        RECT  4.930 2.120 5.090 2.540 ;
        RECT  3.920 2.120 4.930 2.280 ;
        RECT  4.470 2.450 4.710 3.160 ;
        RECT  2.960 2.450 4.470 2.610 ;
        RECT  3.920 1.090 4.340 1.310 ;
        RECT  4.020 2.770 4.300 3.050 ;
        RECT  3.260 2.770 4.020 2.930 ;
        RECT  3.760 1.090 3.920 2.280 ;
        RECT  3.340 2.120 3.760 2.280 ;
        RECT  3.440 0.770 3.600 1.310 ;
        RECT  3.120 1.550 3.340 2.280 ;
        RECT  2.980 2.770 3.260 3.050 ;
        RECT  2.640 2.770 2.980 2.930 ;
        RECT  2.800 0.780 2.960 2.610 ;
        RECT  2.480 0.450 2.640 2.930 ;
        RECT  2.160 0.500 2.320 0.930 ;
        RECT  2.100 2.370 2.320 2.810 ;
        RECT  0.660 0.500 2.160 0.660 ;
        RECT  2.000 1.090 2.140 1.250 ;
        RECT  0.760 2.650 2.100 2.810 ;
        RECT  1.840 0.820 2.000 1.250 ;
        RECT  0.980 0.820 1.840 0.980 ;
        RECT  0.820 0.820 0.980 2.190 ;
        RECT  0.660 2.530 0.760 2.810 ;
        RECT  0.500 0.440 0.660 2.810 ;
    END
END SDFFNSRX4TR

MACRO SDFFNSRX2TR
    CLASS CORE ;
    FOREIGN SDFFNSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 2.440 9.520 2.800 ;
        RECT  8.860 2.520 9.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.540 2.320 1.960 ;
        RECT  1.460 1.540 2.080 1.820 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.410 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 0.520 11.520 3.110 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 2.040 10.720 2.720 ;
        RECT  10.420 1.090 10.550 1.310 ;
        RECT  10.250 1.090 10.420 2.720 ;
        END
        ANTENNADIFFAREA 3.272 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.140 1.680 1.300 ;
        RECT  1.300 2.040 1.520 2.480 ;
        RECT  1.140 1.140 1.300 2.480 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.470 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.030 -0.280 11.600 0.280 ;
        RECT  10.750 -0.280 11.030 0.610 ;
        RECT  9.450 -0.280 10.750 0.280 ;
        RECT  9.170 -0.280 9.450 0.400 ;
        RECT  3.780 -0.280 9.170 0.280 ;
        RECT  3.500 -0.280 3.780 0.290 ;
        RECT  1.540 -0.280 3.500 0.280 ;
        RECT  1.380 -0.280 1.540 0.340 ;
        RECT  0.340 -0.280 1.380 0.280 ;
        RECT  0.180 -0.280 0.340 1.310 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.990 3.320 11.600 3.880 ;
        RECT  10.710 3.260 10.990 3.880 ;
        RECT  9.460 3.320 10.710 3.880 ;
        RECT  9.180 3.200 9.460 3.880 ;
        RECT  7.420 3.320 9.180 3.880 ;
        RECT  7.140 2.990 7.420 3.880 ;
        RECT  5.900 3.320 7.140 3.880 ;
        RECT  4.870 2.890 5.900 3.880 ;
        RECT  3.780 3.320 4.870 3.880 ;
        RECT  3.500 3.150 3.780 3.880 ;
        RECT  1.620 3.320 3.500 3.880 ;
        RECT  1.340 3.200 1.620 3.880 ;
        RECT  0.440 3.320 1.340 3.880 ;
        RECT  0.160 3.200 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.960 0.770 11.120 3.100 ;
        RECT  10.210 0.770 10.960 0.930 ;
        RECT  10.900 1.350 10.960 1.640 ;
        RECT  9.980 2.940 10.960 3.100 ;
        RECT  9.930 0.450 10.210 0.930 ;
        RECT  9.930 1.090 10.090 1.950 ;
        RECT  9.700 2.940 9.980 3.150 ;
        RECT  9.640 1.090 9.930 1.310 ;
        RECT  9.920 1.790 9.930 1.950 ;
        RECT  9.760 1.790 9.920 2.190 ;
        RECT  8.560 1.790 9.760 1.950 ;
        RECT  8.930 1.470 9.580 1.630 ;
        RECT  8.760 1.320 8.930 1.630 ;
        RECT  8.630 0.450 8.910 0.750 ;
        RECT  8.580 2.110 8.860 2.360 ;
        RECT  8.560 1.320 8.760 1.480 ;
        RECT  6.400 0.450 8.630 0.610 ;
        RECT  8.560 2.200 8.580 2.360 ;
        RECT  8.400 1.210 8.560 1.480 ;
        RECT  8.400 1.640 8.560 1.950 ;
        RECT  8.400 2.200 8.560 2.830 ;
        RECT  7.860 1.210 8.400 1.370 ;
        RECT  6.420 2.670 8.400 2.830 ;
        RECT  8.080 1.530 8.240 2.510 ;
        RECT  8.050 0.770 8.210 1.050 ;
        RECT  7.960 1.530 8.080 1.810 ;
        RECT  6.740 2.350 8.080 2.510 ;
        RECT  7.480 0.770 8.050 0.930 ;
        RECT  7.800 1.970 7.920 2.190 ;
        RECT  7.800 1.090 7.860 1.370 ;
        RECT  7.640 1.090 7.800 2.190 ;
        RECT  7.320 0.770 7.480 2.190 ;
        RECT  6.720 0.770 7.320 0.930 ;
        RECT  7.200 1.910 7.320 2.190 ;
        RECT  7.040 1.090 7.160 1.310 ;
        RECT  6.880 1.090 7.040 2.130 ;
        RECT  6.660 1.620 6.880 2.130 ;
        RECT  6.580 2.290 6.740 2.510 ;
        RECT  6.560 0.770 6.720 1.460 ;
        RECT  5.760 1.620 6.660 1.780 ;
        RECT  5.760 2.290 6.580 2.450 ;
        RECT  6.080 1.300 6.560 1.460 ;
        RECT  6.140 2.610 6.420 2.830 ;
        RECT  6.240 0.450 6.400 1.140 ;
        RECT  5.440 1.940 6.230 2.100 ;
        RECT  5.920 0.450 6.080 1.460 ;
        RECT  2.640 0.450 5.920 0.610 ;
        RECT  5.600 0.770 5.760 1.780 ;
        RECT  5.600 2.290 5.760 2.540 ;
        RECT  3.600 0.770 5.600 0.930 ;
        RECT  5.090 2.380 5.600 2.540 ;
        RECT  5.280 1.090 5.440 2.220 ;
        RECT  5.080 1.090 5.280 1.250 ;
        RECT  4.930 2.120 5.090 2.540 ;
        RECT  3.920 2.120 4.930 2.280 ;
        RECT  4.470 2.450 4.710 3.160 ;
        RECT  2.960 2.450 4.470 2.610 ;
        RECT  3.920 1.090 4.340 1.310 ;
        RECT  4.020 2.770 4.300 3.050 ;
        RECT  3.260 2.770 4.020 2.930 ;
        RECT  3.760 1.090 3.920 2.280 ;
        RECT  3.340 2.120 3.760 2.280 ;
        RECT  3.440 0.770 3.600 1.310 ;
        RECT  3.120 1.550 3.340 2.280 ;
        RECT  2.980 2.770 3.260 3.050 ;
        RECT  2.640 2.770 2.980 2.930 ;
        RECT  2.800 0.780 2.960 2.610 ;
        RECT  2.480 0.450 2.640 2.930 ;
        RECT  2.160 0.500 2.320 0.930 ;
        RECT  2.100 2.370 2.320 2.810 ;
        RECT  0.660 0.500 2.160 0.660 ;
        RECT  2.000 1.090 2.140 1.250 ;
        RECT  0.760 2.650 2.100 2.810 ;
        RECT  1.840 0.820 2.000 1.250 ;
        RECT  0.980 0.820 1.840 0.980 ;
        RECT  0.820 0.820 0.980 2.190 ;
        RECT  0.660 2.530 0.760 2.810 ;
        RECT  0.500 0.440 0.660 2.810 ;
    END
END SDFFNSRX2TR

MACRO SDFFNSRX1TR
    CLASS CORE ;
    FOREIGN SDFFNSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 2.440 9.520 2.800 ;
        RECT  8.860 2.520 9.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.540 2.320 1.960 ;
        RECT  1.460 1.540 2.080 1.820 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.410 5.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.280 1.030 11.520 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 2.040 10.720 2.360 ;
        RECT  10.260 1.030 10.420 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.140 1.680 1.300 ;
        RECT  1.300 2.040 1.520 2.480 ;
        RECT  1.140 1.140 1.300 2.480 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.470 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.000 -0.280 11.600 0.280 ;
        RECT  10.720 -0.280 11.000 0.340 ;
        RECT  9.470 -0.280 10.720 0.280 ;
        RECT  9.190 -0.280 9.470 1.140 ;
        RECT  3.780 -0.280 9.190 0.280 ;
        RECT  3.500 -0.280 3.780 0.290 ;
        RECT  1.540 -0.280 3.500 0.280 ;
        RECT  1.380 -0.280 1.540 0.340 ;
        RECT  0.340 -0.280 1.380 0.280 ;
        RECT  0.120 -0.280 0.340 1.310 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.000 3.320 11.600 3.880 ;
        RECT  10.720 3.260 11.000 3.880 ;
        RECT  9.460 3.320 10.720 3.880 ;
        RECT  9.180 3.200 9.460 3.880 ;
        RECT  7.420 3.320 9.180 3.880 ;
        RECT  7.140 2.930 7.420 3.880 ;
        RECT  5.900 3.320 7.140 3.880 ;
        RECT  4.870 2.890 5.900 3.880 ;
        RECT  3.780 3.320 4.870 3.880 ;
        RECT  3.500 3.150 3.780 3.880 ;
        RECT  1.620 3.320 3.500 3.880 ;
        RECT  1.340 3.200 1.620 3.880 ;
        RECT  0.440 3.320 1.340 3.880 ;
        RECT  0.160 3.200 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.960 0.500 11.120 3.070 ;
        RECT  10.440 0.500 10.960 0.660 ;
        RECT  10.420 2.910 10.960 3.070 ;
        RECT  10.160 0.450 10.440 0.660 ;
        RECT  10.110 2.910 10.420 3.130 ;
        RECT  9.940 1.000 10.100 1.920 ;
        RECT  9.740 1.000 9.940 1.160 ;
        RECT  9.920 1.760 9.940 1.920 ;
        RECT  9.760 1.760 9.920 2.190 ;
        RECT  8.560 1.760 9.760 1.920 ;
        RECT  9.480 1.320 9.640 1.600 ;
        RECT  8.560 1.320 9.480 1.480 ;
        RECT  8.820 0.470 8.880 0.750 ;
        RECT  8.580 2.080 8.860 2.360 ;
        RECT  8.720 0.450 8.820 0.750 ;
        RECT  6.400 0.450 8.720 0.610 ;
        RECT  8.560 2.200 8.580 2.360 ;
        RECT  8.400 1.210 8.560 1.480 ;
        RECT  8.400 1.640 8.560 1.920 ;
        RECT  8.400 2.200 8.560 2.770 ;
        RECT  7.920 1.210 8.400 1.370 ;
        RECT  6.140 2.610 8.400 2.770 ;
        RECT  8.080 0.770 8.240 1.050 ;
        RECT  8.080 1.530 8.240 2.450 ;
        RECT  7.480 0.770 8.080 0.930 ;
        RECT  7.960 1.530 8.080 1.810 ;
        RECT  5.760 2.290 8.080 2.450 ;
        RECT  7.800 1.090 7.920 1.370 ;
        RECT  7.800 1.970 7.920 2.130 ;
        RECT  7.640 1.090 7.800 2.130 ;
        RECT  7.320 0.770 7.480 2.130 ;
        RECT  6.720 0.770 7.320 0.930 ;
        RECT  7.200 1.850 7.320 2.130 ;
        RECT  7.040 1.090 7.160 1.310 ;
        RECT  6.880 1.090 7.040 2.130 ;
        RECT  6.660 1.620 6.880 2.130 ;
        RECT  6.560 0.770 6.720 1.460 ;
        RECT  5.760 1.620 6.660 1.780 ;
        RECT  6.080 1.300 6.560 1.460 ;
        RECT  6.240 0.450 6.400 1.140 ;
        RECT  5.440 1.940 6.230 2.100 ;
        RECT  5.920 0.450 6.080 1.460 ;
        RECT  2.640 0.450 5.920 0.610 ;
        RECT  5.600 0.770 5.760 1.780 ;
        RECT  5.600 2.290 5.760 2.540 ;
        RECT  3.600 0.770 5.600 0.930 ;
        RECT  5.090 2.380 5.600 2.540 ;
        RECT  5.280 1.090 5.440 2.220 ;
        RECT  5.080 1.090 5.280 1.250 ;
        RECT  4.930 2.120 5.090 2.540 ;
        RECT  3.920 2.120 4.930 2.280 ;
        RECT  4.470 2.450 4.710 3.160 ;
        RECT  2.960 2.450 4.470 2.610 ;
        RECT  3.920 1.090 4.460 1.310 ;
        RECT  4.020 2.770 4.300 3.050 ;
        RECT  3.260 2.770 4.020 2.930 ;
        RECT  3.760 1.090 3.920 2.280 ;
        RECT  3.340 2.120 3.760 2.280 ;
        RECT  3.440 0.770 3.600 1.310 ;
        RECT  3.120 1.550 3.340 2.280 ;
        RECT  2.980 2.770 3.260 3.050 ;
        RECT  2.640 2.770 2.980 2.930 ;
        RECT  2.800 0.780 2.960 2.610 ;
        RECT  2.480 0.450 2.640 2.930 ;
        RECT  2.160 0.500 2.320 0.930 ;
        RECT  2.100 2.370 2.320 2.810 ;
        RECT  0.660 0.500 2.160 0.660 ;
        RECT  2.000 1.090 2.140 1.250 ;
        RECT  0.760 2.650 2.100 2.810 ;
        RECT  1.840 0.820 2.000 1.250 ;
        RECT  0.980 0.820 1.840 0.980 ;
        RECT  0.820 0.820 0.980 2.190 ;
        RECT  0.660 2.530 0.760 2.810 ;
        RECT  0.500 0.440 0.660 2.810 ;
    END
END SDFFNSRX1TR

MACRO SDFFHQX8TR
    CLASS CORE ;
    FOREIGN SDFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 1.640 6.320 1.960 ;
        RECT  5.950 1.270 6.110 1.960 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.120 1.560 ;
        RECT  2.840 1.400 2.880 1.560 ;
        RECT  2.550 1.400 2.840 1.790 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.950 0.620 16.220 3.090 ;
        RECT  15.230 1.440 15.950 2.160 ;
        RECT  15.230 0.580 15.240 1.140 ;
        RECT  14.950 0.580 15.230 3.100 ;
        END
        ANTENNADIFFAREA 8.612 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.510 3.520 2.090 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.340 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.700 -0.280 16.800 0.280 ;
        RECT  16.430 -0.280 16.700 1.150 ;
        RECT  15.720 -0.280 16.430 0.280 ;
        RECT  15.440 -0.280 15.720 1.140 ;
        RECT  14.720 -0.280 15.440 0.280 ;
        RECT  14.020 -0.280 14.720 0.760 ;
        RECT  11.250 -0.280 14.020 0.280 ;
        RECT  10.970 -0.280 11.250 0.340 ;
        RECT  10.210 -0.280 10.970 0.280 ;
        RECT  9.930 -0.280 10.210 0.340 ;
        RECT  9.040 -0.280 9.930 0.280 ;
        RECT  8.760 -0.280 9.040 0.340 ;
        RECT  7.400 -0.280 8.760 0.280 ;
        RECT  7.240 -0.280 7.400 1.080 ;
        RECT  6.070 -0.280 7.240 0.280 ;
        RECT  7.030 0.800 7.240 1.080 ;
        RECT  5.360 -0.280 6.070 0.780 ;
        RECT  2.560 -0.280 5.360 0.280 ;
        RECT  2.280 -0.280 2.560 0.400 ;
        RECT  0.920 -0.280 2.280 0.280 ;
        RECT  0.620 -0.280 0.920 0.360 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.700 3.320 16.800 3.880 ;
        RECT  16.430 2.400 16.700 3.880 ;
        RECT  15.750 3.320 16.430 3.880 ;
        RECT  15.470 2.400 15.750 3.880 ;
        RECT  14.710 3.320 15.470 3.880 ;
        RECT  14.030 2.920 14.710 3.880 ;
        RECT  11.280 3.320 14.030 3.880 ;
        RECT  11.000 3.200 11.280 3.880 ;
        RECT  10.160 3.320 11.000 3.880 ;
        RECT  9.880 3.200 10.160 3.880 ;
        RECT  8.520 3.320 9.880 3.880 ;
        RECT  8.240 3.200 8.520 3.880 ;
        RECT  7.270 3.320 8.240 3.880 ;
        RECT  6.990 3.200 7.270 3.880 ;
        RECT  6.150 3.320 6.990 3.880 ;
        RECT  5.870 3.200 6.150 3.880 ;
        RECT  4.270 3.320 5.870 3.880 ;
        RECT  3.270 3.020 4.270 3.880 ;
        RECT  2.620 3.320 3.270 3.880 ;
        RECT  2.340 3.020 2.620 3.880 ;
        RECT  0.780 3.320 2.340 3.880 ;
        RECT  0.500 3.200 0.780 3.880 ;
        RECT  0.000 3.320 0.500 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  14.620 1.490 14.740 1.770 ;
        RECT  14.460 1.490 14.620 2.650 ;
        RECT  13.330 2.490 14.460 2.650 ;
        RECT  14.130 1.910 14.250 2.190 ;
        RECT  14.130 1.030 14.240 1.310 ;
        RECT  13.970 1.030 14.130 2.190 ;
        RECT  13.960 1.030 13.970 1.760 ;
        RECT  13.750 1.480 13.960 1.760 ;
        RECT  13.420 0.440 13.580 1.960 ;
        RECT  11.570 0.440 13.420 0.600 ;
        RECT  13.250 1.680 13.420 1.960 ;
        RECT  13.050 2.140 13.330 2.870 ;
        RECT  13.100 0.780 13.260 1.250 ;
        RECT  12.320 1.090 13.100 1.250 ;
        RECT  12.320 2.140 13.050 2.300 ;
        RECT  11.890 0.770 12.830 0.930 ;
        RECT  12.530 2.470 12.810 3.140 ;
        RECT  11.840 2.980 12.530 3.140 ;
        RECT  12.290 1.090 12.320 2.300 ;
        RECT  12.160 1.090 12.290 2.810 ;
        RECT  12.050 1.090 12.160 1.310 ;
        RECT  12.010 2.140 12.160 2.810 ;
        RECT  11.840 0.770 11.890 0.990 ;
        RECT  11.730 0.770 11.840 3.140 ;
        RECT  11.680 0.830 11.730 3.140 ;
        RECT  11.470 0.830 11.680 1.300 ;
        RECT  11.490 2.300 11.680 2.940 ;
        RECT  11.410 0.440 11.570 0.670 ;
        RECT  10.900 0.830 11.470 0.990 ;
        RECT  11.300 1.790 11.460 2.070 ;
        RECT  7.720 0.510 11.410 0.670 ;
        RECT  11.260 1.910 11.300 2.070 ;
        RECT  11.100 1.910 11.260 3.040 ;
        RECT  7.160 2.880 11.100 3.040 ;
        RECT  10.740 0.830 10.900 2.170 ;
        RECT  10.450 0.830 10.740 1.170 ;
        RECT  10.720 1.990 10.740 2.170 ;
        RECT  10.440 1.990 10.720 2.630 ;
        RECT  10.260 1.510 10.570 1.790 ;
        RECT  9.920 1.990 10.440 2.150 ;
        RECT  10.100 1.010 10.260 1.670 ;
        RECT  9.400 1.010 10.100 1.170 ;
        RECT  9.760 1.470 9.920 2.150 ;
        RECT  9.640 1.470 9.760 1.750 ;
        RECT  9.130 0.890 9.400 1.170 ;
        RECT  9.130 2.370 9.400 2.650 ;
        RECT  9.120 0.890 9.130 2.650 ;
        RECT  8.970 0.920 9.120 2.650 ;
        RECT  7.880 0.920 8.970 1.080 ;
        RECT  7.640 2.490 8.970 2.650 ;
        RECT  8.180 1.910 8.300 2.190 ;
        RECT  8.020 1.250 8.180 2.190 ;
        RECT  7.720 1.250 8.020 1.410 ;
        RECT  7.560 0.510 7.720 1.410 ;
        RECT  7.360 2.430 7.640 2.710 ;
        RECT  6.830 1.250 7.560 1.410 ;
        RECT  7.210 1.580 7.490 1.860 ;
        RECT  7.160 1.700 7.210 1.860 ;
        RECT  7.000 1.700 7.160 3.040 ;
        RECT  6.390 0.470 7.070 0.630 ;
        RECT  5.550 2.880 7.000 3.040 ;
        RECT  6.710 0.860 6.830 1.410 ;
        RECT  6.550 0.860 6.710 2.660 ;
        RECT  6.490 2.120 6.550 2.660 ;
        RECT  6.480 2.380 6.490 2.660 ;
        RECT  2.050 2.380 6.480 2.540 ;
        RECT  6.230 0.470 6.390 1.100 ;
        RECT  5.790 0.940 6.230 1.100 ;
        RECT  5.630 0.940 5.790 2.180 ;
        RECT  4.610 0.940 5.630 1.110 ;
        RECT  5.110 2.020 5.630 2.180 ;
        RECT  5.390 2.700 5.550 3.040 ;
        RECT  5.310 1.360 5.470 1.850 ;
        RECT  1.700 2.700 5.390 2.860 ;
        RECT  4.170 1.360 5.310 1.520 ;
        RECT  3.840 2.000 4.870 2.160 ;
        RECT  4.330 0.810 4.610 1.110 ;
        RECT  2.880 0.440 4.540 0.600 ;
        RECT  4.010 0.770 4.170 1.520 ;
        RECT  3.200 0.770 4.010 0.930 ;
        RECT  3.680 1.090 3.840 2.220 ;
        RECT  3.460 1.090 3.680 1.250 ;
        RECT  3.040 0.770 3.200 1.080 ;
        RECT  2.370 0.920 3.040 1.080 ;
        RECT  2.370 2.040 2.970 2.200 ;
        RECT  2.720 0.440 2.880 0.750 ;
        RECT  0.780 0.590 2.720 0.750 ;
        RECT  2.210 0.920 2.370 2.200 ;
        RECT  2.190 0.920 2.210 1.100 ;
        RECT  1.890 1.880 2.050 2.540 ;
        RECT  1.340 1.880 1.890 2.050 ;
        RECT  1.540 2.440 1.700 2.860 ;
        RECT  1.420 2.440 1.540 2.730 ;
        RECT  1.180 0.960 1.460 1.240 ;
        RECT  1.110 2.440 1.420 2.600 ;
        RECT  1.110 1.080 1.180 1.240 ;
        RECT  0.950 1.080 1.110 2.600 ;
        RECT  0.620 0.590 0.780 1.090 ;
        RECT  0.320 0.930 0.620 1.090 ;
        RECT  0.160 0.930 0.320 2.560 ;
    END
END SDFFHQX8TR

MACRO SDFFHQX4TR
    CLASS CORE ;
    FOREIGN SDFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 1.640 6.320 1.960 ;
        RECT  5.950 1.270 6.110 1.960 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.120 1.560 ;
        RECT  2.840 1.400 2.880 1.560 ;
        RECT  2.550 1.400 2.840 1.790 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.340 1.440 15.520 2.160 ;
        RECT  15.230 0.580 15.340 2.160 ;
        RECT  15.060 0.580 15.230 3.100 ;
        RECT  14.950 1.460 15.060 3.100 ;
        END
        ANTENNADIFFAREA 4.46 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.510 3.520 2.090 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.340 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.860 -0.280 16.000 0.280 ;
        RECT  15.580 -0.280 15.860 1.070 ;
        RECT  14.830 -0.280 15.580 0.280 ;
        RECT  14.020 -0.280 14.830 0.760 ;
        RECT  11.250 -0.280 14.020 0.280 ;
        RECT  10.970 -0.280 11.250 0.340 ;
        RECT  10.210 -0.280 10.970 0.280 ;
        RECT  9.930 -0.280 10.210 0.340 ;
        RECT  9.040 -0.280 9.930 0.280 ;
        RECT  8.760 -0.280 9.040 0.340 ;
        RECT  7.400 -0.280 8.760 0.280 ;
        RECT  7.240 -0.280 7.400 1.080 ;
        RECT  6.070 -0.280 7.240 0.280 ;
        RECT  7.030 0.800 7.240 1.080 ;
        RECT  5.360 -0.280 6.070 0.780 ;
        RECT  2.560 -0.280 5.360 0.280 ;
        RECT  2.280 -0.280 2.560 0.400 ;
        RECT  0.920 -0.280 2.280 0.280 ;
        RECT  0.620 -0.280 0.920 0.360 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.750 3.320 16.000 3.880 ;
        RECT  15.470 2.400 15.750 3.880 ;
        RECT  14.710 3.320 15.470 3.880 ;
        RECT  14.030 2.930 14.710 3.880 ;
        RECT  11.280 3.320 14.030 3.880 ;
        RECT  11.000 3.200 11.280 3.880 ;
        RECT  10.160 3.320 11.000 3.880 ;
        RECT  9.880 3.200 10.160 3.880 ;
        RECT  8.520 3.320 9.880 3.880 ;
        RECT  8.240 3.200 8.520 3.880 ;
        RECT  7.270 3.320 8.240 3.880 ;
        RECT  6.990 3.200 7.270 3.880 ;
        RECT  6.150 3.320 6.990 3.880 ;
        RECT  5.870 3.200 6.150 3.880 ;
        RECT  4.270 3.320 5.870 3.880 ;
        RECT  3.270 3.020 4.270 3.880 ;
        RECT  2.620 3.320 3.270 3.880 ;
        RECT  2.340 3.020 2.620 3.880 ;
        RECT  0.780 3.320 2.340 3.880 ;
        RECT  0.500 3.200 0.780 3.880 ;
        RECT  0.000 3.320 0.500 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  14.620 1.490 14.740 1.770 ;
        RECT  14.460 1.490 14.620 2.650 ;
        RECT  13.330 2.490 14.460 2.650 ;
        RECT  14.130 1.910 14.250 2.190 ;
        RECT  14.130 1.030 14.240 1.310 ;
        RECT  13.970 1.030 14.130 2.190 ;
        RECT  13.960 1.030 13.970 1.760 ;
        RECT  13.750 1.480 13.960 1.760 ;
        RECT  13.420 0.440 13.580 1.960 ;
        RECT  11.570 0.440 13.420 0.600 ;
        RECT  13.250 1.680 13.420 1.960 ;
        RECT  13.050 2.140 13.330 2.870 ;
        RECT  13.100 0.780 13.260 1.250 ;
        RECT  12.320 1.090 13.100 1.250 ;
        RECT  12.320 2.140 13.050 2.300 ;
        RECT  11.890 0.770 12.830 0.930 ;
        RECT  12.530 2.470 12.810 3.140 ;
        RECT  11.840 2.980 12.530 3.140 ;
        RECT  12.290 1.090 12.320 2.300 ;
        RECT  12.160 1.090 12.290 2.810 ;
        RECT  12.050 1.090 12.160 1.310 ;
        RECT  12.010 2.140 12.160 2.810 ;
        RECT  11.840 0.770 11.890 0.990 ;
        RECT  11.730 0.770 11.840 3.140 ;
        RECT  11.680 0.830 11.730 3.140 ;
        RECT  11.470 0.830 11.680 1.300 ;
        RECT  11.490 2.300 11.680 2.940 ;
        RECT  11.410 0.440 11.570 0.670 ;
        RECT  10.900 0.830 11.470 0.990 ;
        RECT  11.300 1.790 11.460 2.070 ;
        RECT  7.720 0.510 11.410 0.670 ;
        RECT  11.260 1.910 11.300 2.070 ;
        RECT  11.100 1.910 11.260 3.040 ;
        RECT  7.160 2.880 11.100 3.040 ;
        RECT  10.740 0.830 10.900 2.170 ;
        RECT  10.450 0.830 10.740 1.170 ;
        RECT  10.720 1.990 10.740 2.170 ;
        RECT  10.440 1.990 10.720 2.630 ;
        RECT  10.260 1.510 10.570 1.790 ;
        RECT  9.920 1.990 10.440 2.150 ;
        RECT  10.100 1.010 10.260 1.790 ;
        RECT  9.400 1.010 10.100 1.170 ;
        RECT  9.760 1.470 9.920 2.150 ;
        RECT  9.640 1.470 9.760 1.750 ;
        RECT  9.130 0.890 9.400 1.170 ;
        RECT  9.130 2.370 9.400 2.650 ;
        RECT  9.120 0.890 9.130 2.650 ;
        RECT  8.970 0.920 9.120 2.650 ;
        RECT  7.880 0.920 8.970 1.080 ;
        RECT  7.640 2.490 8.970 2.650 ;
        RECT  8.180 1.910 8.300 2.190 ;
        RECT  8.020 1.250 8.180 2.190 ;
        RECT  7.720 1.250 8.020 1.410 ;
        RECT  7.560 0.510 7.720 1.410 ;
        RECT  7.360 2.430 7.640 2.710 ;
        RECT  6.830 1.250 7.560 1.410 ;
        RECT  7.210 1.580 7.490 1.860 ;
        RECT  7.160 1.700 7.210 1.860 ;
        RECT  7.000 1.700 7.160 3.040 ;
        RECT  6.390 0.470 7.070 0.630 ;
        RECT  5.550 2.880 7.000 3.040 ;
        RECT  6.710 0.860 6.830 1.410 ;
        RECT  6.550 0.860 6.710 2.660 ;
        RECT  6.490 2.120 6.550 2.660 ;
        RECT  6.480 2.380 6.490 2.660 ;
        RECT  2.050 2.380 6.480 2.540 ;
        RECT  6.230 0.470 6.390 1.100 ;
        RECT  5.790 0.940 6.230 1.100 ;
        RECT  5.630 0.940 5.790 2.180 ;
        RECT  4.610 0.940 5.630 1.110 ;
        RECT  5.110 2.020 5.630 2.180 ;
        RECT  5.390 2.700 5.550 3.040 ;
        RECT  5.310 1.360 5.470 1.850 ;
        RECT  1.700 2.700 5.390 2.860 ;
        RECT  4.170 1.360 5.310 1.520 ;
        RECT  3.840 2.000 4.870 2.160 ;
        RECT  4.330 0.810 4.610 1.110 ;
        RECT  2.880 0.440 4.540 0.600 ;
        RECT  4.010 0.770 4.170 1.520 ;
        RECT  3.200 0.770 4.010 0.930 ;
        RECT  3.680 1.090 3.840 2.220 ;
        RECT  3.460 1.090 3.680 1.250 ;
        RECT  3.040 0.770 3.200 1.080 ;
        RECT  2.370 0.920 3.040 1.080 ;
        RECT  2.370 2.040 2.970 2.200 ;
        RECT  2.720 0.440 2.880 0.750 ;
        RECT  0.780 0.590 2.720 0.750 ;
        RECT  2.210 0.920 2.370 2.200 ;
        RECT  2.190 0.920 2.210 1.100 ;
        RECT  1.890 1.880 2.050 2.540 ;
        RECT  1.340 1.880 1.890 2.050 ;
        RECT  1.540 2.440 1.700 2.860 ;
        RECT  1.420 2.440 1.540 2.730 ;
        RECT  1.180 0.960 1.460 1.240 ;
        RECT  1.110 2.440 1.420 2.600 ;
        RECT  1.110 1.080 1.180 1.240 ;
        RECT  0.950 1.080 1.110 2.600 ;
        RECT  0.620 0.590 0.780 1.090 ;
        RECT  0.320 0.930 0.620 1.090 ;
        RECT  0.160 0.930 0.320 2.560 ;
    END
END SDFFHQX4TR

MACRO SDFFHQX2TR
    CLASS CORE ;
    FOREIGN SDFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.310 1.240 4.720 1.620 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.440 1.960 2.760 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.110 0.840 11.120 1.960 ;
        RECT  10.830 0.440 11.110 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.300 2.520 1.580 ;
        RECT  2.080 1.240 2.360 1.580 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.216 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.630 -0.280 11.200 0.280 ;
        RECT  10.350 -0.280 10.630 1.270 ;
        RECT  9.610 -0.280 10.350 0.340 ;
        RECT  9.330 -0.280 9.610 1.260 ;
        RECT  7.570 -0.280 9.330 0.280 ;
        RECT  6.190 -0.280 7.570 0.340 ;
        RECT  4.430 -0.280 6.190 0.280 ;
        RECT  4.150 -0.280 4.430 0.740 ;
        RECT  2.540 -0.280 4.150 0.280 ;
        RECT  2.260 -0.280 2.540 0.290 ;
        RECT  0.380 -0.280 2.260 0.280 ;
        RECT  0.100 -0.280 0.380 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.630 3.320 11.200 3.880 ;
        RECT  9.950 2.930 10.630 3.880 ;
        RECT  7.750 3.260 9.950 3.880 ;
        RECT  7.470 3.200 7.750 3.880 ;
        RECT  6.950 3.320 7.470 3.880 ;
        RECT  6.670 3.200 6.950 3.880 ;
        RECT  5.270 3.260 6.670 3.880 ;
        RECT  4.990 3.200 5.270 3.880 ;
        RECT  4.410 3.320 4.990 3.880 ;
        RECT  4.130 3.200 4.410 3.880 ;
        RECT  2.210 3.260 4.130 3.880 ;
        RECT  1.990 2.930 2.210 3.880 ;
        RECT  0.700 3.320 1.990 3.880 ;
        RECT  0.420 2.710 0.700 3.880 ;
        RECT  0.000 3.320 0.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.510 1.540 10.630 1.820 ;
        RECT  10.350 1.540 10.510 2.660 ;
        RECT  9.170 2.500 10.350 2.660 ;
        RECT  10.070 1.910 10.190 2.190 ;
        RECT  9.910 1.030 10.070 2.190 ;
        RECT  9.790 1.030 9.910 1.710 ;
        RECT  9.710 1.430 9.790 1.710 ;
        RECT  9.330 1.420 9.490 2.340 ;
        RECT  8.890 1.420 9.330 1.580 ;
        RECT  9.050 2.380 9.170 2.660 ;
        RECT  8.890 1.740 9.050 2.660 ;
        RECT  8.730 0.440 8.890 1.580 ;
        RECT  8.570 1.740 8.890 1.900 ;
        RECT  8.210 2.500 8.890 2.660 ;
        RECT  8.210 2.820 8.890 3.100 ;
        RECT  7.890 0.440 8.730 0.660 ;
        RECT  8.410 2.060 8.690 2.340 ;
        RECT  8.410 0.990 8.570 1.900 ;
        RECT  8.290 0.990 8.410 1.270 ;
        RECT  8.090 2.060 8.410 2.220 ;
        RECT  7.930 2.380 8.210 2.660 ;
        RECT  6.550 2.880 8.210 3.040 ;
        RECT  7.930 0.940 8.090 2.220 ;
        RECT  7.810 0.940 7.930 1.220 ;
        RECT  7.350 2.050 7.930 2.220 ;
        RECT  7.730 0.440 7.890 0.720 ;
        RECT  7.650 1.420 7.770 1.700 ;
        RECT  5.740 0.560 7.730 0.720 ;
        RECT  7.490 1.080 7.650 1.700 ;
        RECT  6.810 1.080 7.490 1.240 ;
        RECT  7.070 2.050 7.350 2.720 ;
        RECT  6.730 2.050 7.070 2.210 ;
        RECT  6.530 0.940 6.810 1.240 ;
        RECT  6.570 1.410 6.730 2.210 ;
        RECT  6.450 1.410 6.570 1.660 ;
        RECT  6.270 2.720 6.550 3.040 ;
        RECT  5.990 1.080 6.530 1.240 ;
        RECT  2.530 2.880 6.270 3.040 ;
        RECT  5.990 2.050 6.110 2.720 ;
        RECT  5.830 1.080 5.990 2.720 ;
        RECT  5.310 1.080 5.830 1.270 ;
        RECT  5.580 0.560 5.740 0.920 ;
        RECT  5.130 0.760 5.580 0.920 ;
        RECT  5.130 1.700 5.510 1.980 ;
        RECT  4.750 0.440 5.420 0.600 ;
        RECT  5.070 0.760 5.130 1.980 ;
        RECT  4.930 0.760 5.070 2.260 ;
        RECT  4.910 0.760 4.930 2.380 ;
        RECT  4.810 2.100 4.910 2.380 ;
        RECT  4.650 2.100 4.810 2.700 ;
        RECT  4.590 0.440 4.750 1.080 ;
        RECT  2.850 2.540 4.650 2.700 ;
        RECT  4.150 0.920 4.590 1.080 ;
        RECT  3.990 0.920 4.150 2.320 ;
        RECT  2.860 0.440 3.990 0.600 ;
        RECT  3.490 0.920 3.990 1.200 ;
        RECT  3.430 2.160 3.990 2.320 ;
        RECT  3.550 1.360 3.830 1.960 ;
        RECT  3.310 1.360 3.550 1.520 ;
        RECT  3.150 0.770 3.310 1.520 ;
        RECT  3.010 1.680 3.230 2.320 ;
        RECT  1.880 0.770 3.150 0.930 ;
        RECT  2.970 1.680 3.010 1.840 ;
        RECT  2.810 1.090 2.970 1.840 ;
        RECT  2.700 0.440 2.860 0.610 ;
        RECT  2.690 2.000 2.850 2.700 ;
        RECT  2.690 1.090 2.810 1.310 ;
        RECT  0.700 0.450 2.700 0.610 ;
        RECT  2.600 2.000 2.690 2.160 ;
        RECT  2.440 1.740 2.600 2.160 ;
        RECT  2.370 2.320 2.530 3.040 ;
        RECT  1.800 1.740 2.440 1.900 ;
        RECT  2.280 2.320 2.370 2.480 ;
        RECT  2.120 2.060 2.280 2.480 ;
        RECT  1.360 2.060 2.120 2.280 ;
        RECT  1.720 0.770 1.880 1.140 ;
        RECT  1.520 1.600 1.800 1.900 ;
        RECT  1.040 0.770 1.720 0.930 ;
        RECT  1.040 2.930 1.650 3.150 ;
        RECT  1.360 1.090 1.460 1.310 ;
        RECT  1.200 1.090 1.360 2.280 ;
        RECT  0.880 0.770 1.040 3.150 ;
        RECT  0.540 0.450 0.700 1.270 ;
        RECT  0.250 0.990 0.540 1.270 ;
        RECT  0.250 2.120 0.370 2.400 ;
        RECT  0.090 0.990 0.250 2.400 ;
    END
END SDFFHQX2TR

MACRO SDFFHQX1TR
    CLASS CORE ;
    FOREIGN SDFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.310 1.240 4.720 1.620 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.440 1.960 2.760 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.110 0.840 11.120 1.960 ;
        RECT  10.830 0.840 11.110 2.650 ;
        END
        ANTENNADIFFAREA 1.92 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.520 1.580 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.630 -0.280 11.200 0.280 ;
        RECT  10.350 -0.280 10.630 1.270 ;
        RECT  9.610 -0.280 10.350 0.340 ;
        RECT  9.330 -0.280 9.610 1.260 ;
        RECT  7.570 -0.280 9.330 0.280 ;
        RECT  6.190 -0.280 7.570 0.340 ;
        RECT  4.430 -0.280 6.190 0.280 ;
        RECT  4.150 -0.280 4.430 0.740 ;
        RECT  2.540 -0.280 4.150 0.280 ;
        RECT  2.260 -0.280 2.540 0.290 ;
        RECT  0.380 -0.280 2.260 0.280 ;
        RECT  0.100 -0.280 0.380 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.590 3.320 11.200 3.880 ;
        RECT  9.910 2.960 10.590 3.880 ;
        RECT  6.990 3.320 9.910 3.880 ;
        RECT  6.710 3.260 6.990 3.880 ;
        RECT  5.270 3.320 6.710 3.880 ;
        RECT  4.990 3.260 5.270 3.880 ;
        RECT  4.410 3.320 4.990 3.880 ;
        RECT  2.210 3.260 4.410 3.880 ;
        RECT  1.920 2.930 2.210 3.880 ;
        RECT  0.700 3.320 1.920 3.880 ;
        RECT  0.420 2.650 0.700 3.880 ;
        RECT  0.000 3.320 0.420 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.510 1.510 10.630 1.820 ;
        RECT  10.350 1.510 10.510 2.800 ;
        RECT  9.110 2.640 10.350 2.800 ;
        RECT  10.070 1.910 10.190 2.190 ;
        RECT  9.910 1.030 10.070 2.190 ;
        RECT  9.790 1.030 9.910 1.780 ;
        RECT  9.650 1.430 9.790 1.780 ;
        RECT  9.270 1.420 9.490 2.340 ;
        RECT  8.890 1.420 9.270 1.580 ;
        RECT  8.950 1.740 9.110 2.800 ;
        RECT  8.570 1.740 8.950 1.900 ;
        RECT  8.150 2.640 8.950 2.800 ;
        RECT  8.730 0.440 8.890 1.580 ;
        RECT  7.770 2.960 8.750 3.120 ;
        RECT  7.890 0.440 8.730 0.660 ;
        RECT  8.410 2.060 8.690 2.470 ;
        RECT  8.410 0.990 8.570 1.900 ;
        RECT  8.290 0.990 8.410 1.270 ;
        RECT  8.090 2.060 8.410 2.220 ;
        RECT  7.930 2.410 8.150 2.800 ;
        RECT  7.930 0.940 8.090 2.220 ;
        RECT  7.810 0.940 7.930 1.220 ;
        RECT  7.510 2.050 7.930 2.220 ;
        RECT  7.730 0.440 7.890 0.720 ;
        RECT  7.650 1.560 7.770 1.860 ;
        RECT  7.470 2.900 7.770 3.120 ;
        RECT  6.280 0.560 7.730 0.720 ;
        RECT  7.490 1.080 7.650 1.860 ;
        RECT  7.230 2.050 7.510 2.530 ;
        RECT  6.810 1.080 7.490 1.240 ;
        RECT  6.550 2.900 7.470 3.060 ;
        RECT  6.820 2.050 7.230 2.210 ;
        RECT  6.540 1.530 6.820 2.210 ;
        RECT  6.530 0.940 6.810 1.240 ;
        RECT  6.270 2.790 6.550 3.100 ;
        RECT  5.990 1.080 6.530 1.240 ;
        RECT  6.090 0.560 6.280 0.920 ;
        RECT  2.530 2.900 6.270 3.060 ;
        RECT  5.990 2.050 6.110 2.530 ;
        RECT  5.130 0.760 6.090 0.920 ;
        RECT  5.830 1.080 5.990 2.530 ;
        RECT  5.310 1.080 5.830 1.270 ;
        RECT  4.750 0.440 5.760 0.600 ;
        RECT  5.130 1.660 5.440 1.940 ;
        RECT  5.120 0.760 5.130 1.940 ;
        RECT  4.910 0.760 5.120 2.380 ;
        RECT  4.810 2.120 4.910 2.380 ;
        RECT  4.650 2.120 4.810 2.700 ;
        RECT  4.590 0.440 4.750 1.080 ;
        RECT  2.850 2.540 4.650 2.700 ;
        RECT  4.150 0.920 4.590 1.080 ;
        RECT  3.990 0.920 4.150 2.330 ;
        RECT  2.860 0.440 3.990 0.600 ;
        RECT  3.490 0.920 3.990 1.200 ;
        RECT  3.430 2.120 3.990 2.330 ;
        RECT  3.550 1.360 3.830 1.940 ;
        RECT  3.330 1.360 3.550 1.520 ;
        RECT  3.140 0.770 3.330 1.520 ;
        RECT  3.010 1.680 3.230 2.340 ;
        RECT  1.880 0.770 3.140 0.930 ;
        RECT  2.970 1.680 3.010 1.840 ;
        RECT  2.810 1.090 2.970 1.840 ;
        RECT  2.700 0.440 2.860 0.610 ;
        RECT  2.690 2.000 2.850 2.700 ;
        RECT  2.690 1.090 2.810 1.310 ;
        RECT  0.700 0.450 2.700 0.610 ;
        RECT  2.600 2.000 2.690 2.160 ;
        RECT  2.440 1.740 2.600 2.160 ;
        RECT  2.370 2.320 2.530 3.060 ;
        RECT  1.800 1.740 2.440 1.900 ;
        RECT  2.280 2.320 2.370 2.480 ;
        RECT  2.120 2.060 2.280 2.480 ;
        RECT  1.360 2.060 2.120 2.280 ;
        RECT  1.720 0.770 1.880 1.140 ;
        RECT  1.520 1.600 1.800 1.900 ;
        RECT  1.040 0.770 1.720 0.930 ;
        RECT  1.040 2.930 1.650 3.150 ;
        RECT  1.360 1.090 1.460 1.310 ;
        RECT  1.200 1.090 1.360 2.280 ;
        RECT  0.880 0.770 1.040 3.150 ;
        RECT  0.540 0.450 0.700 1.250 ;
        RECT  0.250 1.090 0.540 1.250 ;
        RECT  0.250 2.120 0.370 2.280 ;
        RECT  0.090 1.090 0.250 2.280 ;
    END
END SDFFHQX1TR

MACRO SDFFXLTR
    CLASS CORE ;
    FOREIGN SDFFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.640 1.520 2.020 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 2.140 1.960 2.360 ;
        RECT  1.840 2.040 1.920 2.360 ;
        RECT  1.680 2.040 1.840 2.720 ;
        RECT  0.250 2.560 1.680 2.720 ;
        RECT  0.250 1.580 0.370 1.860 ;
        RECT  0.090 1.580 0.250 2.720 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.880 1.030 9.120 2.360 ;
        END
        ANTENNADIFFAREA 1.083 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.560 0.690 8.720 2.510 ;
        RECT  8.440 0.690 8.560 1.160 ;
        RECT  8.170 2.350 8.560 2.510 ;
        RECT  8.210 0.690 8.440 0.850 ;
        RECT  7.930 0.550 8.210 0.850 ;
        RECT  7.890 2.350 8.170 2.750 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.320 1.960 ;
        RECT  2.060 1.640 2.080 1.880 ;
        RECT  1.780 1.600 2.060 1.880 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.020 2.040 4.400 2.360 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.670 -0.280 9.200 0.280 ;
        RECT  8.390 -0.280 8.670 0.400 ;
        RECT  7.650 -0.280 8.390 0.280 ;
        RECT  7.370 -0.280 7.650 0.400 ;
        RECT  6.050 -0.280 7.370 0.340 ;
        RECT  5.770 -0.280 6.050 0.890 ;
        RECT  4.650 -0.280 5.770 0.280 ;
        RECT  3.620 -0.280 4.650 0.640 ;
        RECT  1.510 -0.280 3.620 0.340 ;
        RECT  1.230 -0.280 1.510 0.400 ;
        RECT  0.240 -0.280 1.230 0.280 ;
        RECT  0.240 1.030 0.370 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.670 3.320 9.200 3.880 ;
        RECT  8.390 2.670 8.670 3.880 ;
        RECT  7.650 3.320 8.390 3.880 ;
        RECT  7.370 2.800 7.650 3.880 ;
        RECT  6.050 3.320 7.370 3.880 ;
        RECT  5.770 3.200 6.050 3.880 ;
        RECT  5.080 3.320 5.770 3.880 ;
        RECT  4.800 3.200 5.080 3.880 ;
        RECT  4.060 3.260 4.800 3.880 ;
        RECT  3.780 3.200 4.060 3.880 ;
        RECT  1.840 3.260 3.780 3.880 ;
        RECT  1.560 3.200 1.840 3.880 ;
        RECT  0.370 3.320 1.560 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.230 1.470 8.400 1.750 ;
        RECT  8.210 1.030 8.230 2.070 ;
        RECT  8.070 1.030 8.210 2.190 ;
        RECT  7.990 1.030 8.070 1.310 ;
        RECT  7.930 1.910 8.070 2.190 ;
        RECT  7.470 1.910 7.930 2.070 ;
        RECT  7.830 1.470 7.910 1.750 ;
        RECT  7.670 1.260 7.830 1.750 ;
        RECT  7.010 1.260 7.670 1.420 ;
        RECT  7.310 1.580 7.470 2.070 ;
        RECT  7.250 1.580 7.310 1.860 ;
        RECT  6.510 0.500 7.130 0.720 ;
        RECT  6.890 1.260 7.010 2.470 ;
        RECT  6.850 0.880 6.890 2.590 ;
        RECT  6.670 0.880 6.850 1.420 ;
        RECT  6.670 2.310 6.850 2.590 ;
        RECT  6.510 1.870 6.690 2.150 ;
        RECT  6.350 0.500 6.510 3.010 ;
        RECT  5.880 1.170 6.350 1.330 ;
        RECT  4.520 2.850 6.350 3.010 ;
        RECT  5.910 1.620 6.190 2.690 ;
        RECT  5.110 2.410 5.910 2.690 ;
        RECT  5.660 1.050 5.880 1.330 ;
        RECT  5.340 0.440 5.500 2.230 ;
        RECT  5.210 0.440 5.340 0.890 ;
        RECT  4.810 0.440 5.210 0.660 ;
        RECT  5.110 1.070 5.180 1.900 ;
        RECT  4.960 1.070 5.110 2.690 ;
        RECT  4.950 1.700 4.960 2.690 ;
        RECT  3.860 1.700 4.950 1.860 ;
        RECT  3.300 1.380 4.800 1.540 ;
        RECT  4.240 2.520 4.520 3.010 ;
        RECT  4.060 0.860 4.340 1.140 ;
        RECT  3.540 2.850 4.240 3.010 ;
        RECT  3.340 0.860 4.060 1.020 ;
        RECT  3.580 1.700 3.860 2.020 ;
        RECT  3.260 2.850 3.540 3.100 ;
        RECT  3.180 0.620 3.340 1.020 ;
        RECT  3.080 1.380 3.300 2.690 ;
        RECT  2.920 2.850 3.260 3.010 ;
        RECT  2.640 0.620 3.180 0.780 ;
        RECT  3.020 1.380 3.080 1.540 ;
        RECT  2.800 0.940 3.020 1.540 ;
        RECT  2.760 1.840 2.920 3.010 ;
        RECT  2.640 1.840 2.760 2.000 ;
        RECT  2.480 0.620 2.640 2.000 ;
        RECT  2.320 2.410 2.600 3.040 ;
        RECT  2.360 1.160 2.480 1.440 ;
        RECT  2.100 0.560 2.320 1.000 ;
        RECT  0.960 2.880 2.320 3.040 ;
        RECT  0.620 0.560 2.100 0.720 ;
        RECT  1.460 1.060 1.740 1.340 ;
        RECT  0.930 1.150 1.460 1.310 ;
        RECT  0.810 2.180 1.200 2.400 ;
        RECT  0.680 2.880 0.960 3.160 ;
        RECT  0.810 1.030 0.930 1.310 ;
        RECT  0.650 1.030 0.810 2.400 ;
        RECT  0.530 1.910 0.650 2.190 ;
        RECT  0.400 0.440 0.620 0.720 ;
    END
END SDFFXLTR

MACRO SDFFX4TR
    CLASS CORE ;
    FOREIGN SDFFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.630 1.520 1.970 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.960 1.920 2.360 ;
        RECT  1.690 1.960 1.840 2.610 ;
        RECT  1.680 2.040 1.690 2.610 ;
        RECT  0.250 2.450 1.680 2.610 ;
        RECT  0.250 1.680 0.370 1.960 ;
        RECT  0.090 1.680 0.250 2.610 ;
        END
        ANTENNAGATEAREA 0.1512 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.190 1.040 12.320 1.760 ;
        RECT  11.990 0.490 12.190 3.160 ;
        RECT  11.910 0.490 11.990 1.410 ;
        RECT  11.910 2.010 11.990 3.160 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.950 0.490 11.230 2.290 ;
        RECT  10.880 1.040 10.950 1.760 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.370 2.070 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.820 4.760 2.360 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.710 -0.280 12.800 0.280 ;
        RECT  12.490 -0.280 12.710 1.410 ;
        RECT  11.710 -0.280 12.490 0.280 ;
        RECT  11.430 -0.280 11.710 1.410 ;
        RECT  10.690 -0.280 11.430 0.280 ;
        RECT  10.470 -0.280 10.690 1.410 ;
        RECT  9.810 -0.280 10.470 0.280 ;
        RECT  9.590 -0.280 9.810 1.410 ;
        RECT  8.060 -0.280 9.590 0.280 ;
        RECT  7.780 -0.280 8.060 0.600 ;
        RECT  6.340 -0.280 7.780 0.280 ;
        RECT  6.060 -0.280 6.340 0.930 ;
        RECT  4.840 -0.280 6.060 0.280 ;
        RECT  4.560 -0.280 4.840 0.880 ;
        RECT  4.010 -0.280 4.560 0.280 ;
        RECT  3.730 -0.280 4.010 0.950 ;
        RECT  1.770 -0.280 3.730 0.280 ;
        RECT  1.490 -0.280 1.770 0.400 ;
        RECT  0.370 -0.280 1.490 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.670 3.320 12.800 3.880 ;
        RECT  12.390 2.010 12.670 3.880 ;
        RECT  11.710 3.320 12.390 3.880 ;
        RECT  11.430 2.930 11.710 3.880 ;
        RECT  10.750 3.320 11.430 3.880 ;
        RECT  10.470 2.930 10.750 3.880 ;
        RECT  9.810 3.320 10.470 3.880 ;
        RECT  9.530 2.330 9.810 3.880 ;
        RECT  8.020 3.320 9.530 3.880 ;
        RECT  7.740 2.890 8.020 3.880 ;
        RECT  6.300 3.320 7.740 3.880 ;
        RECT  6.020 3.240 6.300 3.880 ;
        RECT  4.790 3.260 6.020 3.880 ;
        RECT  4.090 3.320 4.790 3.880 ;
        RECT  3.810 3.260 4.090 3.880 ;
        RECT  1.850 3.320 3.810 3.880 ;
        RECT  1.570 3.200 1.850 3.880 ;
        RECT  0.370 3.320 1.570 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.710 1.570 11.830 1.850 ;
        RECT  11.550 1.570 11.710 2.610 ;
        RECT  10.310 2.450 11.550 2.610 ;
        RECT  10.290 0.590 10.310 2.610 ;
        RECT  10.150 0.590 10.290 3.160 ;
        RECT  10.010 0.590 10.150 1.410 ;
        RECT  10.010 2.010 10.150 3.160 ;
        RECT  9.370 2.010 10.010 2.170 ;
        RECT  9.710 1.570 9.990 1.850 ;
        RECT  9.430 1.580 9.710 1.740 ;
        RECT  9.270 0.760 9.430 1.740 ;
        RECT  9.210 2.010 9.370 3.130 ;
        RECT  6.940 0.760 9.270 0.980 ;
        RECT  8.940 1.580 9.270 1.740 ;
        RECT  9.090 2.850 9.210 3.130 ;
        RECT  8.830 1.140 9.110 1.420 ;
        RECT  8.820 1.580 8.940 2.540 ;
        RECT  8.500 1.140 8.830 1.300 ;
        RECT  8.780 1.580 8.820 3.160 ;
        RECT  8.540 2.380 8.780 3.160 ;
        RECT  8.500 1.860 8.620 2.220 ;
        RECT  7.220 2.380 8.540 2.540 ;
        RECT  8.340 1.140 8.500 2.220 ;
        RECT  6.180 1.140 8.340 1.300 ;
        RECT  7.060 2.060 8.340 2.220 ;
        RECT  7.540 1.520 8.180 1.800 ;
        RECT  6.620 1.520 7.540 1.680 ;
        RECT  6.940 2.380 7.220 3.160 ;
        RECT  6.780 1.840 7.060 2.220 ;
        RECT  6.540 2.060 6.780 2.220 ;
        RECT  6.340 1.520 6.620 1.900 ;
        RECT  6.380 2.060 6.540 3.070 ;
        RECT  3.570 2.850 6.380 3.070 ;
        RECT  6.220 1.740 6.340 1.900 ;
        RECT  6.060 1.740 6.220 2.690 ;
        RECT  6.020 1.140 6.180 1.580 ;
        RECT  5.370 2.470 6.060 2.690 ;
        RECT  5.850 1.300 6.020 1.580 ;
        RECT  5.690 2.010 5.900 2.290 ;
        RECT  5.690 0.860 5.860 1.140 ;
        RECT  5.530 0.440 5.690 2.290 ;
        RECT  5.330 0.440 5.530 0.720 ;
        RECT  5.190 1.050 5.370 2.690 ;
        RECT  5.090 1.050 5.190 1.330 ;
        RECT  3.970 2.530 5.190 2.690 ;
        RECT  4.650 1.380 4.930 1.660 ;
        RECT  3.330 1.500 4.650 1.660 ;
        RECT  4.210 1.060 4.490 1.340 ;
        RECT  3.530 1.180 4.210 1.340 ;
        RECT  3.810 1.820 3.970 2.690 ;
        RECT  3.690 1.820 3.810 2.100 ;
        RECT  3.290 2.850 3.570 3.130 ;
        RECT  3.370 0.550 3.530 1.340 ;
        RECT  2.750 0.550 3.370 0.710 ;
        RECT  3.210 1.500 3.330 2.570 ;
        RECT  2.890 2.850 3.290 3.010 ;
        RECT  3.130 0.990 3.210 2.570 ;
        RECT  3.050 0.870 3.130 2.570 ;
        RECT  2.910 0.870 3.050 1.150 ;
        RECT  2.750 1.320 2.890 3.010 ;
        RECT  2.730 0.550 2.750 3.010 ;
        RECT  2.590 0.550 2.730 1.480 ;
        RECT  2.470 1.200 2.590 1.480 ;
        RECT  2.290 2.590 2.570 2.930 ;
        RECT  2.210 0.560 2.430 1.010 ;
        RECT  0.970 2.770 2.290 2.930 ;
        RECT  0.830 0.560 2.210 0.720 ;
        RECT  1.610 1.200 1.890 1.480 ;
        RECT  0.810 1.200 1.610 1.360 ;
        RECT  0.810 2.130 1.210 2.290 ;
        RECT  0.690 2.770 0.970 3.050 ;
        RECT  0.550 0.440 0.830 0.720 ;
        RECT  0.690 1.030 0.810 1.360 ;
        RECT  0.690 2.010 0.810 2.290 ;
        RECT  0.530 1.030 0.690 2.290 ;
    END
END SDFFX4TR

MACRO SDFFX2TR
    CLASS CORE ;
    FOREIGN SDFFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.600 1.520 2.080 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 2.120 2.000 2.360 ;
        RECT  1.840 2.040 1.920 2.360 ;
        RECT  1.680 2.040 1.840 2.720 ;
        RECT  0.470 2.560 1.680 2.720 ;
        RECT  0.470 1.470 0.550 1.750 ;
        RECT  0.310 1.470 0.470 2.720 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.680 0.440 9.920 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.600 2.040 8.720 2.360 ;
        RECT  8.480 0.450 8.600 2.360 ;
        RECT  8.440 0.450 8.480 2.210 ;
        RECT  8.340 0.450 8.440 0.670 ;
        RECT  8.320 1.930 8.440 2.210 ;
        END
        ANTENNADIFFAREA 2.536 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.920 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.440 2.040 4.720 2.360 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.380 -0.280 10.000 0.280 ;
        RECT  9.100 -0.280 9.380 0.410 ;
        RECT  8.100 -0.280 9.100 0.280 ;
        RECT  7.740 -0.280 8.100 0.300 ;
        RECT  6.280 -0.280 7.740 0.280 ;
        RECT  6.000 -0.280 6.280 0.340 ;
        RECT  4.870 -0.280 6.000 0.280 ;
        RECT  3.880 -0.280 4.870 0.340 ;
        RECT  1.620 -0.280 3.880 0.280 ;
        RECT  1.290 -0.280 1.620 0.340 ;
        RECT  0.240 -0.280 1.290 0.280 ;
        RECT  0.240 1.030 0.310 1.310 ;
        RECT  0.080 -0.280 0.240 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.360 3.320 10.000 3.880 ;
        RECT  9.200 2.570 9.360 3.880 ;
        RECT  8.030 3.320 9.200 3.880 ;
        RECT  7.810 2.930 8.030 3.880 ;
        RECT  6.120 3.320 7.810 3.880 ;
        RECT  5.840 3.260 6.120 3.880 ;
        RECT  4.980 3.320 5.840 3.880 ;
        RECT  4.700 3.260 4.980 3.880 ;
        RECT  4.000 3.320 4.700 3.880 ;
        RECT  3.720 3.260 4.000 3.880 ;
        RECT  1.880 3.320 3.720 3.880 ;
        RECT  1.600 3.260 1.880 3.880 ;
        RECT  0.410 3.320 1.600 3.880 ;
        RECT  0.130 3.260 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.040 1.330 9.520 1.610 ;
        RECT  8.920 1.330 9.040 2.850 ;
        RECT  8.880 1.000 8.920 2.850 ;
        RECT  8.760 1.000 8.880 1.530 ;
        RECT  8.720 2.570 8.880 2.850 ;
        RECT  7.600 2.570 8.720 2.730 ;
        RECT  8.130 1.330 8.280 1.640 ;
        RECT  7.970 0.460 8.130 2.330 ;
        RECT  6.840 0.460 7.970 0.620 ;
        RECT  7.000 2.170 7.970 2.330 ;
        RECT  7.650 0.810 7.810 1.930 ;
        RECT  5.830 0.810 7.650 0.970 ;
        RECT  6.400 1.770 7.650 1.930 ;
        RECT  7.440 2.570 7.600 2.970 ;
        RECT  7.210 1.130 7.490 1.530 ;
        RECT  5.700 1.130 7.210 1.290 ;
        RECT  6.650 2.170 7.000 3.160 ;
        RECT  6.240 1.770 6.400 3.100 ;
        RECT  6.080 1.450 6.360 1.610 ;
        RECT  4.400 2.940 6.240 3.100 ;
        RECT  5.920 1.450 6.080 2.780 ;
        RECT  5.320 2.620 5.920 2.780 ;
        RECT  5.660 0.480 5.720 0.640 ;
        RECT  5.660 1.130 5.700 2.190 ;
        RECT  5.500 0.480 5.660 2.190 ;
        RECT  5.440 0.480 5.500 0.670 ;
        RECT  3.100 0.510 5.440 0.670 ;
        RECT  5.160 0.940 5.320 2.780 ;
        RECT  3.740 1.670 5.160 1.830 ;
        RECT  5.090 2.620 5.160 2.780 ;
        RECT  3.180 1.350 5.000 1.510 ;
        RECT  2.760 0.830 4.520 0.990 ;
        RECT  4.240 2.760 4.400 3.100 ;
        RECT  3.420 2.830 4.240 3.100 ;
        RECT  3.580 1.670 3.740 1.950 ;
        RECT  3.260 2.830 3.420 3.110 ;
        RECT  2.860 2.830 3.260 2.990 ;
        RECT  3.080 1.350 3.180 2.670 ;
        RECT  3.020 1.150 3.080 2.670 ;
        RECT  2.920 1.150 3.020 1.510 ;
        RECT  2.760 1.670 2.860 2.990 ;
        RECT  2.700 0.830 2.760 2.990 ;
        RECT  2.600 0.830 2.700 1.830 ;
        RECT  2.480 1.380 2.600 1.540 ;
        RECT  2.380 2.430 2.540 3.040 ;
        RECT  2.280 0.560 2.440 1.080 ;
        RECT  0.940 2.880 2.380 3.040 ;
        RECT  0.560 0.560 2.280 0.720 ;
        RECT  0.870 1.150 1.860 1.310 ;
        RECT  0.870 2.240 1.240 2.400 ;
        RECT  0.780 2.880 0.940 3.160 ;
        RECT  0.710 1.030 0.870 2.400 ;
        RECT  0.630 1.910 0.710 2.190 ;
        RECT  0.400 0.440 0.560 0.720 ;
    END
END SDFFX2TR

MACRO SDFFX1TR
    CLASS CORE ;
    FOREIGN SDFFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.580 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 2.140 1.980 2.360 ;
        RECT  1.840 2.040 1.920 2.360 ;
        RECT  1.680 2.040 1.840 2.700 ;
        RECT  0.430 2.540 1.680 2.700 ;
        RECT  0.270 1.580 0.430 2.700 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.440 1.240 9.520 2.360 ;
        RECT  9.280 1.030 9.440 2.550 ;
        END
        ANTENNADIFFAREA 1.98 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.040 0.840 9.120 2.630 ;
        RECT  8.960 0.690 9.040 2.630 ;
        RECT  8.880 0.690 8.960 1.160 ;
        RECT  8.520 2.470 8.960 2.630 ;
        RECT  8.500 0.690 8.880 0.850 ;
        RECT  8.360 2.470 8.520 2.850 ;
        RECT  8.340 0.490 8.500 0.850 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.320 1.980 ;
        RECT  1.940 1.640 2.080 1.870 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.250 2.080 4.700 2.240 ;
        RECT  4.090 2.080 4.250 2.600 ;
        RECT  3.920 2.440 4.090 2.600 ;
        RECT  3.680 2.440 3.920 2.760 ;
        END
        ANTENNAGATEAREA 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.060 -0.280 9.600 0.280 ;
        RECT  8.780 -0.280 9.060 0.340 ;
        RECT  8.040 -0.280 8.780 0.280 ;
        RECT  7.760 -0.280 8.040 0.900 ;
        RECT  6.280 -0.280 7.760 0.280 ;
        RECT  6.120 -0.280 6.280 0.820 ;
        RECT  4.910 -0.280 6.120 0.280 ;
        RECT  3.970 -0.280 4.910 0.660 ;
        RECT  1.780 -0.280 3.970 0.280 ;
        RECT  1.500 -0.280 1.780 0.340 ;
        RECT  0.310 -0.280 1.500 0.280 ;
        RECT  0.150 -0.280 0.310 1.310 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.090 3.320 9.600 3.880 ;
        RECT  8.790 2.860 9.090 3.880 ;
        RECT  8.040 3.320 8.790 3.880 ;
        RECT  7.700 2.800 8.040 3.880 ;
        RECT  6.220 3.320 7.700 3.880 ;
        RECT  5.940 3.260 6.220 3.880 ;
        RECT  5.160 3.320 5.940 3.880 ;
        RECT  4.880 3.260 5.160 3.880 ;
        RECT  4.180 3.320 4.880 3.880 ;
        RECT  3.900 3.260 4.180 3.880 ;
        RECT  1.860 3.320 3.900 3.880 ;
        RECT  1.580 3.260 1.860 3.880 ;
        RECT  0.370 3.320 1.580 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.540 1.490 8.800 1.650 ;
        RECT  8.520 1.030 8.540 2.070 ;
        RECT  8.380 1.030 8.520 2.310 ;
        RECT  8.360 1.910 8.380 2.310 ;
        RECT  7.640 1.910 8.360 2.070 ;
        RECT  8.060 1.380 8.220 1.750 ;
        RECT  7.180 1.380 8.060 1.540 ;
        RECT  7.480 1.700 7.640 2.070 ;
        RECT  6.680 0.710 7.520 0.870 ;
        RECT  7.020 1.030 7.180 2.240 ;
        RECT  6.960 1.030 7.020 1.310 ;
        RECT  7.000 2.080 7.020 2.240 ;
        RECT  6.840 2.080 7.000 2.830 ;
        RECT  6.680 1.760 6.860 1.920 ;
        RECT  6.520 0.710 6.680 3.100 ;
        RECT  6.110 0.980 6.520 1.140 ;
        RECT  4.580 2.940 6.520 3.100 ;
        RECT  6.200 1.420 6.360 2.700 ;
        RECT  5.350 2.540 6.200 2.700 ;
        RECT  5.950 0.980 6.110 1.260 ;
        RECT  5.630 0.440 5.790 2.220 ;
        RECT  5.560 0.440 5.630 0.930 ;
        RECT  5.510 2.060 5.630 2.220 ;
        RECT  5.100 0.440 5.560 0.600 ;
        RECT  5.350 1.110 5.470 1.900 ;
        RECT  5.310 1.110 5.350 2.700 ;
        RECT  5.190 1.740 5.310 2.700 ;
        RECT  3.920 1.740 5.190 1.900 ;
        RECT  3.250 1.420 5.150 1.580 ;
        RECT  4.420 2.660 4.580 3.100 ;
        RECT  4.410 0.970 4.570 1.250 ;
        RECT  2.930 2.940 4.420 3.100 ;
        RECT  3.570 0.970 4.410 1.130 ;
        RECT  3.760 1.740 3.920 2.020 ;
        RECT  3.410 0.710 3.570 1.130 ;
        RECT  2.930 0.710 3.410 0.870 ;
        RECT  3.090 1.030 3.250 2.690 ;
        RECT  2.770 0.710 2.930 3.100 ;
        RECT  2.500 1.390 2.770 1.550 ;
        RECT  2.400 2.410 2.560 3.020 ;
        RECT  2.320 0.560 2.480 1.230 ;
        RECT  0.920 2.860 2.400 3.020 ;
        RECT  0.840 0.560 2.320 0.720 ;
        RECT  1.680 1.200 1.840 1.480 ;
        RECT  0.870 1.200 1.680 1.360 ;
        RECT  0.870 2.220 1.220 2.380 ;
        RECT  0.760 2.860 0.920 3.140 ;
        RECT  0.710 1.030 0.870 2.380 ;
        RECT  0.680 0.440 0.840 0.720 ;
        RECT  0.590 1.910 0.710 2.190 ;
    END
END SDFFX1TR

MACRO RF1R1WX1TR
    CLASS CORE ;
    FOREIGN RF1R1WX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.280 2.350 1.560 2.760 ;
        RECT  1.250 2.480 1.280 2.760 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.360 0.350 2.760 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.640 3.520 2.760 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 0.870 3.200 1.160 ;
        RECT  2.880 0.840 3.160 1.160 ;
        END
        ANTENNAGATEAREA 0.0504 ;
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.450 3.520 1.480 ;
        RECT  3.110 2.920 3.470 3.150 ;
        RECT  3.230 0.450 3.360 0.670 ;
        RECT  3.110 1.320 3.360 1.480 ;
        RECT  2.950 1.320 3.110 3.150 ;
        RECT  2.440 2.440 2.950 2.760 ;
        END
        ANTENNAGATEAREA 1.801 ;
    END RB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 -0.280 3.600 0.280 ;
        RECT  2.300 -0.280 2.580 0.800 ;
        RECT  0.370 -0.280 2.300 0.280 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 3.320 3.600 3.880 ;
        RECT  2.180 3.200 2.580 3.880 ;
        RECT  1.900 2.860 2.180 3.880 ;
        RECT  0.370 3.320 1.900 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.700 1.430 2.790 1.710 ;
        RECT  2.620 1.240 2.700 2.280 ;
        RECT  2.540 1.030 2.620 2.280 ;
        RECT  2.340 1.030 2.540 1.400 ;
        RECT  2.410 2.000 2.540 2.280 ;
        RECT  2.250 1.560 2.380 1.840 ;
        RECT  1.930 1.240 2.340 1.400 ;
        RECT  2.090 1.560 2.250 1.960 ;
        RECT  1.210 1.800 2.090 1.960 ;
        RECT  1.650 1.240 1.930 1.640 ;
        RECT  0.930 0.500 1.610 0.800 ;
        RECT  0.710 2.920 1.330 3.140 ;
        RECT  1.090 1.030 1.210 1.960 ;
        RECT  0.930 1.030 1.090 2.570 ;
        RECT  0.710 0.640 0.930 0.800 ;
        RECT  0.870 1.880 0.930 2.570 ;
        RECT  0.550 0.640 0.710 3.140 ;
    END
END RF1R1WX1TR

MACRO RF2R1WX1TR
    CLASS CORE ;
    FOREIGN RF2R1WX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.260 2.440 2.320 2.760 ;
        RECT  2.020 2.440 2.260 2.860 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.480 1.240 6.720 2.760 ;
        RECT  6.360 1.240 6.480 1.620 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  5.560 0.990 5.860 1.270 ;
        RECT  5.440 2.880 5.820 3.160 ;
        RECT  5.440 0.840 5.560 1.270 ;
        RECT  5.280 0.840 5.440 3.160 ;
        END
        ANTENNAGATEAREA 2.784 ;
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.720 1.760 4.800 2.040 ;
        RECT  4.480 1.640 4.720 2.040 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.920 2.880 4.060 3.160 ;
        RECT  3.920 1.000 4.000 1.280 ;
        RECT  3.760 1.000 3.920 3.160 ;
        RECT  3.640 2.840 3.760 3.160 ;
        END
        ANTENNAGATEAREA 2.866 ;
    END R1B
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.320 -0.280 6.800 0.280 ;
        RECT  6.040 -0.280 6.320 0.580 ;
        RECT  5.020 -0.280 6.040 0.280 ;
        RECT  4.740 -0.280 5.020 0.400 ;
        RECT  3.260 -0.280 4.740 0.280 ;
        RECT  2.980 -0.280 3.260 0.800 ;
        RECT  1.880 -0.280 2.980 0.280 ;
        RECT  1.600 -0.280 1.880 0.730 ;
        RECT  0.380 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.340 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.320 3.320 6.800 3.880 ;
        RECT  6.050 2.540 6.320 3.880 ;
        RECT  5.020 3.320 6.050 3.880 ;
        RECT  4.250 2.930 5.020 3.880 ;
        RECT  3.260 3.320 4.250 3.880 ;
        RECT  2.980 2.290 3.260 3.880 ;
        RECT  1.860 3.320 2.980 3.880 ;
        RECT  1.580 2.500 1.860 3.880 ;
        RECT  0.380 3.320 1.580 3.880 ;
        RECT  0.100 3.200 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.180 0.860 6.380 1.080 ;
        RECT  6.180 2.060 6.320 2.340 ;
        RECT  6.020 0.860 6.180 2.340 ;
        RECT  5.750 1.660 6.020 1.940 ;
        RECT  5.060 1.320 5.120 1.600 ;
        RECT  4.900 0.680 5.060 1.600 ;
        RECT  3.580 0.680 4.900 0.840 ;
        RECT  4.320 1.030 4.650 1.310 ;
        RECT  4.300 2.360 4.530 2.640 ;
        RECT  4.300 1.030 4.320 1.600 ;
        RECT  4.160 1.030 4.300 2.640 ;
        RECT  4.080 1.440 4.160 2.640 ;
        RECT  3.460 0.680 3.580 1.370 ;
        RECT  3.420 0.680 3.460 1.890 ;
        RECT  3.340 1.210 3.420 1.890 ;
        RECT  3.180 1.210 3.340 2.130 ;
        RECT  2.780 1.210 3.180 1.370 ;
        RECT  2.780 1.970 3.180 2.130 ;
        RECT  2.060 1.530 2.980 1.810 ;
        RECT  2.500 1.030 2.780 1.370 ;
        RECT  2.620 1.970 2.780 3.080 ;
        RECT  2.500 2.800 2.620 3.080 ;
        RECT  1.740 1.210 2.500 1.370 ;
        RECT  2.320 0.520 2.440 0.800 ;
        RECT  2.220 1.970 2.440 2.250 ;
        RECT  2.160 0.520 2.320 1.050 ;
        RECT  1.420 2.090 2.220 2.250 ;
        RECT  1.420 0.890 2.160 1.050 ;
        RECT  1.900 1.530 2.060 1.900 ;
        RECT  1.100 1.740 1.900 1.900 ;
        RECT  1.460 1.210 1.740 1.580 ;
        RECT  1.260 0.530 1.420 1.050 ;
        RECT  1.260 2.090 1.420 2.980 ;
        RECT  0.660 0.530 1.260 0.810 ;
        RECT  0.900 2.820 1.260 2.980 ;
        RECT  0.820 0.970 1.100 2.660 ;
        RECT  0.660 2.820 0.900 3.100 ;
        RECT  0.620 0.530 0.660 3.100 ;
        RECT  0.500 0.530 0.620 2.980 ;
    END
END RF2R1WX1TR

MACRO RFRDX4TR
    CLASS CORE ;
    FOREIGN RFRDX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.520 2.310 1.400 ;
        RECT  2.050 1.910 2.170 2.190 ;
        RECT  2.030 0.520 2.150 0.800 ;
        RECT  2.050 1.240 2.150 1.400 ;
        RECT  1.890 1.240 2.050 2.190 ;
        RECT  1.520 1.240 1.890 1.400 ;
        RECT  1.290 0.840 1.520 1.400 ;
        RECT  1.280 0.840 1.290 1.640 ;
        RECT  0.970 1.240 1.280 1.640 ;
        RECT  0.930 1.360 0.970 1.640 ;
        END
        ANTENNAGATEAREA 0.528 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.580 1.730 1.860 ;
        RECT  1.450 1.580 1.610 2.000 ;
        RECT  1.120 1.840 1.450 2.000 ;
        RECT  0.810 1.840 1.120 2.560 ;
        RECT  0.770 0.440 0.810 1.200 ;
        RECT  0.770 1.840 0.810 3.160 ;
        RECT  0.530 0.440 0.770 3.160 ;
        END
        ANTENNADIFFAREA 0.2584 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.280 2.400 0.280 ;
        RECT  1.090 -0.280 1.370 0.590 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 3.320 2.400 3.880 ;
        RECT  1.090 2.800 1.370 3.880 ;
        RECT  0.350 3.320 1.090 3.880 ;
        RECT  0.090 1.910 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END RFRDX4TR

MACRO RFRDX2TR
    CLASS CORE ;
    FOREIGN RFRDX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.520 1.840 1.400 ;
        RECT  1.560 0.520 1.680 0.800 ;
        RECT  1.520 1.240 1.680 1.400 ;
        RECT  1.520 1.910 1.640 2.190 ;
        RECT  1.360 1.240 1.520 2.190 ;
        RECT  0.760 1.240 1.360 1.400 ;
        RECT  0.480 1.240 0.760 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.580 1.200 1.860 ;
        RECT  0.920 1.580 1.080 2.070 ;
        RECT  0.380 1.910 0.920 2.070 ;
        RECT  0.240 1.910 0.380 3.160 ;
        RECT  0.240 0.500 0.320 1.310 ;
        RECT  0.080 0.500 0.240 3.160 ;
        END
        ANTENNADIFFAREA 0.2584 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.280 2.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.800 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 3.320 2.000 3.880 ;
        RECT  0.620 2.800 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
END RFRDX2TR

MACRO RFRDX1TR
    CLASS CORE ;
    FOREIGN RFRDX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 0.520 1.820 1.000 ;
        RECT  1.520 1.910 1.640 2.190 ;
        RECT  1.520 0.840 1.600 1.000 ;
        RECT  1.360 0.840 1.520 2.190 ;
        RECT  0.740 0.840 1.360 1.000 ;
        RECT  0.480 0.840 0.740 1.730 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.520 1.200 2.220 ;
        RECT  0.400 2.060 0.920 2.220 ;
        RECT  0.320 2.060 0.400 2.550 ;
        RECT  0.240 0.930 0.320 1.260 ;
        RECT  0.240 1.640 0.320 2.760 ;
        RECT  0.080 0.930 0.240 2.760 ;
        END
        ANTENNADIFFAREA 0.2584 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 3.320 2.000 3.880 ;
        RECT  0.640 2.800 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
END RFRDX1TR

MACRO BENCX4TR
    CLASS CORE ;
    FOREIGN BENCX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 32.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  22.050 0.900 22.370 2.080 ;
        RECT  21.290 0.900 22.050 1.140 ;
        RECT  18.930 1.860 22.050 2.080 ;
        RECT  21.010 0.810 21.290 1.140 ;
        RECT  20.250 0.810 21.010 1.050 ;
        RECT  18.930 0.770 20.250 1.050 ;
        END
        ANTENNADIFFAREA 15.624 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  31.870 1.040 31.920 1.760 ;
        RECT  31.830 0.950 31.870 2.070 ;
        RECT  31.570 0.950 31.830 3.160 ;
        RECT  31.550 1.070 31.570 3.160 ;
        RECT  30.890 1.070 31.550 1.310 ;
        RECT  30.870 1.910 31.550 2.150 ;
        RECT  30.610 0.440 30.890 1.310 ;
        RECT  30.590 1.910 30.870 3.160 ;
        RECT  29.930 1.070 30.610 1.310 ;
        RECT  29.910 1.910 30.590 2.150 ;
        RECT  29.650 0.440 29.930 1.310 ;
        RECT  29.630 1.910 29.910 3.160 ;
        RECT  28.970 1.070 29.650 1.310 ;
        RECT  28.950 1.910 29.630 2.150 ;
        RECT  28.690 0.440 28.970 1.310 ;
        RECT  28.670 1.910 28.950 3.160 ;
        END
        ANTENNADIFFAREA 15.871 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  23.010 2.880 23.290 3.160 ;
        RECT  15.270 2.880 23.010 3.040 ;
        RECT  15.110 2.880 15.270 3.150 ;
        RECT  12.550 2.990 15.110 3.150 ;
        RECT  12.390 2.840 12.550 3.150 ;
        RECT  9.160 2.840 12.390 3.000 ;
        RECT  8.840 2.840 9.160 3.160 ;
        RECT  8.810 2.840 8.840 3.120 ;
        END
        ANTENNAGATEAREA 0.372 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.740 1.640 12.860 1.920 ;
        RECT  12.580 1.640 12.740 2.680 ;
        RECT  8.510 2.520 12.580 2.680 ;
        RECT  8.350 1.990 8.510 2.680 ;
        RECT  7.510 1.990 8.350 2.150 ;
        RECT  7.350 1.550 7.510 2.150 ;
        RECT  7.230 1.550 7.350 1.960 ;
        RECT  6.320 1.800 7.230 1.960 ;
        RECT  6.030 1.580 6.320 1.960 ;
        END
        ANTENNAGATEAREA 1.008 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.510 1.640 10.670 1.920 ;
        RECT  10.350 0.640 10.510 1.920 ;
        RECT  9.650 0.640 10.350 0.800 ;
        RECT  9.490 0.640 9.650 1.390 ;
        RECT  6.760 1.230 9.490 1.390 ;
        RECT  6.480 1.230 6.760 1.640 ;
        END
        ANTENNAGATEAREA 1.008 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.440 3.730 1.310 ;
        RECT  3.450 1.910 3.730 3.160 ;
        RECT  2.770 1.070 3.450 1.310 ;
        RECT  2.770 1.910 3.450 2.150 ;
        RECT  2.490 0.440 2.770 1.310 ;
        RECT  2.490 1.910 2.770 3.160 ;
        RECT  1.810 1.070 2.490 1.310 ;
        RECT  1.810 1.910 2.490 2.150 ;
        RECT  1.530 0.440 1.810 1.310 ;
        RECT  1.530 1.910 1.810 3.160 ;
        RECT  0.850 1.070 1.530 1.310 ;
        RECT  0.850 1.910 1.530 2.150 ;
        RECT  0.570 0.440 0.850 3.160 ;
        RECT  0.530 1.040 0.570 2.070 ;
        RECT  0.480 1.040 0.530 1.760 ;
        END
        ANTENNADIFFAREA 15.984 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  31.370 -0.280 32.400 0.280 ;
        RECT  31.090 -0.280 31.370 0.670 ;
        RECT  30.410 -0.280 31.090 0.280 ;
        RECT  30.130 -0.280 30.410 0.670 ;
        RECT  29.450 -0.280 30.130 0.280 ;
        RECT  29.170 -0.280 29.450 0.670 ;
        RECT  28.450 -0.280 29.170 0.280 ;
        RECT  28.170 -0.280 28.450 0.350 ;
        RECT  24.330 -0.280 28.170 0.340 ;
        RECT  22.850 -0.280 24.330 0.280 ;
        RECT  22.570 -0.280 22.850 0.290 ;
        RECT  21.810 -0.280 22.570 0.280 ;
        RECT  21.530 -0.280 21.810 0.290 ;
        RECT  20.770 -0.280 21.530 0.280 ;
        RECT  20.490 -0.280 20.770 0.290 ;
        RECT  19.730 -0.280 20.490 0.280 ;
        RECT  19.450 -0.280 19.730 0.290 ;
        RECT  18.690 -0.280 19.450 0.280 ;
        RECT  18.410 -0.280 18.690 0.290 ;
        RECT  17.790 -0.280 18.410 0.280 ;
        RECT  17.510 -0.280 17.790 0.290 ;
        RECT  16.750 -0.280 17.510 0.280 ;
        RECT  16.470 -0.280 16.750 0.290 ;
        RECT  12.890 -0.280 16.470 0.280 ;
        RECT  12.610 -0.280 12.890 0.400 ;
        RECT  11.430 -0.280 12.610 0.280 ;
        RECT  11.150 -0.280 11.430 1.240 ;
        RECT  10.430 -0.280 11.150 0.280 ;
        RECT  10.150 -0.280 10.430 0.400 ;
        RECT  8.090 -0.280 10.150 0.280 ;
        RECT  7.810 -0.280 8.090 0.310 ;
        RECT  7.050 -0.280 7.810 0.280 ;
        RECT  6.770 -0.280 7.050 0.310 ;
        RECT  6.010 -0.280 6.770 0.280 ;
        RECT  5.730 -0.280 6.010 0.370 ;
        RECT  5.130 -0.280 5.730 0.340 ;
        RECT  4.850 -0.280 5.130 0.960 ;
        RECT  4.250 -0.280 4.850 0.340 ;
        RECT  3.970 -0.280 4.250 0.370 ;
        RECT  3.250 -0.280 3.970 0.280 ;
        RECT  2.970 -0.280 3.250 0.670 ;
        RECT  2.290 -0.280 2.970 0.280 ;
        RECT  2.010 -0.280 2.290 0.670 ;
        RECT  1.330 -0.280 2.010 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.320 -0.280 0.370 0.880 ;
        RECT  0.090 -0.280 0.320 1.140 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  32.310 3.320 32.400 3.880 ;
        RECT  32.030 1.920 32.310 3.880 ;
        RECT  31.350 3.320 32.030 3.880 ;
        RECT  31.070 2.450 31.350 3.880 ;
        RECT  30.390 3.320 31.070 3.880 ;
        RECT  30.110 2.440 30.390 3.880 ;
        RECT  29.430 3.320 30.110 3.880 ;
        RECT  29.150 2.390 29.430 3.880 ;
        RECT  28.470 3.320 29.150 3.880 ;
        RECT  28.190 1.910 28.470 3.880 ;
        RECT  27.510 3.260 28.190 3.880 ;
        RECT  27.230 2.120 27.510 3.880 ;
        RECT  26.550 3.260 27.230 3.880 ;
        RECT  26.270 2.140 26.550 3.880 ;
        RECT  25.890 3.260 26.270 3.880 ;
        RECT  25.610 2.140 25.890 3.880 ;
        RECT  24.210 3.320 25.610 3.880 ;
        RECT  23.930 2.780 24.210 3.880 ;
        RECT  22.850 3.320 23.930 3.880 ;
        RECT  22.570 3.200 22.850 3.880 ;
        RECT  21.810 3.320 22.570 3.880 ;
        RECT  21.530 3.200 21.810 3.880 ;
        RECT  20.770 3.320 21.530 3.880 ;
        RECT  20.490 3.200 20.770 3.880 ;
        RECT  19.730 3.320 20.490 3.880 ;
        RECT  19.450 3.200 19.730 3.880 ;
        RECT  18.690 3.320 19.450 3.880 ;
        RECT  18.410 3.200 18.690 3.880 ;
        RECT  17.710 3.260 18.410 3.880 ;
        RECT  17.430 3.200 17.710 3.880 ;
        RECT  16.630 3.320 17.430 3.880 ;
        RECT  16.350 3.200 16.630 3.880 ;
        RECT  15.710 3.260 16.350 3.880 ;
        RECT  15.430 3.200 15.710 3.880 ;
        RECT  12.230 3.320 15.430 3.880 ;
        RECT  11.950 3.200 12.230 3.880 ;
        RECT  11.190 3.320 11.950 3.880 ;
        RECT  10.910 3.200 11.190 3.880 ;
        RECT  10.150 3.320 10.910 3.880 ;
        RECT  9.870 3.200 10.150 3.880 ;
        RECT  8.650 3.320 9.870 3.880 ;
        RECT  8.370 2.840 8.650 3.880 ;
        RECT  7.710 3.320 8.370 3.880 ;
        RECT  7.430 2.630 7.710 3.880 ;
        RECT  6.070 3.320 7.430 3.880 ;
        RECT  5.790 3.200 6.070 3.880 ;
        RECT  5.130 3.260 5.790 3.880 ;
        RECT  4.850 2.400 5.130 3.880 ;
        RECT  4.250 3.260 4.850 3.880 ;
        RECT  3.970 3.180 4.250 3.880 ;
        RECT  3.250 3.320 3.970 3.880 ;
        RECT  2.970 2.440 3.250 3.880 ;
        RECT  2.290 3.320 2.970 3.880 ;
        RECT  2.010 2.480 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.490 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 1.910 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  28.470 1.470 31.390 1.750 ;
        RECT  28.050 1.470 28.470 1.630 ;
        RECT  28.030 0.900 28.050 1.630 ;
        RECT  27.890 0.900 28.030 2.680 ;
        RECT  27.770 0.900 27.890 1.180 ;
        RECT  27.870 1.530 27.890 2.680 ;
        RECT  27.710 1.800 27.870 2.680 ;
        RECT  27.130 0.900 27.770 1.060 ;
        RECT  26.530 1.360 27.710 1.640 ;
        RECT  27.030 1.800 27.710 1.960 ;
        RECT  26.850 0.840 27.130 1.120 ;
        RECT  26.870 1.800 27.030 2.680 ;
        RECT  26.750 2.140 26.870 2.680 ;
        RECT  26.370 0.500 26.530 1.980 ;
        RECT  23.450 0.500 26.370 0.780 ;
        RECT  25.210 1.820 26.370 1.980 ;
        RECT  22.970 0.940 26.210 1.220 ;
        RECT  25.730 1.380 26.010 1.660 ;
        RECT  24.890 1.380 25.730 1.540 ;
        RECT  25.090 1.820 25.210 2.310 ;
        RECT  25.050 1.820 25.090 3.060 ;
        RECT  24.810 2.150 25.050 3.060 ;
        RECT  24.650 1.380 24.890 1.990 ;
        RECT  23.730 2.460 24.810 2.620 ;
        RECT  24.490 1.380 24.650 2.300 ;
        RECT  22.690 1.380 24.490 1.540 ;
        RECT  23.010 2.140 24.490 2.300 ;
        RECT  24.050 1.700 24.330 1.980 ;
        RECT  22.690 1.820 24.050 1.980 ;
        RECT  23.450 2.460 23.730 2.740 ;
        RECT  22.850 2.140 23.010 2.720 ;
        RECT  15.110 2.560 22.850 2.720 ;
        RECT  22.530 0.450 22.690 1.540 ;
        RECT  22.530 1.820 22.690 2.400 ;
        RECT  15.750 0.450 22.530 0.610 ;
        RECT  16.230 2.240 22.530 2.400 ;
        RECT  18.350 1.340 21.890 1.620 ;
        RECT  18.190 0.980 18.350 2.080 ;
        RECT  18.030 0.980 18.190 1.260 ;
        RECT  16.910 1.860 18.190 2.080 ;
        RECT  17.270 0.980 18.030 1.140 ;
        RECT  16.830 1.420 18.030 1.700 ;
        RECT  16.990 0.860 17.270 1.140 ;
        RECT  16.670 0.770 16.830 1.700 ;
        RECT  15.750 0.770 16.670 0.930 ;
        RECT  16.190 2.120 16.230 2.400 ;
        RECT  15.950 1.090 16.190 2.400 ;
        RECT  15.910 1.090 15.950 1.740 ;
        RECT  14.350 1.580 15.910 1.740 ;
        RECT  15.590 0.440 15.750 0.610 ;
        RECT  15.590 0.770 15.750 1.360 ;
        RECT  13.210 0.440 15.590 0.600 ;
        RECT  15.010 1.200 15.590 1.360 ;
        RECT  15.210 0.760 15.430 1.040 ;
        RECT  13.530 0.760 15.210 0.920 ;
        RECT  14.950 1.970 15.110 2.720 ;
        RECT  14.850 1.080 15.010 1.360 ;
        RECT  14.790 1.970 14.950 2.830 ;
        RECT  13.850 1.080 14.850 1.300 ;
        RECT  12.910 2.610 14.790 2.830 ;
        RECT  14.350 1.970 14.630 2.250 ;
        RECT  14.070 1.460 14.350 1.740 ;
        RECT  13.850 1.970 14.350 2.130 ;
        RECT  13.230 2.290 14.150 2.450 ;
        RECT  13.690 1.080 13.850 2.130 ;
        RECT  13.390 1.910 13.690 2.130 ;
        RECT  13.370 0.760 13.530 1.160 ;
        RECT  13.230 0.880 13.370 1.160 ;
        RECT  13.130 0.880 13.230 2.450 ;
        RECT  13.050 0.440 13.210 0.720 ;
        RECT  13.070 1.000 13.130 2.450 ;
        RECT  12.370 1.000 13.070 1.160 ;
        RECT  11.910 0.560 13.050 0.720 ;
        RECT  12.250 0.970 12.370 1.250 ;
        RECT  12.090 0.970 12.250 2.240 ;
        RECT  11.710 2.080 12.090 2.240 ;
        RECT  11.790 1.640 11.930 1.920 ;
        RECT  11.790 0.530 11.910 1.240 ;
        RECT  11.630 0.530 11.790 1.920 ;
        RECT  11.430 2.080 11.710 2.360 ;
        RECT  10.990 1.640 11.630 1.920 ;
        RECT  10.830 0.530 10.990 2.240 ;
        RECT  10.670 0.530 10.830 1.240 ;
        RECT  10.670 2.080 10.830 2.240 ;
        RECT  10.390 2.080 10.670 2.360 ;
        RECT  9.630 2.080 10.390 2.240 ;
        RECT  9.810 0.960 10.030 1.830 ;
        RECT  9.170 1.670 9.810 1.830 ;
        RECT  9.350 2.050 9.630 2.330 ;
        RECT  9.110 0.440 9.330 1.070 ;
        RECT  8.890 1.670 9.170 2.360 ;
        RECT  5.870 0.850 9.110 1.070 ;
        RECT  6.250 0.470 8.910 0.690 ;
        RECT  8.320 1.670 8.890 1.830 ;
        RECT  8.040 1.550 8.320 1.830 ;
        RECT  7.910 2.310 8.190 2.910 ;
        RECT  6.910 2.310 7.910 2.470 ;
        RECT  6.630 2.120 6.910 2.910 ;
        RECT  5.870 2.120 6.630 2.280 ;
        RECT  5.710 0.850 5.870 2.280 ;
        RECT  4.210 1.440 5.710 1.720 ;
        RECT  5.330 0.960 5.550 1.280 ;
        RECT  5.330 1.910 5.550 2.680 ;
        RECT  4.650 1.120 5.330 1.280 ;
        RECT  4.650 1.910 5.330 2.070 ;
        RECT  4.370 0.960 4.650 1.280 ;
        RECT  4.370 1.910 4.650 2.680 ;
        RECT  4.050 1.120 4.370 1.280 ;
        RECT  4.050 1.910 4.370 2.070 ;
        RECT  3.890 1.120 4.050 2.070 ;
        RECT  1.010 1.470 3.890 1.750 ;
    END
END BENCX4TR

MACRO BENCX2TR
    CLASS CORE ;
    FOREIGN BENCX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.800 1.800 12.820 2.080 ;
        RECT  12.640 0.840 12.800 2.080 ;
        RECT  11.440 0.840 12.640 1.120 ;
        RECT  12.440 1.640 12.640 2.080 ;
        RECT  11.560 1.800 12.440 2.080 ;
        END
        ANTENNADIFFAREA 7.596 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.820 1.150 17.920 2.070 ;
        RECT  17.640 0.440 17.820 3.160 ;
        RECT  17.540 0.440 17.640 1.310 ;
        RECT  17.540 1.910 17.640 3.160 ;
        RECT  16.860 1.150 17.540 1.310 ;
        RECT  16.860 1.910 17.540 2.070 ;
        RECT  16.580 0.440 16.860 1.310 ;
        RECT  16.580 1.910 16.860 3.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.440 2.840 14.760 3.160 ;
        RECT  13.840 2.840 14.440 3.000 ;
        RECT  13.720 2.840 13.840 3.160 ;
        RECT  13.560 2.880 13.720 3.160 ;
        RECT  10.880 2.880 13.560 3.040 ;
        RECT  10.720 2.880 10.880 3.160 ;
        RECT  7.780 3.000 10.720 3.160 ;
        RECT  7.620 2.820 7.780 3.160 ;
        RECT  6.050 2.820 7.620 3.040 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.940 2.480 8.160 2.760 ;
        RECT  5.890 2.480 7.940 2.640 ;
        RECT  5.610 2.480 5.890 2.840 ;
        RECT  5.030 2.480 5.610 2.640 ;
        RECT  4.870 2.350 5.030 2.640 ;
        RECT  4.070 2.350 4.870 2.510 ;
        RECT  3.680 1.580 4.070 2.510 ;
        END
        ANTENNAGATEAREA 0.5136 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.700 0.520 6.860 1.320 ;
        RECT  5.390 0.520 6.700 0.680 ;
        RECT  6.580 1.040 6.700 1.320 ;
        RECT  5.230 0.520 5.390 0.920 ;
        RECT  4.870 0.760 5.230 0.920 ;
        RECT  4.710 0.760 4.870 1.400 ;
        RECT  3.520 1.240 4.710 1.400 ;
        RECT  3.490 1.240 3.520 1.560 ;
        RECT  3.270 1.240 3.490 1.690 ;
        END
        ANTENNAGATEAREA 0.5112 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.440 1.810 1.310 ;
        RECT  1.530 1.910 1.810 3.160 ;
        RECT  0.850 1.150 1.530 1.310 ;
        RECT  0.850 1.910 1.530 2.070 ;
        RECT  0.760 0.440 0.850 1.310 ;
        RECT  0.760 1.910 0.850 3.160 ;
        RECT  0.570 0.440 0.760 3.160 ;
        RECT  0.480 1.150 0.570 2.070 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.300 -0.280 18.400 0.280 ;
        RECT  18.080 -0.280 18.300 1.310 ;
        RECT  17.340 -0.280 18.080 0.280 ;
        RECT  17.060 -0.280 17.340 0.990 ;
        RECT  16.340 -0.280 17.060 0.280 ;
        RECT  16.060 -0.280 16.340 0.400 ;
        RECT  15.540 -0.280 16.060 0.280 ;
        RECT  15.260 -0.280 15.540 0.400 ;
        RECT  14.500 -0.280 15.260 0.280 ;
        RECT  14.220 -0.280 14.500 0.340 ;
        RECT  13.320 -0.280 14.220 0.280 ;
        RECT  13.040 -0.280 13.320 0.360 ;
        RECT  12.200 -0.280 13.040 0.280 ;
        RECT  11.920 -0.280 12.200 0.360 ;
        RECT  11.160 -0.280 11.920 0.280 ;
        RECT  10.880 -0.280 11.160 0.360 ;
        RECT  10.040 -0.280 10.880 0.340 ;
        RECT  9.760 -0.280 10.040 0.360 ;
        RECT  7.820 -0.280 9.760 0.280 ;
        RECT  7.540 -0.280 7.820 0.360 ;
        RECT  6.780 -0.280 7.540 0.280 ;
        RECT  6.500 -0.280 6.780 0.360 ;
        RECT  5.530 -0.280 6.500 0.340 ;
        RECT  4.210 -0.280 5.530 0.280 ;
        RECT  3.930 -0.280 4.210 0.320 ;
        RECT  3.170 -0.280 3.930 0.280 ;
        RECT  2.890 -0.280 3.170 0.400 ;
        RECT  2.290 -0.280 2.890 0.280 ;
        RECT  2.010 -0.280 2.290 0.860 ;
        RECT  1.330 -0.280 2.010 0.280 ;
        RECT  1.050 -0.280 1.330 0.990 ;
        RECT  0.310 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.310 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.300 3.320 18.400 3.880 ;
        RECT  18.080 1.910 18.300 3.880 ;
        RECT  17.340 3.320 18.080 3.880 ;
        RECT  17.060 2.230 17.340 3.880 ;
        RECT  16.340 3.320 17.060 3.880 ;
        RECT  16.060 3.200 16.340 3.880 ;
        RECT  15.580 3.320 16.060 3.880 ;
        RECT  15.300 3.200 15.580 3.880 ;
        RECT  14.280 3.320 15.300 3.880 ;
        RECT  14.000 3.200 14.280 3.880 ;
        RECT  13.400 3.320 14.000 3.880 ;
        RECT  13.120 3.200 13.400 3.880 ;
        RECT  12.360 3.320 13.120 3.880 ;
        RECT  12.080 3.200 12.360 3.880 ;
        RECT  11.320 3.320 12.080 3.880 ;
        RECT  11.040 3.200 11.320 3.880 ;
        RECT  7.460 3.320 11.040 3.880 ;
        RECT  7.180 3.200 7.460 3.880 ;
        RECT  6.660 3.320 7.180 3.880 ;
        RECT  6.380 3.200 6.660 3.880 ;
        RECT  5.450 3.320 6.380 3.880 ;
        RECT  5.170 2.800 5.450 3.880 ;
        RECT  4.310 3.320 5.170 3.880 ;
        RECT  4.030 3.200 4.310 3.880 ;
        RECT  3.290 3.320 4.030 3.880 ;
        RECT  3.010 3.200 3.290 3.880 ;
        RECT  2.290 3.320 3.010 3.880 ;
        RECT  2.010 2.120 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.230 1.330 3.880 ;
        RECT  0.310 3.320 1.050 3.880 ;
        RECT  0.090 1.910 0.310 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.380 1.470 17.480 1.750 ;
        RECT  16.060 1.470 16.380 1.630 ;
        RECT  15.980 1.030 16.060 2.070 ;
        RECT  15.900 1.030 15.980 2.690 ;
        RECT  15.660 1.030 15.900 1.310 ;
        RECT  15.700 1.910 15.900 2.690 ;
        RECT  15.280 1.470 15.740 1.750 ;
        RECT  15.120 0.880 15.280 2.560 ;
        RECT  13.880 0.880 15.120 1.160 ;
        RECT  14.840 2.400 15.120 2.680 ;
        RECT  13.680 0.500 15.020 0.720 ;
        RECT  14.680 1.320 14.960 2.240 ;
        RECT  13.880 2.400 14.840 2.560 ;
        RECT  13.120 1.320 14.680 1.480 ;
        RECT  13.460 2.080 14.680 2.240 ;
        RECT  13.140 1.640 14.520 1.920 ;
        RECT  13.660 2.400 13.880 2.680 ;
        RECT  13.520 0.500 13.680 1.160 ;
        RECT  13.400 0.880 13.520 1.160 ;
        RECT  13.300 2.080 13.460 2.720 ;
        RECT  10.560 2.560 13.300 2.720 ;
        RECT  12.980 1.640 13.140 2.400 ;
        RECT  12.960 0.520 13.120 1.480 ;
        RECT  10.240 2.240 12.980 2.400 ;
        RECT  9.340 0.520 12.960 0.680 ;
        RECT  11.200 1.280 12.280 1.560 ;
        RECT  10.800 1.280 11.200 1.440 ;
        RECT  10.640 1.280 10.800 2.080 ;
        RECT  10.520 0.920 10.640 2.080 ;
        RECT  10.400 2.560 10.560 2.840 ;
        RECT  10.360 0.920 10.520 1.440 ;
        RECT  8.320 2.680 10.400 2.840 ;
        RECT  9.920 1.600 10.360 1.880 ;
        RECT  10.080 2.240 10.240 2.520 ;
        RECT  8.480 2.360 10.080 2.520 ;
        RECT  9.760 0.960 9.920 2.200 ;
        RECT  8.860 0.960 9.760 1.120 ;
        RECT  8.800 2.040 9.760 2.200 ;
        RECT  8.440 1.660 9.600 1.880 ;
        RECT  9.060 0.520 9.340 0.800 ;
        RECT  7.300 0.520 9.060 0.680 ;
        RECT  8.580 0.840 8.860 1.120 ;
        RECT  8.320 2.160 8.480 2.520 ;
        RECT  8.220 1.660 8.440 1.820 ;
        RECT  8.220 0.840 8.340 1.120 ;
        RECT  6.090 2.160 8.320 2.320 ;
        RECT  8.060 0.840 8.220 2.000 ;
        RECT  7.700 1.720 8.060 2.000 ;
        RECT  7.300 1.280 7.900 1.560 ;
        RECT  7.180 0.520 7.300 1.560 ;
        RECT  7.140 0.520 7.180 2.000 ;
        RECT  7.020 0.690 7.140 2.000 ;
        RECT  6.780 1.720 7.020 2.000 ;
        RECT  6.090 0.840 6.330 1.120 ;
        RECT  6.050 0.840 6.090 2.320 ;
        RECT  5.930 0.960 6.050 2.320 ;
        RECT  5.810 2.040 5.930 2.320 ;
        RECT  5.190 1.080 5.370 1.300 ;
        RECT  5.030 1.080 5.190 1.730 ;
        RECT  4.530 0.440 5.070 0.600 ;
        RECT  5.010 1.570 5.030 1.730 ;
        RECT  4.730 1.570 5.010 2.190 ;
        RECT  4.230 1.570 4.730 1.790 ;
        RECT  3.470 2.670 4.710 2.890 ;
        RECT  3.110 0.860 4.550 1.080 ;
        RECT  4.370 0.440 4.530 0.700 ;
        RECT  3.410 0.480 4.370 0.700 ;
        RECT  3.310 1.910 3.470 2.890 ;
        RECT  3.190 1.910 3.310 2.700 ;
        RECT  3.110 1.910 3.190 2.070 ;
        RECT  2.950 0.860 3.110 2.070 ;
        RECT  2.290 1.360 2.950 1.640 ;
        RECT  2.650 0.820 2.770 1.100 ;
        RECT  2.650 2.880 2.770 3.160 ;
        RECT  2.490 0.820 2.650 1.180 ;
        RECT  2.490 1.800 2.650 3.160 ;
        RECT  2.130 1.020 2.490 1.180 ;
        RECT  2.130 1.800 2.490 1.960 ;
        RECT  1.970 1.020 2.130 1.960 ;
        RECT  0.920 1.470 1.970 1.750 ;
    END
END BENCX2TR

MACRO BENCX1TR
    CLASS CORE ;
    FOREIGN BENCX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.660 0.840 9.920 1.160 ;
        RECT  9.500 0.840 9.660 2.040 ;
        RECT  9.320 1.880 9.500 2.040 ;
        END
        ANTENNADIFFAREA 3.834 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.280 0.440 13.520 3.160 ;
        RECT  13.200 0.440 13.280 1.310 ;
        RECT  13.200 1.910 13.280 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.500 2.630 10.880 3.160 ;
        RECT  10.480 2.840 10.500 3.160 ;
        RECT  6.260 2.840 10.480 3.000 ;
        RECT  6.100 2.840 6.260 3.160 ;
        RECT  5.600 3.000 6.100 3.160 ;
        RECT  5.440 2.880 5.600 3.160 ;
        RECT  4.620 2.880 5.440 3.040 ;
        RECT  4.430 2.880 4.620 3.160 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.760 2.520 5.940 2.840 ;
        RECT  3.120 2.520 5.760 2.680 ;
        RECT  3.040 2.040 3.120 2.680 ;
        RECT  2.960 1.720 3.040 2.680 ;
        RECT  2.880 1.720 2.960 2.360 ;
        RECT  2.820 1.720 2.880 2.000 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.330 1.190 4.500 1.560 ;
        RECT  2.720 1.400 4.330 1.560 ;
        RECT  2.500 1.240 2.720 1.560 ;
        RECT  2.340 1.240 2.500 1.890 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.440 0.860 1.250 ;
        RECT  0.580 1.880 0.860 3.160 ;
        RECT  0.320 1.090 0.580 1.250 ;
        RECT  0.320 1.880 0.580 2.040 ;
        RECT  0.080 0.840 0.320 2.040 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.900 -0.280 14.000 0.280 ;
        RECT  13.680 -0.280 13.900 1.310 ;
        RECT  12.900 -0.280 13.680 0.280 ;
        RECT  11.880 -0.280 12.900 0.340 ;
        RECT  11.120 -0.280 11.880 0.280 ;
        RECT  10.840 -0.280 11.120 0.340 ;
        RECT  9.240 -0.280 10.840 0.280 ;
        RECT  8.960 -0.280 9.240 0.340 ;
        RECT  8.260 -0.280 8.960 0.280 ;
        RECT  7.980 -0.280 8.260 0.340 ;
        RECT  5.760 -0.280 7.980 0.280 ;
        RECT  5.480 -0.280 5.760 0.340 ;
        RECT  3.840 -0.280 5.480 0.280 ;
        RECT  3.100 -0.280 3.840 0.340 ;
        RECT  2.320 -0.280 3.100 0.280 ;
        RECT  1.330 -0.280 2.320 0.340 ;
        RECT  1.060 -0.280 1.330 0.760 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 0.670 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.900 3.320 14.000 3.880 ;
        RECT  13.680 1.910 13.900 3.880 ;
        RECT  12.900 3.320 13.680 3.880 ;
        RECT  12.620 3.260 12.900 3.880 ;
        RECT  11.320 3.320 12.620 3.880 ;
        RECT  11.040 3.260 11.320 3.880 ;
        RECT  10.120 3.320 11.040 3.880 ;
        RECT  9.840 3.260 10.120 3.880 ;
        RECT  9.080 3.320 9.840 3.880 ;
        RECT  8.800 3.260 9.080 3.880 ;
        RECT  7.970 3.320 8.800 3.880 ;
        RECT  7.690 3.260 7.970 3.880 ;
        RECT  5.280 3.320 7.690 3.880 ;
        RECT  5.000 3.260 5.280 3.880 ;
        RECT  4.260 3.320 5.000 3.880 ;
        RECT  4.020 2.840 4.260 3.880 ;
        RECT  3.180 3.320 4.020 3.880 ;
        RECT  2.900 3.260 3.180 3.880 ;
        RECT  1.380 3.320 2.900 3.880 ;
        RECT  1.100 2.920 1.380 3.880 ;
        RECT  0.410 3.320 1.100 3.880 ;
        RECT  0.100 2.200 0.410 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.000 1.470 13.120 1.630 ;
        RECT  12.840 1.150 13.000 2.070 ;
        RECT  12.440 1.150 12.840 1.310 ;
        RECT  12.440 1.910 12.840 2.070 ;
        RECT  12.100 1.470 12.680 1.630 ;
        RECT  12.280 1.030 12.440 1.310 ;
        RECT  12.280 1.910 12.440 2.690 ;
        RECT  11.940 1.000 12.100 2.470 ;
        RECT  10.840 1.000 11.940 1.160 ;
        RECT  10.460 2.310 11.940 2.470 ;
        RECT  11.620 1.350 11.780 2.150 ;
        RECT  10.240 1.350 11.620 1.510 ;
        RECT  10.300 1.990 11.620 2.150 ;
        RECT  11.420 0.450 11.580 0.730 ;
        RECT  10.650 0.570 11.420 0.730 ;
        RECT  9.980 1.670 11.360 1.830 ;
        RECT  10.400 0.570 10.650 1.190 ;
        RECT  10.140 1.990 10.300 2.680 ;
        RECT  10.080 0.500 10.240 1.510 ;
        RECT  6.100 2.520 10.140 2.680 ;
        RECT  7.180 0.500 10.080 0.660 ;
        RECT  9.820 1.670 9.980 2.360 ;
        RECT  8.280 2.200 9.820 2.360 ;
        RECT  8.720 1.270 9.340 1.550 ;
        RECT  8.660 1.270 8.720 2.040 ;
        RECT  8.500 0.940 8.660 2.040 ;
        RECT  8.440 1.880 8.500 2.040 ;
        RECT  8.120 0.820 8.280 2.360 ;
        RECT  7.500 0.820 8.120 0.980 ;
        RECT  7.710 2.200 8.120 2.360 ;
        RECT  7.800 1.550 7.960 1.860 ;
        RECT  6.900 1.700 7.800 1.860 ;
        RECT  7.340 0.820 7.500 1.420 ;
        RECT  7.120 1.260 7.340 1.420 ;
        RECT  7.160 2.020 7.320 2.360 ;
        RECT  7.020 0.500 7.180 1.100 ;
        RECT  6.160 2.200 7.160 2.360 ;
        RECT  6.960 1.260 7.120 1.540 ;
        RECT  5.150 0.500 7.020 0.660 ;
        RECT  6.780 1.700 6.900 2.040 ;
        RECT  6.620 0.940 6.780 2.040 ;
        RECT  6.480 0.940 6.620 1.100 ;
        RECT  6.160 0.940 6.280 1.100 ;
        RECT  6.050 0.940 6.160 2.360 ;
        RECT  6.000 0.940 6.050 2.330 ;
        RECT  5.540 2.170 6.000 2.330 ;
        RECT  5.160 1.610 5.620 1.770 ;
        RECT  5.150 1.610 5.160 2.240 ;
        RECT  4.990 0.500 5.150 2.240 ;
        RECT  4.720 2.080 4.990 2.240 ;
        RECT  4.660 0.520 4.820 1.920 ;
        RECT  4.560 2.080 4.720 2.360 ;
        RECT  4.190 0.520 4.660 0.680 ;
        RECT  3.680 1.740 4.660 1.920 ;
        RECT  3.680 1.030 3.840 1.190 ;
        RECT  3.480 2.840 3.700 3.120 ;
        RECT  3.520 0.510 3.680 1.190 ;
        RECT  3.520 1.740 3.680 2.360 ;
        RECT  2.560 0.510 3.520 0.670 ;
        RECT  3.280 1.740 3.520 1.900 ;
        RECT  2.300 2.840 3.480 3.000 ;
        RECT  3.080 0.920 3.360 1.190 ;
        RECT  2.180 0.920 3.080 1.080 ;
        RECT  2.180 2.050 2.300 3.000 ;
        RECT  2.140 0.920 2.180 3.000 ;
        RECT  2.020 0.920 2.140 2.210 ;
        RECT  1.560 1.360 2.020 1.640 ;
        RECT  1.400 2.470 1.920 2.630 ;
        RECT  1.680 0.850 1.840 1.130 ;
        RECT  1.400 0.970 1.680 1.130 ;
        RECT  1.240 0.970 1.400 2.630 ;
        RECT  0.580 1.560 1.240 1.720 ;
    END
END BENCX1TR

MACRO BMXIX4TR
    CLASS CORE ;
    FOREIGN BMXIX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.410 2.720 12.510 3.000 ;
        RECT  12.230 2.720 12.410 3.160 ;
        RECT  12.080 2.840 12.230 3.160 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.120 1.240 9.160 1.640 ;
        END
        ANTENNAGATEAREA 0.6312 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.430 1.240 13.520 2.360 ;
        RECT  13.150 0.440 13.430 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.510 7.960 1.960 ;
        RECT  7.580 1.510 7.640 1.790 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 1.210 3.080 2.720 ;
        RECT  0.720 2.560 2.800 2.720 ;
        RECT  0.560 1.640 0.720 2.760 ;
        RECT  0.400 1.640 0.560 1.920 ;
        RECT  0.480 2.440 0.560 2.760 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.640 1.940 1.920 ;
        RECT  0.880 1.640 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.6336 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.910 -0.280 14.000 0.280 ;
        RECT  13.690 -0.280 13.910 1.310 ;
        RECT  12.910 -0.280 13.690 0.280 ;
        RECT  12.630 -0.280 12.910 0.400 ;
        RECT  9.070 -0.280 12.630 0.280 ;
        RECT  8.790 -0.280 9.070 0.320 ;
        RECT  8.030 -0.280 8.790 0.280 ;
        RECT  7.750 -0.280 8.030 0.320 ;
        RECT  1.780 -0.280 7.750 0.280 ;
        RECT  1.500 -0.280 1.780 0.750 ;
        RECT  0.780 -0.280 1.500 0.280 ;
        RECT  0.500 -0.280 0.780 0.400 ;
        RECT  0.000 -0.280 0.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.910 3.320 14.000 3.880 ;
        RECT  13.690 1.910 13.910 3.880 ;
        RECT  12.950 3.320 13.690 3.880 ;
        RECT  12.670 1.910 12.950 3.880 ;
        RECT  9.070 3.320 12.670 3.880 ;
        RECT  8.790 3.260 9.070 3.880 ;
        RECT  8.030 3.320 8.790 3.880 ;
        RECT  7.750 3.260 8.030 3.880 ;
        RECT  1.780 3.320 7.750 3.880 ;
        RECT  1.500 2.880 1.780 3.880 ;
        RECT  0.780 3.320 1.500 3.880 ;
        RECT  0.500 3.180 0.780 3.880 ;
        RECT  0.000 3.320 0.500 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.910 1.470 12.990 1.750 ;
        RECT  12.750 0.560 12.910 1.750 ;
        RECT  11.970 0.560 12.750 0.760 ;
        RECT  12.310 0.970 12.430 1.190 ;
        RECT  12.310 2.000 12.430 2.280 ;
        RECT  12.150 0.970 12.310 2.280 ;
        RECT  11.980 1.510 12.150 1.790 ;
        RECT  11.820 0.560 11.970 0.990 ;
        RECT  11.820 2.490 11.920 2.780 ;
        RECT  11.660 0.560 11.820 2.780 ;
        RECT  11.010 0.560 11.660 0.720 ;
        RECT  11.370 2.010 11.500 2.670 ;
        RECT  11.370 0.920 11.490 1.200 ;
        RECT  11.210 0.920 11.370 3.100 ;
        RECT  7.300 2.940 11.210 3.100 ;
        RECT  10.890 2.180 11.020 2.780 ;
        RECT  10.890 0.560 11.010 0.930 ;
        RECT  10.730 0.560 10.890 2.780 ;
        RECT  10.060 2.620 10.730 2.780 ;
        RECT  10.410 0.610 10.540 2.460 ;
        RECT  10.380 0.480 10.410 2.460 ;
        RECT  10.250 0.480 10.380 0.890 ;
        RECT  10.260 2.180 10.380 2.460 ;
        RECT  6.620 0.480 10.250 0.640 ;
        RECT  9.900 0.880 10.060 2.780 ;
        RECT  9.770 0.880 9.900 1.200 ;
        RECT  9.780 2.180 9.900 2.780 ;
        RECT  9.480 1.910 9.600 2.780 ;
        RECT  9.480 0.920 9.590 1.230 ;
        RECT  9.320 0.920 9.480 2.780 ;
        RECT  8.550 0.920 9.320 1.080 ;
        RECT  8.550 2.620 9.320 2.780 ;
        RECT  8.270 0.800 8.550 1.080 ;
        RECT  8.270 1.910 8.550 2.780 ;
        RECT  7.140 2.620 8.270 2.780 ;
        RECT  7.420 1.030 7.630 1.310 ;
        RECT  7.420 1.930 7.480 2.210 ;
        RECT  7.260 1.030 7.420 2.210 ;
        RECT  7.140 2.940 7.300 3.160 ;
        RECT  7.200 1.530 7.260 2.210 ;
        RECT  7.110 1.530 7.200 1.810 ;
        RECT  6.980 2.500 7.140 2.780 ;
        RECT  3.400 3.000 7.140 3.160 ;
        RECT  6.950 0.980 7.100 1.260 ;
        RECT  6.950 1.970 6.980 2.840 ;
        RECT  6.820 0.980 6.950 2.840 ;
        RECT  6.790 1.100 6.820 2.130 ;
        RECT  5.140 2.680 6.820 2.840 ;
        RECT  6.500 2.240 6.660 2.520 ;
        RECT  6.500 0.480 6.620 0.990 ;
        RECT  6.460 0.480 6.500 2.520 ;
        RECT  6.340 0.710 6.460 2.520 ;
        RECT  5.620 2.360 6.340 2.520 ;
        RECT  6.020 0.710 6.140 0.990 ;
        RECT  6.020 1.920 6.140 2.200 ;
        RECT  5.860 0.440 6.020 2.200 ;
        RECT  4.680 0.440 5.860 0.720 ;
        RECT  5.620 0.980 5.660 1.260 ;
        RECT  5.460 0.980 5.620 2.520 ;
        RECT  5.380 0.980 5.460 1.260 ;
        RECT  5.340 2.240 5.460 2.520 ;
        RECT  5.140 1.030 5.180 1.310 ;
        RECT  4.980 1.030 5.140 2.840 ;
        RECT  4.900 1.030 4.980 1.310 ;
        RECT  4.860 2.560 4.980 2.840 ;
        RECT  3.780 2.680 4.860 2.840 ;
        RECT  4.680 1.910 4.800 2.190 ;
        RECT  4.520 0.440 4.680 2.190 ;
        RECT  2.640 0.440 4.520 0.600 ;
        RECT  4.260 1.030 4.360 1.310 ;
        RECT  4.240 1.030 4.260 2.480 ;
        RECT  4.080 0.770 4.240 2.480 ;
        RECT  3.400 0.770 4.080 0.930 ;
        RECT  3.980 2.200 4.080 2.480 ;
        RECT  3.780 1.090 3.840 1.310 ;
        RECT  3.560 1.090 3.780 2.840 ;
        RECT  3.240 0.770 3.400 3.160 ;
        RECT  3.000 0.770 3.240 1.050 ;
        RECT  2.520 2.880 3.240 3.160 ;
        RECT  2.480 0.440 2.640 2.280 ;
        RECT  2.360 0.440 2.480 1.160 ;
        RECT  2.260 2.120 2.480 2.280 ;
        RECT  1.300 1.000 2.360 1.160 ;
        RECT  2.100 1.320 2.320 1.890 ;
        RECT  1.980 2.120 2.260 2.400 ;
        RECT  0.380 1.320 2.100 1.480 ;
        RECT  1.300 2.120 1.980 2.280 ;
        RECT  1.020 0.440 1.300 1.160 ;
        RECT  1.020 2.120 1.300 2.400 ;
        RECT  0.240 0.880 0.380 1.480 ;
        RECT  0.240 2.080 0.320 2.360 ;
        RECT  0.080 0.880 0.240 2.360 ;
    END
END BMXIX4TR

MACRO BMXIX2TR
    CLASS CORE ;
    FOREIGN BMXIX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.040 2.440 8.360 2.840 ;
        END
        ANTENNAGATEAREA 0.2208 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.240 6.360 1.640 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.360 0.440 9.520 3.160 ;
        RECT  9.130 0.440 9.360 1.310 ;
        RECT  9.110 1.910 9.360 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.240 5.560 1.840 ;
        RECT  5.180 1.560 5.280 1.840 ;
        END
        ANTENNAGATEAREA 0.2208 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.420 1.520 2.580 2.920 ;
        RECT  2.350 1.520 2.420 1.800 ;
        RECT  2.230 2.760 2.420 2.920 ;
        RECT  1.950 2.760 2.230 3.040 ;
        RECT  0.720 2.880 1.950 3.040 ;
        RECT  0.560 1.640 0.720 3.040 ;
        RECT  0.410 1.640 0.560 1.960 ;
        RECT  0.480 2.440 0.560 2.760 ;
        END
        ANTENNAGATEAREA 0.2184 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.890 -0.280 9.600 0.280 ;
        RECT  8.610 -0.280 8.890 0.400 ;
        RECT  6.460 -0.280 8.610 0.340 ;
        RECT  5.380 -0.280 6.460 0.380 ;
        RECT  1.850 -0.280 5.380 0.340 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  0.810 -0.280 1.570 0.340 ;
        RECT  0.530 -0.280 0.810 0.780 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.940 3.320 9.600 3.880 ;
        RECT  8.650 2.020 8.940 3.880 ;
        RECT  6.460 3.260 8.650 3.880 ;
        RECT  5.380 3.200 6.460 3.880 ;
        RECT  1.850 3.260 5.380 3.880 ;
        RECT  1.570 3.200 1.850 3.880 ;
        RECT  0.810 3.260 1.570 3.880 ;
        RECT  0.530 3.200 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.860 1.470 9.130 1.750 ;
        RECT  8.700 0.560 8.860 1.750 ;
        RECT  7.440 0.560 8.700 0.720 ;
        RECT  8.240 0.880 8.380 1.160 ;
        RECT  8.240 2.000 8.340 2.280 ;
        RECT  8.080 0.880 8.240 2.280 ;
        RECT  8.060 1.550 8.080 2.280 ;
        RECT  7.920 1.550 8.060 1.830 ;
        RECT  7.760 0.880 7.920 1.160 ;
        RECT  7.760 1.990 7.880 2.670 ;
        RECT  7.600 0.880 7.760 3.040 ;
        RECT  5.120 2.880 7.600 3.040 ;
        RECT  7.400 0.560 7.440 0.930 ;
        RECT  7.280 0.560 7.400 2.670 ;
        RECT  7.240 0.650 7.280 2.670 ;
        RECT  7.160 0.650 7.240 0.930 ;
        RECT  7.120 2.140 7.240 2.670 ;
        RECT  6.840 0.650 6.960 0.930 ;
        RECT  6.840 2.140 6.920 2.720 ;
        RECT  6.680 0.540 6.840 2.720 ;
        RECT  4.160 0.540 6.680 0.700 ;
        RECT  6.640 2.140 6.680 2.720 ;
        RECT  5.880 0.860 6.060 1.080 ;
        RECT  5.880 1.980 6.060 2.720 ;
        RECT  5.720 0.860 5.880 2.720 ;
        RECT  4.800 2.460 5.720 2.720 ;
        RECT  5.020 2.000 5.140 2.280 ;
        RECT  4.960 2.880 5.120 3.100 ;
        RECT  5.020 0.910 5.100 1.190 ;
        RECT  4.800 0.910 5.020 2.280 ;
        RECT  2.900 2.940 4.960 3.100 ;
        RECT  4.640 2.460 4.800 2.780 ;
        RECT  4.420 0.990 4.640 2.780 ;
        RECT  3.440 2.620 4.420 2.780 ;
        RECT  4.160 2.010 4.260 2.350 ;
        RECT  4.000 0.540 4.160 2.350 ;
        RECT  3.880 0.710 4.000 0.990 ;
        RECT  3.980 2.010 4.000 2.350 ;
        RECT  3.620 1.930 3.780 2.210 ;
        RECT  3.460 0.500 3.620 2.210 ;
        RECT  2.190 0.500 3.460 0.660 ;
        RECT  3.300 2.500 3.440 2.780 ;
        RECT  3.140 0.820 3.300 2.780 ;
        RECT  2.890 0.820 3.140 1.040 ;
        RECT  2.740 1.200 2.900 3.100 ;
        RECT  2.690 1.200 2.740 1.360 ;
        RECT  2.410 1.030 2.690 1.360 ;
        RECT  2.190 2.190 2.260 2.470 ;
        RECT  2.030 0.500 2.190 2.470 ;
        RECT  1.910 0.760 2.030 1.040 ;
        RECT  1.980 2.230 2.030 2.470 ;
        RECT  1.330 2.230 1.980 2.390 ;
        RECT  1.330 0.880 1.910 1.040 ;
        RECT  1.710 1.320 1.870 2.070 ;
        RECT  0.370 1.320 1.710 1.480 ;
        RECT  1.050 0.760 1.330 1.040 ;
        RECT  1.050 2.230 1.330 2.510 ;
        RECT  0.250 1.030 0.370 1.480 ;
        RECT  0.250 2.120 0.320 2.400 ;
        RECT  0.090 1.030 0.250 2.400 ;
    END
END BMXIX2TR

MACRO BMXX4TR
    CLASS CORE ;
    FOREIGN BMXX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.320 2.840 14.850 3.120 ;
        RECT  14.080 2.840 14.320 3.160 ;
        END
        ANTENNAGATEAREA 0.5976 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.360 1.560 9.010 1.840 ;
        RECT  8.080 1.560 8.360 1.960 ;
        END
        ANTENNAGATEAREA 0.6768 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.490 0.440 15.770 3.160 ;
        RECT  15.280 0.640 15.490 1.360 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.530 1.240 7.920 1.610 ;
        END
        ANTENNAGATEAREA 0.4656 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.790 1.250 3.070 2.720 ;
        RECT  0.720 2.560 2.790 2.720 ;
        RECT  0.560 1.640 0.720 2.720 ;
        RECT  0.480 1.640 0.560 2.360 ;
        RECT  0.400 1.640 0.480 1.920 ;
        END
        ANTENNAGATEAREA 0.4704 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.640 1.930 1.920 ;
        RECT  0.880 1.640 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.6816 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.250 -0.280 16.400 0.280 ;
        RECT  15.970 -0.280 16.250 1.310 ;
        RECT  15.250 -0.280 15.970 0.280 ;
        RECT  14.970 -0.280 15.250 0.400 ;
        RECT  11.850 -0.280 14.970 0.280 ;
        RECT  11.570 -0.280 11.850 0.340 ;
        RECT  10.810 -0.280 11.570 0.280 ;
        RECT  10.530 -0.280 10.810 0.320 ;
        RECT  9.770 -0.280 10.530 0.280 ;
        RECT  9.490 -0.280 9.770 0.320 ;
        RECT  8.950 -0.280 9.490 0.280 ;
        RECT  8.670 -0.280 8.950 0.320 ;
        RECT  7.910 -0.280 8.670 0.280 ;
        RECT  7.630 -0.280 7.910 0.320 ;
        RECT  1.770 -0.280 7.630 0.280 ;
        RECT  1.490 -0.280 1.770 0.690 ;
        RECT  0.770 -0.280 1.490 0.280 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.250 3.320 16.400 3.880 ;
        RECT  15.970 1.910 16.250 3.880 ;
        RECT  15.290 3.320 15.970 3.880 ;
        RECT  15.010 1.910 15.290 3.880 ;
        RECT  11.850 3.320 15.010 3.880 ;
        RECT  11.570 3.200 11.850 3.880 ;
        RECT  10.810 3.320 11.570 3.880 ;
        RECT  10.530 3.200 10.810 3.880 ;
        RECT  9.770 3.320 10.530 3.880 ;
        RECT  9.490 3.200 9.770 3.880 ;
        RECT  8.930 3.320 9.490 3.880 ;
        RECT  8.650 3.200 8.930 3.880 ;
        RECT  7.890 3.320 8.650 3.880 ;
        RECT  7.610 3.200 7.890 3.880 ;
        RECT  1.770 3.320 7.610 3.880 ;
        RECT  1.490 2.880 1.770 3.880 ;
        RECT  0.770 3.320 1.490 3.880 ;
        RECT  0.490 3.180 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.120 1.530 15.330 1.750 ;
        RECT  14.960 0.710 15.120 1.750 ;
        RECT  14.270 0.710 14.960 0.870 ;
        RECT  14.610 1.030 14.730 1.310 ;
        RECT  14.610 1.910 14.730 2.680 ;
        RECT  14.450 1.030 14.610 2.680 ;
        RECT  14.270 1.450 14.450 1.730 ;
        RECT  14.110 0.440 14.270 1.140 ;
        RECT  14.110 1.910 14.270 2.680 ;
        RECT  13.950 0.440 14.110 2.680 ;
        RECT  13.310 0.440 13.950 0.600 ;
        RECT  13.670 0.860 13.790 1.140 ;
        RECT  13.670 1.910 13.790 2.890 ;
        RECT  13.510 0.860 13.670 3.160 ;
        RECT  12.330 3.000 13.510 3.160 ;
        RECT  13.190 0.440 13.310 1.140 ;
        RECT  13.190 2.120 13.310 2.840 ;
        RECT  13.030 0.440 13.190 2.840 ;
        RECT  12.350 2.560 13.030 2.720 ;
        RECT  12.670 0.500 12.830 2.400 ;
        RECT  12.550 0.500 12.670 1.140 ;
        RECT  12.550 2.120 12.670 2.400 ;
        RECT  11.370 0.500 12.550 0.660 ;
        RECT  12.190 0.860 12.350 2.720 ;
        RECT  12.170 2.880 12.330 3.160 ;
        RECT  12.070 0.860 12.190 1.140 ;
        RECT  12.070 2.120 12.190 2.720 ;
        RECT  10.330 2.880 12.170 3.040 ;
        RECT  11.210 0.500 11.370 2.720 ;
        RECT  11.050 0.570 11.210 0.850 ;
        RECT  11.050 1.910 11.210 2.720 ;
        RECT  10.770 1.360 11.050 1.640 ;
        RECT  10.650 1.360 10.770 1.520 ;
        RECT  10.490 0.480 10.650 1.520 ;
        RECT  6.570 0.480 10.490 0.640 ;
        RECT  10.170 0.950 10.330 3.040 ;
        RECT  10.010 0.950 10.170 1.230 ;
        RECT  10.010 1.910 10.170 3.040 ;
        RECT  9.850 1.470 10.010 1.750 ;
        RECT  9.690 1.470 9.850 3.040 ;
        RECT  7.290 2.880 9.690 3.040 ;
        RECT  9.330 1.000 9.470 1.280 ;
        RECT  9.330 1.910 9.450 2.280 ;
        RECT  9.190 1.000 9.330 2.280 ;
        RECT  9.170 1.070 9.190 2.280 ;
        RECT  8.430 1.070 9.170 1.230 ;
        RECT  8.410 2.120 9.170 2.280 ;
        RECT  8.150 0.950 8.430 1.230 ;
        RECT  8.130 2.120 8.410 2.720 ;
        RECT  7.130 2.560 8.130 2.720 ;
        RECT  7.370 0.800 7.510 1.080 ;
        RECT  7.370 1.910 7.480 2.190 ;
        RECT  7.210 0.800 7.370 2.190 ;
        RECT  7.130 2.880 7.290 3.160 ;
        RECT  7.200 1.480 7.210 2.190 ;
        RECT  7.050 1.480 7.200 1.760 ;
        RECT  6.970 2.440 7.130 2.720 ;
        RECT  3.390 3.000 7.130 3.160 ;
        RECT  6.890 0.980 7.050 1.260 ;
        RECT  6.890 1.920 6.970 2.840 ;
        RECT  6.810 0.980 6.890 2.840 ;
        RECT  6.770 0.980 6.810 2.080 ;
        RECT  5.130 2.680 6.810 2.840 ;
        RECT  6.730 1.100 6.770 2.080 ;
        RECT  6.450 2.240 6.650 2.520 ;
        RECT  6.450 0.480 6.570 0.990 ;
        RECT  6.410 0.480 6.450 2.520 ;
        RECT  6.290 0.710 6.410 2.520 ;
        RECT  5.610 2.360 6.290 2.520 ;
        RECT  5.970 1.920 6.130 2.200 ;
        RECT  5.970 0.660 6.090 0.990 ;
        RECT  5.810 0.660 5.970 2.200 ;
        RECT  4.790 0.660 5.810 0.820 ;
        RECT  5.450 0.980 5.610 2.520 ;
        RECT  5.330 0.980 5.450 1.260 ;
        RECT  5.330 2.240 5.450 2.520 ;
        RECT  4.970 1.020 5.130 2.840 ;
        RECT  4.850 1.020 4.970 1.310 ;
        RECT  4.850 2.560 4.970 2.840 ;
        RECT  3.830 2.680 4.850 2.840 ;
        RECT  4.670 0.440 4.790 0.820 ;
        RECT  4.670 1.920 4.790 2.200 ;
        RECT  4.510 0.440 4.670 2.200 ;
        RECT  2.630 0.440 4.510 0.600 ;
        RECT  4.190 1.030 4.350 1.310 ;
        RECT  4.190 2.240 4.310 2.520 ;
        RECT  4.030 0.770 4.190 2.520 ;
        RECT  3.390 0.770 4.030 0.930 ;
        RECT  3.550 1.090 3.830 2.840 ;
        RECT  3.230 0.770 3.390 3.160 ;
        RECT  2.990 0.770 3.230 1.050 ;
        RECT  2.550 2.880 3.230 3.160 ;
        RECT  2.470 0.440 2.630 2.280 ;
        RECT  2.350 0.440 2.470 1.160 ;
        RECT  2.250 2.120 2.470 2.280 ;
        RECT  1.290 1.000 2.350 1.160 ;
        RECT  2.090 1.320 2.310 1.930 ;
        RECT  1.970 2.120 2.250 2.400 ;
        RECT  0.370 1.320 2.090 1.480 ;
        RECT  1.290 2.120 1.970 2.280 ;
        RECT  1.010 0.440 1.290 1.160 ;
        RECT  1.010 2.120 1.290 2.400 ;
        RECT  0.240 0.920 0.370 1.480 ;
        RECT  0.240 2.080 0.310 2.360 ;
        RECT  0.080 0.920 0.240 2.360 ;
    END
END BMXX4TR

MACRO BMXX2TR
    CLASS CORE ;
    FOREIGN BMXX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 2.670 9.560 3.160 ;
        END
        ANTENNAGATEAREA 0.3 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.480 0.840 6.720 1.640 ;
        RECT  6.400 1.360 6.480 1.640 ;
        END
        ANTENNAGATEAREA 0.3384 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.560 0.440 10.720 3.160 ;
        RECT  10.340 0.440 10.560 1.310 ;
        RECT  10.300 1.910 10.560 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 1.240 5.920 1.700 ;
        RECT  5.420 1.420 5.640 1.700 ;
        END
        ANTENNAGATEAREA 0.24 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.460 1.460 2.620 2.920 ;
        RECT  2.350 1.460 2.460 1.740 ;
        RECT  2.270 2.760 2.460 2.920 ;
        RECT  1.990 2.760 2.270 3.040 ;
        RECT  0.720 2.880 1.990 3.040 ;
        RECT  0.560 1.640 0.720 3.040 ;
        RECT  0.470 1.640 0.560 1.960 ;
        RECT  0.480 2.440 0.560 2.760 ;
        END
        ANTENNAGATEAREA 0.24 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.3384 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.100 -0.280 10.800 0.280 ;
        RECT  9.820 -0.280 10.100 0.400 ;
        RECT  7.720 -0.280 9.820 0.340 ;
        RECT  7.440 -0.280 7.720 0.360 ;
        RECT  5.620 -0.280 7.440 0.340 ;
        RECT  1.850 -0.280 5.620 0.280 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  0.810 -0.280 1.570 0.340 ;
        RECT  0.530 -0.280 0.810 0.760 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.100 3.320 10.800 3.880 ;
        RECT  9.820 2.320 10.100 3.880 ;
        RECT  7.680 3.320 9.820 3.880 ;
        RECT  7.400 2.890 7.680 3.880 ;
        RECT  6.700 3.320 7.400 3.880 ;
        RECT  5.620 3.200 6.700 3.880 ;
        RECT  1.850 3.260 5.620 3.880 ;
        RECT  1.570 3.200 1.850 3.880 ;
        RECT  0.810 3.260 1.570 3.880 ;
        RECT  0.530 3.200 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.180 1.470 10.340 1.750 ;
        RECT  10.020 0.560 10.180 1.750 ;
        RECT  9.600 0.560 10.020 0.720 ;
        RECT  9.600 0.880 9.740 1.160 ;
        RECT  9.600 2.180 9.620 2.460 ;
        RECT  9.440 0.550 9.600 0.720 ;
        RECT  9.440 0.880 9.600 2.460 ;
        RECT  8.740 0.550 9.440 0.710 ;
        RECT  9.340 1.540 9.440 2.460 ;
        RECT  9.220 1.540 9.340 1.820 ;
        RECT  9.060 0.870 9.280 1.150 ;
        RECT  9.060 1.980 9.120 2.730 ;
        RECT  8.900 0.870 9.060 2.730 ;
        RECT  7.200 2.570 8.900 2.730 ;
        RECT  8.640 0.550 8.740 0.870 ;
        RECT  8.580 0.550 8.640 2.410 ;
        RECT  8.480 0.590 8.580 2.410 ;
        RECT  8.360 2.130 8.480 2.410 ;
        RECT  8.200 0.590 8.320 1.310 ;
        RECT  8.040 0.590 8.200 2.410 ;
        RECT  7.880 2.130 8.040 2.410 ;
        RECT  7.820 1.380 7.880 1.660 ;
        RECT  7.660 0.520 7.820 1.660 ;
        RECT  4.400 0.520 7.660 0.680 ;
        RECT  7.340 1.150 7.500 2.290 ;
        RECT  7.200 1.150 7.340 1.310 ;
        RECT  7.200 2.130 7.340 2.290 ;
        RECT  6.920 1.030 7.200 1.310 ;
        RECT  6.920 2.130 7.200 3.160 ;
        RECT  7.060 1.590 7.180 1.870 ;
        RECT  6.900 1.590 7.060 1.960 ;
        RECT  6.620 1.800 6.900 1.960 ;
        RECT  6.460 1.800 6.620 3.040 ;
        RECT  5.300 2.880 6.460 3.040 ;
        RECT  6.240 0.920 6.300 1.200 ;
        RECT  6.240 1.910 6.300 2.720 ;
        RECT  6.080 0.920 6.240 2.720 ;
        RECT  4.980 2.500 6.080 2.720 ;
        RECT  5.260 2.080 5.380 2.240 ;
        RECT  5.260 0.980 5.340 1.260 ;
        RECT  5.140 2.880 5.300 3.100 ;
        RECT  5.040 0.980 5.260 2.240 ;
        RECT  3.000 2.940 5.140 3.100 ;
        RECT  4.880 2.500 4.980 2.780 ;
        RECT  4.660 1.030 4.880 2.780 ;
        RECT  3.480 2.620 4.660 2.780 ;
        RECT  4.400 2.120 4.500 2.420 ;
        RECT  4.240 0.520 4.400 2.420 ;
        RECT  3.970 0.790 4.240 1.120 ;
        RECT  4.220 2.120 4.240 2.420 ;
        RECT  3.640 1.910 4.020 2.190 ;
        RECT  3.640 0.710 3.700 0.990 ;
        RECT  3.480 0.440 3.640 2.190 ;
        RECT  2.190 0.440 3.480 0.600 ;
        RECT  3.320 2.500 3.480 2.780 ;
        RECT  3.160 0.760 3.320 2.780 ;
        RECT  2.890 0.760 3.160 0.980 ;
        RECT  2.780 1.140 3.000 3.100 ;
        RECT  2.690 1.140 2.780 1.300 ;
        RECT  2.410 1.020 2.690 1.300 ;
        RECT  2.190 2.130 2.300 2.410 ;
        RECT  2.030 0.440 2.190 2.410 ;
        RECT  1.910 0.720 2.030 1.000 ;
        RECT  2.020 2.220 2.030 2.410 ;
        RECT  1.330 2.220 2.020 2.380 ;
        RECT  1.330 0.840 1.910 1.000 ;
        RECT  1.650 1.320 1.870 2.060 ;
        RECT  0.370 1.320 1.650 1.480 ;
        RECT  1.050 0.720 1.330 1.000 ;
        RECT  1.050 2.220 1.330 2.500 ;
        RECT  0.250 1.030 0.370 1.480 ;
        RECT  0.250 2.120 0.320 2.400 ;
        RECT  0.090 1.030 0.250 2.400 ;
    END
END BMXX2TR

MACRO OR4XLTR
    CLASS CORE ;
    FOREIGN OR4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.440 2.720 2.660 ;
        RECT  2.460 2.320 2.480 2.660 ;
        END
        ANTENNADIFFAREA 1.12 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.280 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.620 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.640 0.720 2.200 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 -0.280 2.800 0.280 ;
        RECT  2.030 -0.280 2.310 0.620 ;
        RECT  1.240 -0.280 2.030 0.280 ;
        RECT  0.180 -0.280 1.240 0.380 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 3.320 2.800 3.880 ;
        RECT  2.000 2.380 2.260 3.880 ;
        RECT  0.000 3.320 2.000 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.720 2.320 2.000 ;
        RECT  1.680 1.720 1.840 2.540 ;
        RECT  1.640 0.440 1.760 0.720 ;
        RECT  0.320 2.380 1.680 2.540 ;
        RECT  1.480 0.440 1.640 1.080 ;
        RECT  0.860 0.920 1.480 1.080 ;
        RECT  0.530 0.800 0.860 1.080 ;
        RECT  0.320 0.910 0.530 1.080 ;
        RECT  0.160 0.910 0.320 2.540 ;
    END
END OR4XLTR

MACRO OR4X8TR
    CLASS CORE ;
    FOREIGN OR4X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.640 0.440 6.920 2.820 ;
        RECT  5.960 1.040 6.640 1.760 ;
        RECT  5.740 0.440 5.960 3.160 ;
        RECT  5.680 0.440 5.740 1.310 ;
        RECT  5.680 1.910 5.740 3.160 ;
        END
        ANTENNADIFFAREA 7.784 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.080 1.680 5.200 1.960 ;
        RECT  4.920 1.680 5.080 2.620 ;
        RECT  1.960 2.460 4.920 2.620 ;
        RECT  1.680 1.740 1.960 2.620 ;
        END
        ANTENNAGATEAREA 0.5736 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 1.360 4.720 1.960 ;
        RECT  4.480 1.360 4.640 2.300 ;
        RECT  2.560 2.140 4.480 2.300 ;
        RECT  2.400 1.420 2.560 2.300 ;
        RECT  1.200 1.420 2.400 1.580 ;
        END
        ANTENNAGATEAREA 0.5736 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.240 4.320 1.640 ;
        RECT  4.040 1.240 4.200 1.980 ;
        RECT  3.000 1.820 4.040 1.980 ;
        RECT  2.880 1.360 3.000 1.980 ;
        RECT  2.840 1.100 2.880 1.980 ;
        RECT  2.720 1.100 2.840 1.640 ;
        RECT  1.160 1.100 2.720 1.260 ;
        RECT  0.880 0.960 1.160 1.260 ;
        END
        ANTENNAGATEAREA 0.5736 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.380 3.840 1.660 ;
        RECT  3.240 1.240 3.560 1.660 ;
        END
        ANTENNAGATEAREA 0.5736 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.400 -0.280 7.600 0.280 ;
        RECT  7.120 -0.280 7.400 1.310 ;
        RECT  6.440 -0.280 7.120 0.280 ;
        RECT  6.160 -0.280 6.440 0.670 ;
        RECT  5.440 -0.280 6.160 0.280 ;
        RECT  4.240 -0.280 5.440 0.340 ;
        RECT  3.720 -0.280 4.240 0.280 ;
        RECT  3.440 -0.280 3.720 0.340 ;
        RECT  2.680 -0.280 3.440 0.280 ;
        RECT  2.400 -0.280 2.680 0.620 ;
        RECT  1.680 -0.280 2.400 0.280 ;
        RECT  1.400 -0.280 1.680 0.940 ;
        RECT  0.000 -0.280 1.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.400 3.320 7.600 3.880 ;
        RECT  7.120 1.910 7.400 3.880 ;
        RECT  6.440 3.320 7.120 3.880 ;
        RECT  6.160 2.180 6.440 3.880 ;
        RECT  5.440 3.320 6.160 3.880 ;
        RECT  5.160 3.180 5.440 3.880 ;
        RECT  2.040 3.320 5.160 3.880 ;
        RECT  1.760 3.180 2.040 3.880 ;
        RECT  0.000 3.320 1.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.520 1.470 5.580 1.750 ;
        RECT  5.360 0.900 5.520 2.940 ;
        RECT  5.040 0.900 5.360 1.060 ;
        RECT  3.800 2.780 5.360 2.940 ;
        RECT  4.760 0.780 5.040 1.060 ;
        RECT  4.120 0.900 4.760 1.060 ;
        RECT  3.840 0.780 4.120 1.060 ;
        RECT  1.880 0.780 3.840 0.940 ;
        RECT  3.240 2.780 3.800 3.060 ;
        RECT  0.560 2.780 3.240 2.940 ;
        RECT  0.280 2.030 0.560 3.160 ;
    END
END OR4X8TR

MACRO OR4X6TR
    CLASS CORE ;
    FOREIGN OR4X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.130 0.440 5.410 2.950 ;
        RECT  4.450 1.040 5.130 1.760 ;
        RECT  4.230 0.540 4.450 3.160 ;
        RECT  4.170 0.540 4.230 1.310 ;
        RECT  4.170 1.910 4.230 3.160 ;
        END
        ANTENNADIFFAREA 7.132 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 1.560 3.690 2.720 ;
        RECT  0.820 2.560 3.410 2.720 ;
        RECT  0.660 1.720 0.820 2.720 ;
        RECT  0.510 1.720 0.660 1.960 ;
        RECT  0.320 1.550 0.510 1.960 ;
        RECT  0.080 0.830 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.240 3.250 1.520 ;
        RECT  2.970 1.240 3.130 2.400 ;
        RECT  1.140 2.240 2.970 2.400 ;
        RECT  0.980 1.240 1.140 2.400 ;
        RECT  0.770 1.240 0.980 1.560 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.240 2.810 1.560 ;
        RECT  2.440 1.240 2.600 2.080 ;
        RECT  1.520 1.920 2.440 2.080 ;
        RECT  1.300 1.240 1.520 2.080 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.480 2.130 1.760 ;
        RECT  1.680 1.240 1.960 1.760 ;
        END
        ANTENNAGATEAREA 0.4416 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 -0.280 5.600 0.280 ;
        RECT  4.650 -0.280 4.930 0.670 ;
        RECT  3.930 -0.280 4.650 0.280 ;
        RECT  2.730 -0.280 3.930 0.340 ;
        RECT  0.000 -0.280 2.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 3.320 5.600 3.880 ;
        RECT  4.650 2.230 4.930 3.880 ;
        RECT  3.930 3.320 4.650 3.880 ;
        RECT  3.650 3.200 3.930 3.880 ;
        RECT  0.500 3.320 3.650 3.880 ;
        RECT  0.220 2.120 0.500 3.880 ;
        RECT  0.000 3.320 0.220 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.010 1.470 4.070 1.750 ;
        RECT  3.850 0.920 4.010 3.040 ;
        RECT  3.530 0.920 3.850 1.080 ;
        RECT  2.160 2.880 3.850 3.040 ;
        RECT  3.250 0.800 3.530 1.080 ;
        RECT  2.610 0.920 3.250 1.080 ;
        RECT  2.330 0.800 2.610 1.080 ;
        RECT  1.690 0.920 2.330 1.080 ;
        RECT  1.860 2.880 2.160 3.160 ;
        RECT  1.410 0.800 1.690 1.080 ;
        RECT  0.770 0.920 1.410 1.080 ;
        RECT  0.490 0.800 0.770 1.080 ;
    END
END OR4X6TR

MACRO OR4X4TR
    CLASS CORE ;
    FOREIGN OR4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.030 3.920 2.240 ;
        RECT  3.680 0.550 3.830 3.160 ;
        RECT  3.550 0.550 3.680 1.390 ;
        RECT  3.550 1.990 3.680 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.840 3.070 2.120 ;
        RECT  2.850 1.840 3.010 2.600 ;
        RECT  0.320 2.440 2.850 2.600 ;
        RECT  0.080 1.640 0.320 2.770 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.180 2.700 1.460 ;
        RECT  2.480 1.180 2.640 2.280 ;
        RECT  0.830 2.120 2.480 2.280 ;
        RECT  0.670 1.240 0.830 2.280 ;
        RECT  0.480 1.240 0.670 1.560 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.560 ;
        RECT  1.270 1.240 2.080 1.400 ;
        RECT  0.990 1.240 1.270 1.600 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.640 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 -0.280 4.400 0.280 ;
        RECT  4.030 -0.280 4.310 0.750 ;
        RECT  3.350 -0.280 4.030 0.280 ;
        RECT  3.070 -0.280 3.350 0.610 ;
        RECT  2.390 -0.280 3.070 0.280 ;
        RECT  2.110 -0.280 2.390 0.610 ;
        RECT  1.430 -0.280 2.110 0.280 ;
        RECT  1.150 -0.280 1.430 1.010 ;
        RECT  0.000 -0.280 1.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.400 3.880 ;
        RECT  4.030 2.490 4.310 3.880 ;
        RECT  3.310 3.320 4.030 3.880 ;
        RECT  3.030 3.180 3.310 3.880 ;
        RECT  0.390 3.310 3.030 3.880 ;
        RECT  0.110 3.200 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.390 1.550 3.460 1.830 ;
        RECT  3.230 0.860 3.390 2.920 ;
        RECT  2.860 0.860 3.230 1.020 ;
        RECT  1.830 2.760 3.230 2.920 ;
        RECT  2.590 0.450 2.860 1.020 ;
        RECT  1.910 0.860 2.590 1.020 ;
        RECT  1.620 0.450 1.910 1.020 ;
        RECT  1.550 2.760 1.830 3.040 ;
    END
END OR4X4TR

MACRO OR4X2TR
    CLASS CORE ;
    FOREIGN OR4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.440 2.720 2.360 ;
        RECT  2.480 0.440 2.700 3.100 ;
        RECT  2.420 0.440 2.480 1.220 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 2.040 2.320 2.360 ;
        RECT  1.720 1.740 1.880 2.360 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.560 ;
        RECT  1.380 1.240 1.640 1.520 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.200 1.220 1.560 ;
        RECT  0.880 1.200 1.060 1.580 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.740 0.860 2.020 ;
        RECT  0.440 1.640 0.720 2.020 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.320 2.800 3.880 ;
        RECT  1.940 2.650 2.220 3.880 ;
        RECT  0.000 3.320 1.940 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.240 1.420 2.320 1.700 ;
        RECT  2.080 0.880 2.240 1.700 ;
        RECT  1.780 0.880 2.080 1.040 ;
        RECT  1.500 0.760 1.780 1.040 ;
        RECT  0.860 0.880 1.500 1.040 ;
        RECT  0.580 0.760 0.860 1.040 ;
        RECT  0.380 2.180 0.660 3.010 ;
        RECT  0.280 0.880 0.580 1.040 ;
        RECT  0.280 2.180 0.380 2.340 ;
        RECT  0.120 0.880 0.280 2.340 ;
    END
END OR4X2TR

MACRO OR4X1TR
    CLASS CORE ;
    FOREIGN OR4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.530 0.440 2.720 2.660 ;
        RECT  2.480 0.440 2.530 1.560 ;
        RECT  2.460 2.320 2.530 2.660 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.280 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.640 0.720 2.200 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.280 2.800 0.280 ;
        RECT  0.180 -0.280 1.240 0.380 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 3.320 2.800 3.880 ;
        RECT  2.000 2.480 2.260 3.880 ;
        RECT  0.000 3.320 2.000 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.720 2.320 2.000 ;
        RECT  1.680 1.720 1.840 2.540 ;
        RECT  1.480 0.440 1.760 1.080 ;
        RECT  0.320 2.380 1.680 2.540 ;
        RECT  0.860 0.920 1.480 1.080 ;
        RECT  0.530 0.800 0.860 1.080 ;
        RECT  0.320 0.910 0.530 1.080 ;
        RECT  0.160 0.910 0.320 2.540 ;
    END
END OR4X1TR

MACRO OR3XLTR
    CLASS CORE ;
    FOREIGN OR3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.030 2.320 3.160 ;
        RECT  2.060 1.030 2.160 1.310 ;
        RECT  2.080 2.040 2.160 3.160 ;
        RECT  1.940 2.040 2.080 2.390 ;
        END
        ANTENNADIFFAREA 1.174 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.560 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.440 1.120 3.020 ;
        RECT  0.790 2.860 0.880 3.020 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.640 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.280 2.400 0.280 ;
        RECT  1.590 -0.280 1.880 0.730 ;
        RECT  0.830 -0.280 1.590 0.280 ;
        RECT  0.550 -0.280 0.830 0.800 ;
        RECT  0.000 -0.280 0.550 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.320 2.400 3.880 ;
        RECT  1.460 2.190 1.740 3.880 ;
        RECT  0.000 3.320 1.460 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.880 1.480 2.000 1.780 ;
        RECT  1.720 1.060 1.880 1.780 ;
        RECT  1.290 1.060 1.720 1.240 ;
        RECT  1.080 0.520 1.290 1.240 ;
        RECT  1.010 0.520 1.080 2.280 ;
        RECT  0.920 1.090 1.010 2.280 ;
        RECT  0.110 1.090 0.920 1.250 ;
        RECT  0.580 2.120 0.920 2.280 ;
        RECT  0.290 2.120 0.580 2.400 ;
    END
END OR3XLTR

MACRO OR3X8TR
    CLASS CORE ;
    FOREIGN OR3X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.300 0.440 5.320 1.870 ;
        RECT  5.140 0.440 5.300 3.160 ;
        RECT  4.340 1.040 5.140 1.950 ;
        RECT  4.180 0.440 4.340 3.160 ;
        END
        ANTENNADIFFAREA 7.92 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.000 3.580 1.480 ;
        RECT  1.560 1.000 3.420 1.160 ;
        RECT  1.520 1.000 1.560 1.480 ;
        RECT  1.280 0.840 1.520 1.480 ;
        END
        ANTENNAGATEAREA 0.5592 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.190 1.640 3.330 1.800 ;
        RECT  3.030 1.320 3.190 1.800 ;
        RECT  1.880 1.320 3.030 1.480 ;
        RECT  1.720 1.320 1.880 1.800 ;
        RECT  1.120 1.640 1.720 1.800 ;
        RECT  0.870 1.240 1.120 1.800 ;
        RECT  0.720 1.640 0.870 1.800 ;
        END
        ANTENNAGATEAREA 0.5592 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.640 2.720 1.800 ;
        RECT  2.040 1.640 2.200 2.120 ;
        RECT  0.560 1.960 2.040 2.120 ;
        RECT  0.320 1.600 0.560 2.120 ;
        RECT  0.080 0.840 0.320 2.120 ;
        END
        ANTENNAGATEAREA 0.5592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.840 -0.280 6.000 0.280 ;
        RECT  5.560 -0.280 5.840 1.310 ;
        RECT  4.880 -0.280 5.560 0.280 ;
        RECT  4.590 -0.280 4.880 0.670 ;
        RECT  3.880 -0.280 4.590 0.280 ;
        RECT  3.600 -0.280 3.880 0.340 ;
        RECT  2.840 -0.280 3.600 0.280 ;
        RECT  2.560 -0.280 2.840 0.340 ;
        RECT  1.800 -0.280 2.560 0.280 ;
        RECT  1.520 -0.280 1.800 0.340 ;
        RECT  0.740 -0.280 1.520 0.280 ;
        RECT  0.530 -0.280 0.740 1.010 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.850 3.320 6.000 3.880 ;
        RECT  5.530 1.910 5.850 3.880 ;
        RECT  4.900 3.320 5.530 3.880 ;
        RECT  4.590 2.110 4.900 3.880 ;
        RECT  3.940 3.320 4.590 3.880 ;
        RECT  3.630 2.430 3.940 3.880 ;
        RECT  1.600 3.320 3.630 3.880 ;
        RECT  1.320 2.660 1.600 3.880 ;
        RECT  0.000 3.320 1.320 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.900 1.410 3.980 1.690 ;
        RECT  3.740 0.680 3.900 2.120 ;
        RECT  3.300 0.680 3.740 0.840 ;
        RECT  2.700 1.960 3.740 2.120 ;
        RECT  3.140 0.560 3.300 0.840 ;
        RECT  2.260 0.680 3.140 0.840 ;
        RECT  2.460 1.960 2.700 2.690 ;
        RECT  0.340 2.290 2.460 2.450 ;
        RECT  2.100 0.500 2.260 0.840 ;
        RECT  1.000 0.500 2.100 0.660 ;
        RECT  0.180 2.290 0.340 2.660 ;
    END
END OR3X8TR

MACRO OR3X6TR
    CLASS CORE ;
    FOREIGN OR3X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.190 0.500 4.310 1.370 ;
        RECT  4.010 0.500 4.190 2.980 ;
        RECT  3.910 1.040 4.010 2.980 ;
        RECT  3.480 1.040 3.910 2.350 ;
        RECT  3.330 1.040 3.480 1.380 ;
        RECT  3.230 1.980 3.480 2.350 ;
        RECT  3.050 0.440 3.330 1.380 ;
        RECT  3.010 1.980 3.230 3.160 ;
        END
        ANTENNADIFFAREA 6.992 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.590 2.530 2.280 ;
        RECT  0.570 2.120 2.250 2.280 ;
        RECT  0.320 1.640 0.570 2.280 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.320 2.090 1.710 ;
        RECT  0.890 1.320 1.810 1.480 ;
        RECT  0.630 0.840 0.890 1.480 ;
        RECT  0.480 0.840 0.630 1.160 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.640 1.640 1.960 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.810 -0.280 4.400 0.280 ;
        RECT  3.530 -0.280 3.810 0.670 ;
        RECT  2.850 -0.280 3.530 0.280 ;
        RECT  2.570 -0.280 2.850 0.670 ;
        RECT  1.890 -0.280 2.570 0.280 ;
        RECT  1.610 -0.280 1.890 0.670 ;
        RECT  0.000 -0.280 1.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.710 3.320 4.400 3.880 ;
        RECT  3.430 2.700 3.710 3.880 ;
        RECT  2.730 3.320 3.430 3.880 ;
        RECT  2.450 2.930 2.730 3.880 ;
        RECT  0.370 3.320 2.450 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 1.540 3.190 1.820 ;
        RECT  2.690 1.000 2.850 2.600 ;
        RECT  2.370 1.000 2.690 1.160 ;
        RECT  1.490 2.440 2.690 2.600 ;
        RECT  2.090 0.440 2.370 1.160 ;
        RECT  1.410 1.000 2.090 1.160 ;
        RECT  1.210 2.440 1.490 3.160 ;
        RECT  1.130 0.500 1.410 1.160 ;
    END
END OR3X6TR

MACRO OR3X4TR
    CLASS CORE ;
    FOREIGN OR3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.390 1.040 3.520 2.070 ;
        RECT  3.250 0.440 3.390 3.160 ;
        RECT  3.170 0.440 3.250 1.290 ;
        RECT  3.170 1.910 3.250 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.580 2.490 2.280 ;
        RECT  0.720 2.120 2.300 2.280 ;
        RECT  0.470 1.640 0.720 2.280 ;
        RECT  0.260 1.640 0.470 1.930 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.240 2.030 1.420 ;
        RECT  0.880 1.240 1.120 1.600 ;
        RECT  0.590 1.240 0.880 1.420 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.640 1.800 1.960 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.280 4.000 0.280 ;
        RECT  3.590 -0.280 3.870 0.760 ;
        RECT  2.870 -0.280 3.590 0.280 ;
        RECT  2.590 -0.280 2.870 0.690 ;
        RECT  1.910 -0.280 2.590 0.280 ;
        RECT  1.630 -0.280 1.910 0.690 ;
        RECT  0.000 -0.280 1.630 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 3.320 4.000 3.880 ;
        RECT  3.590 2.230 3.870 3.880 ;
        RECT  2.870 3.320 3.590 3.880 ;
        RECT  2.570 2.840 2.870 3.880 ;
        RECT  0.540 3.260 2.570 3.880 ;
        RECT  0.210 2.580 0.540 3.880 ;
        RECT  0.000 3.320 0.210 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.990 1.470 3.070 1.750 ;
        RECT  2.830 0.880 2.990 2.600 ;
        RECT  2.390 0.880 2.830 1.040 ;
        RECT  1.630 2.440 2.830 2.600 ;
        RECT  2.110 0.560 2.390 1.040 ;
        RECT  1.430 0.880 2.110 1.040 ;
        RECT  1.350 2.440 1.630 2.720 ;
        RECT  1.150 0.500 1.430 1.040 ;
    END
END OR3X4TR

MACRO OR3X2TR
    CLASS CORE ;
    FOREIGN OR3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 0.440 2.720 1.560 ;
        RECT  2.520 0.440 2.640 2.070 ;
        RECT  2.480 0.440 2.520 3.100 ;
        RECT  2.400 0.440 2.480 1.310 ;
        RECT  2.240 1.910 2.480 3.100 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.530 1.920 2.000 ;
        RECT  1.550 1.720 1.680 2.000 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.240 1.520 1.560 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.240 0.760 1.560 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 -0.280 2.800 0.280 ;
        RECT  1.880 -0.280 2.160 0.760 ;
        RECT  1.120 -0.280 1.880 0.280 ;
        RECT  0.840 -0.280 1.120 0.640 ;
        RECT  0.000 -0.280 0.840 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 3.320 2.800 3.880 ;
        RECT  1.720 2.280 2.000 3.880 ;
        RECT  0.000 3.320 1.720 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.240 1.470 2.320 1.750 ;
        RECT  2.080 0.920 2.240 1.750 ;
        RECT  1.640 0.920 2.080 1.080 ;
        RECT  1.080 0.800 1.640 1.080 ;
        RECT  0.920 0.800 1.080 2.210 ;
        RECT  0.320 0.800 0.920 1.080 ;
        RECT  0.840 2.050 0.920 2.210 ;
        RECT  0.560 2.050 0.840 2.850 ;
    END
END OR3X2TR

MACRO OR3X1TR
    CLASS CORE ;
    FOREIGN OR3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.950 2.320 3.160 ;
        RECT  2.070 0.950 2.160 1.210 ;
        RECT  2.080 2.040 2.160 3.160 ;
        RECT  1.940 2.040 2.080 2.520 ;
        END
        ANTENNADIFFAREA 1.829 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.560 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.780 1.160 3.160 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.640 0.760 1.960 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.890 -0.280 2.400 0.280 ;
        RECT  1.600 -0.280 1.890 0.550 ;
        RECT  0.840 -0.280 1.600 0.280 ;
        RECT  0.560 -0.280 0.840 0.800 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.740 3.320 2.400 3.880 ;
        RECT  1.460 2.210 1.740 3.880 ;
        RECT  0.000 3.320 1.460 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.880 1.480 2.000 1.780 ;
        RECT  1.720 1.060 1.880 1.780 ;
        RECT  1.300 1.060 1.720 1.240 ;
        RECT  1.080 0.520 1.300 1.240 ;
        RECT  1.020 0.520 1.080 2.280 ;
        RECT  0.920 1.090 1.020 2.280 ;
        RECT  0.120 1.090 0.920 1.250 ;
        RECT  0.580 2.120 0.920 2.280 ;
        RECT  0.300 2.120 0.580 2.400 ;
    END
END OR3X1TR

MACRO OR2XLTR
    CLASS CORE ;
    FOREIGN OR2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.870 1.920 2.760 ;
        RECT  1.600 0.870 1.760 1.090 ;
        RECT  1.660 1.640 1.760 2.760 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.230 1.120 1.560 ;
        RECT  0.900 1.230 1.060 1.710 ;
        RECT  0.880 1.240 0.900 1.710 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.510 0.640 1.770 ;
        RECT  0.080 0.440 0.320 1.770 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.450 -0.280 2.000 0.280 ;
        RECT  1.170 -0.280 1.450 0.500 ;
        RECT  0.000 -0.280 1.170 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.340 3.320 2.000 3.880 ;
        RECT  1.020 2.310 1.340 3.880 ;
        RECT  0.000 3.320 1.020 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.260 1.600 1.480 ;
        RECT  1.280 0.910 1.440 2.150 ;
        RECT  0.890 0.910 1.280 1.070 ;
        RECT  0.440 1.990 1.280 2.150 ;
        RECT  0.610 0.790 0.890 1.070 ;
        RECT  0.160 1.990 0.440 2.270 ;
    END
END OR2XLTR

MACRO OR2X8TR
    CLASS CORE ;
    FOREIGN OR2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 0.820 3.760 2.950 ;
        RECT  3.080 0.820 3.480 2.380 ;
        RECT  2.840 0.820 3.080 1.300 ;
        RECT  2.760 1.900 3.080 2.380 ;
        RECT  2.560 0.440 2.840 1.300 ;
        RECT  2.480 1.900 2.760 3.160 ;
        END
        ANTENNADIFFAREA 7.42 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.590 2.000 2.280 ;
        RECT  0.760 2.120 1.720 2.280 ;
        RECT  0.600 1.590 0.760 2.280 ;
        RECT  0.440 1.590 0.600 1.960 ;
        END
        ANTENNAGATEAREA 0.4704 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.590 1.560 1.960 ;
        RECT  0.920 1.590 1.240 1.870 ;
        END
        ANTENNAGATEAREA 0.4704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.280 -0.280 4.400 0.280 ;
        RECT  3.980 -0.280 4.280 1.030 ;
        RECT  3.320 -0.280 3.980 0.280 ;
        RECT  3.040 -0.280 3.320 0.610 ;
        RECT  2.360 -0.280 3.040 0.280 ;
        RECT  2.080 -0.280 2.360 0.930 ;
        RECT  1.400 -0.280 2.080 0.340 ;
        RECT  1.120 -0.280 1.400 0.930 ;
        RECT  0.440 -0.280 1.120 0.340 ;
        RECT  0.160 -0.280 0.440 1.110 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 3.320 4.400 3.880 ;
        RECT  3.960 1.920 4.240 3.880 ;
        RECT  3.240 3.260 3.960 3.880 ;
        RECT  2.960 2.590 3.240 3.880 ;
        RECT  2.200 3.320 2.960 3.880 ;
        RECT  1.920 2.930 2.200 3.880 ;
        RECT  0.600 3.320 1.920 3.880 ;
        RECT  0.320 2.440 0.600 3.880 ;
        RECT  0.000 3.320 0.320 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.320 1.460 2.900 1.740 ;
        RECT  2.160 1.160 2.320 2.600 ;
        RECT  1.880 1.160 2.160 1.320 ;
        RECT  1.400 2.440 2.160 2.600 ;
        RECT  1.600 1.040 1.880 1.320 ;
        RECT  0.920 1.160 1.600 1.320 ;
        RECT  1.120 2.440 1.400 3.160 ;
        RECT  0.640 1.040 0.920 1.320 ;
    END
END OR2X8TR

MACRO OR2X6TR
    CLASS CORE ;
    FOREIGN OR2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 0.440 3.720 3.160 ;
        RECT  3.400 0.950 3.480 3.160 ;
        RECT  3.080 0.950 3.400 2.280 ;
        RECT  2.800 0.950 3.080 1.310 ;
        RECT  2.720 1.910 3.080 2.280 ;
        RECT  2.520 0.530 2.800 1.310 ;
        RECT  2.440 1.910 2.720 3.160 ;
        END
        ANTENNADIFFAREA 7.48 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.580 1.960 1.860 ;
        RECT  1.680 1.580 1.840 2.280 ;
        RECT  0.720 2.120 1.680 2.280 ;
        RECT  0.440 1.580 0.720 2.280 ;
        END
        ANTENNAGATEAREA 0.372 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.580 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.372 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.280 4.000 0.280 ;
        RECT  3.000 -0.280 3.280 0.670 ;
        RECT  2.320 -0.280 3.000 0.280 ;
        RECT  2.040 -0.280 2.320 1.040 ;
        RECT  1.360 -0.280 2.040 0.340 ;
        RECT  1.080 -0.280 1.360 1.040 ;
        RECT  0.400 -0.280 1.080 0.340 ;
        RECT  0.120 -0.280 0.400 1.040 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.200 3.320 4.000 3.880 ;
        RECT  2.920 2.470 3.200 3.880 ;
        RECT  2.240 3.320 2.920 3.880 ;
        RECT  1.960 2.910 2.240 3.880 ;
        RECT  0.560 3.260 1.960 3.880 ;
        RECT  0.280 2.630 0.560 3.880 ;
        RECT  0.000 3.320 0.280 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 1.470 2.920 1.750 ;
        RECT  2.120 1.200 2.280 2.600 ;
        RECT  1.840 1.200 2.120 1.360 ;
        RECT  1.360 2.440 2.120 2.600 ;
        RECT  1.560 1.030 1.840 1.360 ;
        RECT  0.880 1.200 1.560 1.360 ;
        RECT  1.080 2.440 1.360 2.720 ;
        RECT  0.600 1.030 0.880 1.360 ;
    END
END OR2X6TR

MACRO OR2X4TR
    CLASS CORE ;
    FOREIGN OR2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.440 2.140 2.160 ;
        RECT  1.850 0.440 1.920 3.080 ;
        RECT  1.640 1.920 1.850 3.080 ;
        END
        ANTENNADIFFAREA 3.94 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.160 1.760 ;
        END
        ANTENNAGATEAREA 0.2352 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.370 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2352 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.640 -0.280 2.800 0.280 ;
        RECT  2.360 -0.280 2.640 1.250 ;
        RECT  1.620 -0.280 2.360 0.280 ;
        RECT  1.340 -0.280 1.620 0.760 ;
        RECT  0.560 -0.280 1.340 0.340 ;
        RECT  0.280 -0.280 0.560 0.930 ;
        RECT  0.000 -0.280 0.280 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 3.320 2.800 3.880 ;
        RECT  2.120 2.450 2.400 3.880 ;
        RECT  1.400 3.320 2.120 3.880 ;
        RECT  1.120 2.730 1.400 3.880 ;
        RECT  0.000 3.320 1.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.480 1.660 1.760 ;
        RECT  1.320 0.920 1.480 2.470 ;
        RECT  1.040 0.920 1.320 1.080 ;
        RECT  0.560 2.310 1.320 2.470 ;
        RECT  0.760 0.800 1.040 1.080 ;
        RECT  0.280 2.310 0.560 3.100 ;
    END
END OR2X4TR

MACRO OR2X2TR
    CLASS CORE ;
    FOREIGN OR2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.570 1.920 3.110 ;
        RECT  1.600 0.570 1.760 1.320 ;
        RECT  1.680 1.640 1.760 3.110 ;
        RECT  1.610 2.090 1.680 3.110 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.230 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.240 0.720 1.770 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.080 -0.280 1.360 0.470 ;
        RECT  0.370 -0.280 1.080 0.280 ;
        RECT  0.100 -0.280 0.370 1.040 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 3.320 2.000 3.880 ;
        RECT  1.080 2.470 1.360 3.880 ;
        RECT  0.000 3.320 1.080 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.450 1.580 1.520 1.860 ;
        RECT  1.440 1.580 1.450 2.310 ;
        RECT  1.280 0.910 1.440 2.310 ;
        RECT  0.890 0.910 1.280 1.070 ;
        RECT  0.400 2.150 1.280 2.310 ;
        RECT  0.610 0.790 0.890 1.070 ;
        RECT  0.120 1.990 0.400 2.620 ;
    END
END OR2X2TR

MACRO OR2X1TR
    CLASS CORE ;
    FOREIGN OR2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.760 1.920 2.760 ;
        RECT  1.600 0.760 1.760 1.040 ;
        RECT  1.660 1.640 1.760 2.760 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.230 1.120 1.710 ;
        RECT  0.880 1.240 0.900 1.710 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.550 0.640 1.770 ;
        RECT  0.080 0.440 0.360 1.770 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 3.320 2.000 3.880 ;
        RECT  1.080 2.320 1.360 3.880 ;
        RECT  0.000 3.320 1.080 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.200 1.600 1.480 ;
        RECT  1.280 0.910 1.440 2.150 ;
        RECT  0.890 0.910 1.280 1.070 ;
        RECT  0.440 1.990 1.280 2.150 ;
        RECT  0.610 0.790 0.890 1.070 ;
        RECT  0.160 1.990 0.440 2.270 ;
    END
END OR2X1TR

MACRO OAI33XLTR
    CLASS CORE ;
    FOREIGN OAI33XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.840 3.120 1.960 ;
        RECT  2.880 0.840 3.040 2.680 ;
        RECT  2.870 1.000 2.880 1.280 ;
        RECT  1.640 2.520 2.880 2.680 ;
        RECT  2.110 1.120 2.870 1.280 ;
        RECT  1.950 1.000 2.110 1.280 ;
        RECT  1.380 2.380 1.640 2.680 ;
        END
        ANTENNADIFFAREA 2.548 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.620 1.010 1.780 ;
        RECT  0.480 1.620 0.720 1.980 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.760 1.350 2.100 ;
        RECT  1.120 1.940 1.190 2.100 ;
        RECT  0.880 1.940 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.560 2.720 2.040 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.440 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.640 1.920 2.040 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.280 3.200 0.280 ;
        RECT  0.950 -0.280 1.280 1.190 ;
        RECT  0.370 -0.280 0.950 0.280 ;
        RECT  0.090 -0.280 0.370 0.600 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.850 3.320 3.200 3.880 ;
        RECT  2.570 2.840 2.850 3.880 ;
        RECT  0.430 3.320 2.570 3.880 ;
        RECT  0.270 2.520 0.430 3.880 ;
        RECT  0.000 3.320 0.270 3.880 ;
        END
    END VDD
END OAI33XLTR

MACRO OAI33X4TR
    CLASS CORE ;
    FOREIGN OAI33X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.990 1.920 2.100 ;
        RECT  1.190 0.990 1.640 1.320 ;
        RECT  1.470 1.940 1.640 2.100 ;
        RECT  1.190 1.940 1.470 2.690 ;
        END
        ANTENNADIFFAREA 3.861 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.550 2.200 0.770 ;
        RECT  1.240 0.440 1.560 0.770 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.430 2.590 1.710 ;
        RECT  2.080 1.430 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.580 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.510 4.720 2.760 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.430 3.960 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.700 3.520 2.370 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.790 -0.280 4.800 0.280 ;
        RECT  2.510 -0.280 2.790 0.400 ;
        RECT  2.000 -0.280 2.510 0.280 ;
        RECT  1.720 -0.280 2.000 0.390 ;
        RECT  0.950 -0.280 1.720 0.280 ;
        RECT  0.630 -0.280 0.950 0.910 ;
        RECT  0.000 -0.280 0.630 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.660 3.320 4.800 3.880 ;
        RECT  4.440 2.920 4.660 3.880 ;
        RECT  1.990 3.260 4.440 3.880 ;
        RECT  1.710 3.200 1.990 3.880 ;
        RECT  0.950 3.320 1.710 3.880 ;
        RECT  0.670 3.200 0.950 3.880 ;
        RECT  0.000 3.320 0.670 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.430 0.990 4.710 1.270 ;
        RECT  4.280 1.110 4.430 1.270 ;
        RECT  4.120 1.110 4.280 2.740 ;
        RECT  3.790 1.110 4.120 1.270 ;
        RECT  2.240 2.540 4.120 2.740 ;
        RECT  3.510 0.990 3.790 1.270 ;
        RECT  3.030 0.990 3.310 1.270 ;
        RECT  2.390 1.110 3.030 1.270 ;
        RECT  2.110 0.990 2.390 1.270 ;
        RECT  2.080 2.540 2.240 3.040 ;
        RECT  0.710 2.880 2.080 3.040 ;
        RECT  1.030 1.570 1.480 1.730 ;
        RECT  0.870 1.320 1.030 1.730 ;
        RECT  0.430 1.320 0.870 1.480 ;
        RECT  0.490 1.640 0.710 3.040 ;
        RECT  0.330 0.630 0.430 1.480 ;
        RECT  0.110 0.630 0.330 2.990 ;
    END
END OAI33X4TR

MACRO OAI33X2TR
    CLASS CORE ;
    FOREIGN OAI33X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 0.440 5.920 1.560 ;
        RECT  5.630 2.390 5.890 3.010 ;
        RECT  5.210 0.730 5.680 1.010 ;
        RECT  5.620 2.520 5.630 3.010 ;
        RECT  3.030 2.520 5.620 2.680 ;
        RECT  4.560 0.850 5.210 1.010 ;
        RECT  4.280 0.730 4.560 1.010 ;
        RECT  3.640 0.850 4.280 1.010 ;
        RECT  3.450 0.730 3.640 1.010 ;
        RECT  3.290 0.730 3.450 1.330 ;
        RECT  2.990 1.170 3.290 1.330 ;
        RECT  2.990 2.520 3.030 2.800 ;
        RECT  2.830 1.170 2.990 2.800 ;
        RECT  2.710 2.520 2.830 2.800 ;
        RECT  0.370 2.520 2.710 2.680 ;
        RECT  0.090 2.520 0.370 2.870 ;
        END
        ANTENNADIFFAREA 10.204 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.570 1.660 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.360 2.330 1.640 ;
        RECT  2.050 1.360 2.210 1.980 ;
        RECT  1.120 1.820 2.050 1.980 ;
        RECT  0.880 1.240 1.120 1.980 ;
        RECT  0.730 1.240 0.880 1.640 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.680 2.670 2.360 ;
        RECT  0.510 2.200 2.510 2.360 ;
        RECT  0.320 1.640 0.510 2.360 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.220 4.360 1.660 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.000 1.360 5.250 1.640 ;
        RECT  4.680 1.480 5.000 1.640 ;
        RECT  4.520 1.480 4.680 1.980 ;
        RECT  3.920 1.820 4.520 1.980 ;
        RECT  3.760 1.360 3.920 1.980 ;
        RECT  3.610 1.360 3.760 1.960 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.410 1.760 5.690 2.200 ;
        RECT  5.160 2.040 5.410 2.200 ;
        RECT  4.840 2.040 5.160 2.360 ;
        RECT  3.370 2.200 4.840 2.360 ;
        RECT  3.150 1.700 3.370 2.360 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.280 6.000 0.280 ;
        RECT  2.330 -0.280 2.610 0.400 ;
        RECT  1.690 -0.280 2.330 0.340 ;
        RECT  1.410 -0.280 1.690 0.380 ;
        RECT  0.770 -0.280 1.410 0.280 ;
        RECT  0.490 -0.280 0.770 0.360 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.730 3.320 6.000 3.880 ;
        RECT  4.050 2.850 4.730 3.880 ;
        RECT  1.630 3.320 4.050 3.880 ;
        RECT  1.350 2.850 1.630 3.880 ;
        RECT  0.000 3.320 1.350 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 0.730 3.130 1.010 ;
        RECT  2.210 0.850 2.850 1.010 ;
        RECT  1.930 0.730 2.210 1.010 ;
        RECT  1.290 0.850 1.930 1.010 ;
        RECT  1.010 0.730 1.290 1.010 ;
        RECT  0.370 0.850 1.010 1.010 ;
        RECT  0.090 0.730 0.370 1.010 ;
    END
END OAI33X2TR

MACRO OAI33X1TR
    CLASS CORE ;
    FOREIGN OAI33X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.840 3.520 1.960 ;
        RECT  3.280 0.840 3.440 2.680 ;
        RECT  3.180 1.030 3.280 1.310 ;
        RECT  2.020 2.520 3.280 2.680 ;
        RECT  2.500 1.150 3.180 1.310 ;
        RECT  2.280 1.030 2.500 1.310 ;
        RECT  1.740 2.250 2.020 3.160 ;
        END
        ANTENNADIFFAREA 4.08 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.400 0.720 1.680 ;
        RECT  0.080 1.400 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.470 1.320 1.770 ;
        RECT  0.880 1.470 1.120 1.970 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.810 1.780 2.090 ;
        RECT  1.500 1.810 1.560 2.360 ;
        RECT  1.280 1.930 1.500 2.360 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.640 3.120 2.070 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.470 2.720 2.360 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.100 1.480 2.320 1.960 ;
        RECT  2.040 1.240 2.100 1.960 ;
        RECT  1.940 1.240 2.040 1.900 ;
        RECT  1.680 1.240 1.940 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.540 -0.280 3.600 0.280 ;
        RECT  1.260 -0.280 1.540 0.350 ;
        RECT  0.580 -0.280 1.260 0.280 ;
        RECT  0.300 -0.280 0.580 0.990 ;
        RECT  0.000 -0.280 0.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 3.320 3.600 3.880 ;
        RECT  2.860 2.870 3.140 3.880 ;
        RECT  0.860 3.320 2.860 3.880 ;
        RECT  0.580 2.350 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.710 2.980 0.990 ;
        RECT  2.020 0.710 2.660 0.870 ;
        RECT  1.900 0.710 2.020 0.990 ;
        RECT  1.740 0.710 1.900 1.080 ;
        RECT  1.080 0.920 1.740 1.080 ;
        RECT  0.780 0.920 1.080 1.240 ;
    END
END OAI33X1TR

MACRO OAI32XLTR
    CLASS CORE ;
    FOREIGN OAI32XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.840 2.720 2.600 ;
        RECT  1.970 1.090 2.480 1.250 ;
        RECT  1.650 2.440 2.480 2.600 ;
        RECT  1.370 2.200 1.650 2.600 ;
        END
        ANTENNADIFFAREA 1.2335 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.840 2.040 3.160 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.640 2.320 1.960 ;
        RECT  1.640 1.420 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.420 1.040 1.580 ;
        RECT  0.480 1.420 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.760 1.480 1.920 ;
        RECT  0.880 1.760 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.280 2.800 0.280 ;
        RECT  0.970 -0.280 1.250 0.580 ;
        RECT  0.390 -0.280 0.970 0.280 ;
        RECT  0.090 -0.280 0.390 1.240 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.500 3.320 2.800 3.880 ;
        RECT  2.220 2.800 2.500 3.880 ;
        RECT  0.460 3.320 2.220 3.880 ;
        RECT  0.180 2.920 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.570 1.020 1.770 1.180 ;
    END
END OAI32XLTR

MACRO OAI32X4TR
    CLASS CORE ;
    FOREIGN OAI32X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.180 0.440 4.320 1.370 ;
        RECT  3.940 0.440 4.180 3.160 ;
        RECT  3.900 0.440 3.940 1.310 ;
        RECT  3.900 1.910 3.940 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.720 2.720 2.360 ;
        RECT  2.040 1.720 2.440 2.000 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 2.440 1.960 2.800 ;
        RECT  1.640 2.440 1.920 2.920 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.600 0.620 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.240 1.120 1.660 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.520 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.280 4.800 0.280 ;
        RECT  4.480 -0.280 4.700 1.310 ;
        RECT  3.660 -0.280 4.480 0.280 ;
        RECT  3.380 -0.280 3.660 0.770 ;
        RECT  1.300 -0.280 3.380 0.340 ;
        RECT  1.020 -0.280 1.300 0.400 ;
        RECT  0.380 -0.280 1.020 0.340 ;
        RECT  0.100 -0.280 0.380 1.080 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.420 1.910 4.700 3.880 ;
        RECT  3.660 3.320 4.420 3.880 ;
        RECT  3.380 2.040 3.660 3.880 ;
        RECT  2.560 3.260 3.380 3.880 ;
        RECT  2.280 2.800 2.560 3.880 ;
        RECT  0.380 3.260 2.280 3.880 ;
        RECT  0.100 2.520 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.660 1.470 3.780 1.750 ;
        RECT  3.500 0.930 3.660 1.880 ;
        RECT  3.180 0.930 3.500 1.090 ;
        RECT  3.140 1.720 3.500 1.880 ;
        RECT  3.060 1.280 3.340 1.560 ;
        RECT  3.020 0.500 3.180 1.090 ;
        RECT  2.980 1.720 3.140 2.770 ;
        RECT  2.320 1.400 3.060 1.560 ;
        RECT  2.900 0.500 3.020 0.780 ;
        RECT  2.920 1.910 2.980 2.770 ;
        RECT  2.640 0.960 2.800 1.240 ;
        RECT  2.480 0.710 2.640 1.240 ;
        RECT  1.840 0.710 2.480 0.870 ;
        RECT  2.040 1.030 2.320 1.560 ;
        RECT  1.880 1.400 2.040 1.560 ;
        RECT  1.720 1.400 1.880 2.280 ;
        RECT  1.680 0.710 1.840 1.210 ;
        RECT  1.480 2.120 1.720 2.280 ;
        RECT  1.560 0.800 1.680 1.210 ;
        RECT  0.620 0.800 1.560 1.080 ;
        RECT  1.260 2.120 1.480 2.400 ;
    END
END OAI32X4TR

MACRO OAI32X2TR
    CLASS CORE ;
    FOREIGN OAI32X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.000 0.840 5.120 1.960 ;
        RECT  4.880 0.840 5.000 2.320 ;
        RECT  4.840 1.030 4.880 2.320 ;
        RECT  4.330 1.030 4.840 1.330 ;
        RECT  4.690 2.160 4.840 2.320 ;
        RECT  4.410 2.160 4.690 2.900 ;
        RECT  3.010 2.520 4.410 2.680 ;
        RECT  3.650 1.170 4.330 1.330 ;
        RECT  3.490 1.030 3.650 1.330 ;
        RECT  3.370 1.030 3.490 1.310 ;
        RECT  2.730 2.160 3.010 3.100 ;
        RECT  2.690 2.500 2.730 3.100 ;
        RECT  0.650 2.500 2.690 2.660 ;
        RECT  0.370 2.240 0.650 3.100 ;
        END
        ANTENNADIFFAREA 7.4 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.770 1.810 4.050 2.360 ;
        RECT  3.680 2.040 3.770 2.360 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.370 1.720 4.490 2.000 ;
        RECT  4.210 1.490 4.370 2.000 ;
        RECT  3.520 1.490 4.210 1.650 ;
        RECT  3.090 1.490 3.520 1.960 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.640 1.980 1.990 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.240 2.430 1.400 ;
        RECT  0.880 1.240 1.120 1.620 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 1.720 2.770 2.000 ;
        RECT  2.410 1.720 2.570 2.310 ;
        RECT  0.970 2.150 2.410 2.310 ;
        RECT  0.810 1.780 0.970 2.310 ;
        RECT  0.720 1.780 0.810 1.960 ;
        RECT  0.370 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.770 -0.280 5.200 0.280 ;
        RECT  2.490 -0.280 2.770 0.400 ;
        RECT  1.770 -0.280 2.490 0.280 ;
        RECT  1.490 -0.280 1.770 0.670 ;
        RECT  0.000 -0.280 1.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.850 3.320 5.200 3.880 ;
        RECT  3.570 2.840 3.850 3.880 ;
        RECT  1.770 3.320 3.570 3.880 ;
        RECT  1.490 2.820 1.770 3.880 ;
        RECT  0.000 3.320 1.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.010 0.730 4.130 1.010 ;
        RECT  3.850 0.710 4.010 1.010 ;
        RECT  3.170 0.710 3.850 0.870 ;
        RECT  3.010 0.710 3.170 1.010 ;
        RECT  2.890 0.730 3.010 1.010 ;
        RECT  2.250 0.850 2.890 1.010 ;
        RECT  1.970 0.720 2.250 1.010 ;
        RECT  1.290 0.850 1.970 1.010 ;
        RECT  1.010 0.720 1.290 1.010 ;
        RECT  0.370 0.850 1.010 1.010 ;
        RECT  0.090 0.730 0.370 1.010 ;
    END
END OAI32X2TR

MACRO OAI32X1TR
    CLASS CORE ;
    FOREIGN OAI32X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.870 2.320 1.560 ;
        RECT  2.080 0.870 2.240 2.280 ;
        RECT  2.010 0.870 2.080 1.150 ;
        RECT  1.460 2.120 2.080 2.280 ;
        RECT  1.300 2.120 1.460 2.890 ;
        END
        ANTENNADIFFAREA 3.174 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 1.380 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.360 1.000 1.580 ;
        RECT  0.480 1.360 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.620 1.410 1.900 ;
        RECT  1.120 1.740 1.250 1.900 ;
        RECT  0.880 1.740 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 3.320 2.800 3.880 ;
        RECT  2.150 2.660 2.430 3.880 ;
        RECT  0.430 3.320 2.150 3.880 ;
        RECT  0.120 2.240 0.430 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.550 2.650 0.990 ;
        RECT  1.690 0.550 2.490 0.710 ;
        RECT  1.530 0.550 1.690 0.990 ;
        RECT  0.770 0.830 1.530 0.990 ;
        RECT  0.610 0.710 0.770 0.990 ;
    END
END OAI32X1TR

MACRO OAI31XLTR
    CLASS CORE ;
    FOREIGN OAI31XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.440 2.320 2.280 ;
        RECT  1.900 0.850 2.080 1.010 ;
        RECT  1.580 2.120 2.080 2.280 ;
        RECT  1.290 2.120 1.580 2.530 ;
        END
        ANTENNADIFFAREA 1.664 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.800 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.720 0.440 2.000 ;
        RECT  0.080 0.440 0.320 2.000 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.360 0.920 1.640 ;
        RECT  0.670 1.240 0.720 1.640 ;
        RECT  0.480 1.240 0.670 1.560 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.410 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 3.320 2.400 3.880 ;
        RECT  1.780 2.440 2.060 3.880 ;
        RECT  0.460 3.320 1.780 3.880 ;
        RECT  0.190 2.340 0.460 3.880 ;
        RECT  0.000 3.320 0.190 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 0.710 1.640 0.990 ;
        RECT  0.720 0.830 1.480 0.990 ;
        RECT  0.560 0.710 0.720 0.990 ;
    END
END OAI31XLTR

MACRO OAI31X4TR
    CLASS CORE ;
    FOREIGN OAI31X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.030 4.060 1.950 ;
        RECT  3.840 1.030 3.920 3.160 ;
        RECT  3.820 0.470 3.840 3.160 ;
        RECT  3.530 0.470 3.820 1.310 ;
        RECT  3.600 1.790 3.820 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.140 2.040 1.560 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.620 0.640 1.780 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.240 1.120 1.630 ;
        RECT  0.800 1.230 1.060 1.630 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.280 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.280 4.400 0.280 ;
        RECT  4.020 -0.280 4.290 0.750 ;
        RECT  3.330 -0.280 4.020 0.280 ;
        RECT  3.040 -0.280 3.330 0.950 ;
        RECT  1.260 -0.280 3.040 0.280 ;
        RECT  1.100 -0.280 1.260 0.400 ;
        RECT  0.460 -0.280 1.100 0.280 ;
        RECT  0.150 -0.280 0.460 1.080 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 3.320 4.400 3.880 ;
        RECT  4.080 2.110 4.240 3.880 ;
        RECT  3.350 3.320 4.080 3.880 ;
        RECT  3.060 2.360 3.350 3.880 ;
        RECT  2.250 3.320 3.060 3.880 ;
        RECT  2.000 2.090 2.250 3.880 ;
        RECT  0.550 3.320 2.000 3.880 ;
        RECT  0.230 2.680 0.550 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.340 1.470 3.660 1.630 ;
        RECT  3.180 1.150 3.340 2.200 ;
        RECT  2.790 1.150 3.180 1.310 ;
        RECT  2.840 2.040 3.180 2.200 ;
        RECT  2.370 1.640 3.020 1.880 ;
        RECT  2.540 2.040 2.840 2.740 ;
        RECT  2.630 0.790 2.790 1.310 ;
        RECT  2.210 0.760 2.370 1.880 ;
        RECT  2.040 0.760 2.210 0.920 ;
        RECT  1.840 1.720 2.210 1.880 ;
        RECT  1.680 1.720 1.840 2.360 ;
        RECT  1.620 0.660 1.780 0.980 ;
        RECT  1.410 2.200 1.680 2.360 ;
        RECT  0.920 0.820 1.620 0.980 ;
        RECT  0.760 0.820 0.920 1.070 ;
        RECT  0.640 0.910 0.760 1.070 ;
    END
END OAI31X4TR

MACRO OAI31X2TR
    CLASS CORE ;
    FOREIGN OAI31X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.640 3.920 2.230 ;
        RECT  3.680 0.800 3.840 2.230 ;
        RECT  3.440 0.800 3.680 1.080 ;
        RECT  3.480 2.070 3.680 2.230 ;
        RECT  3.320 2.070 3.480 2.600 ;
        RECT  3.200 2.320 3.320 2.600 ;
        RECT  1.800 2.440 3.200 2.600 ;
        RECT  1.520 2.440 1.800 3.070 ;
        END
        ANTENNADIFFAREA 4.122 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.240 3.520 1.910 ;
        END
        ANTENNAGATEAREA 0.3 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.640 3.120 1.960 ;
        RECT  2.760 1.680 2.840 1.960 ;
        RECT  2.600 1.680 2.760 2.280 ;
        RECT  1.000 2.120 2.600 2.280 ;
        RECT  0.840 1.800 1.000 2.280 ;
        RECT  0.680 1.800 0.840 1.960 ;
        RECT  0.400 1.680 0.680 1.960 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.360 2.440 1.640 ;
        RECT  2.160 1.240 2.320 1.640 ;
        RECT  1.200 1.240 2.160 1.400 ;
        RECT  0.840 1.240 1.200 1.640 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.680 2.000 1.960 ;
        RECT  1.640 1.640 1.960 1.960 ;
        RECT  1.360 1.680 1.640 1.960 ;
        END
        ANTENNAGATEAREA 0.396 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 -0.280 4.400 0.280 ;
        RECT  2.480 -0.280 2.760 0.390 ;
        RECT  1.840 -0.280 2.480 0.340 ;
        RECT  1.560 -0.280 1.840 0.390 ;
        RECT  0.920 -0.280 1.560 0.340 ;
        RECT  0.640 -0.280 0.920 0.390 ;
        RECT  0.000 -0.280 0.640 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.960 3.320 4.400 3.880 ;
        RECT  3.680 2.390 3.960 3.880 ;
        RECT  2.960 3.320 3.680 3.880 ;
        RECT  2.680 2.760 2.960 3.880 ;
        RECT  0.680 3.320 2.680 3.880 ;
        RECT  0.400 2.120 0.680 3.880 ;
        RECT  0.000 3.320 0.400 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.160 0.700 4.280 0.980 ;
        RECT  4.000 0.480 4.160 0.980 ;
        RECT  3.160 0.480 4.000 0.640 ;
        RECT  3.000 0.480 3.160 0.980 ;
        RECT  2.880 0.700 3.000 0.980 ;
        RECT  2.240 0.820 2.880 0.980 ;
        RECT  1.960 0.700 2.240 0.980 ;
        RECT  1.320 0.820 1.960 0.980 ;
        RECT  1.040 0.700 1.320 0.980 ;
        RECT  0.400 0.820 1.040 0.980 ;
        RECT  0.120 0.820 0.400 1.100 ;
    END
END OAI31X2TR

MACRO OAI31X1TR
    CLASS CORE ;
    FOREIGN OAI31X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.440 2.320 2.280 ;
        RECT  1.900 0.920 2.080 1.080 ;
        RECT  1.580 2.120 2.080 2.280 ;
        RECT  1.290 2.120 1.580 2.530 ;
        END
        ANTENNADIFFAREA 2.587 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.800 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.720 0.440 2.000 ;
        RECT  0.080 0.440 0.320 2.000 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.360 0.920 1.640 ;
        RECT  0.670 1.240 0.720 1.640 ;
        RECT  0.480 1.240 0.670 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.410 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 3.320 2.400 3.880 ;
        RECT  1.780 2.440 2.060 3.880 ;
        RECT  0.460 3.320 1.780 3.880 ;
        RECT  0.190 2.340 0.460 3.880 ;
        RECT  0.000 3.320 0.190 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 0.710 1.640 0.990 ;
        RECT  0.720 0.830 1.480 0.990 ;
        RECT  0.560 0.710 0.720 0.990 ;
    END
END OAI31X1TR

MACRO OAI2BB2XLTR
    CLASS CORE ;
    FOREIGN OAI2BB2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.900 2.720 2.800 ;
        RECT  2.410 0.900 2.480 1.140 ;
        RECT  1.910 2.520 2.480 2.800 ;
        END
        ANTENNADIFFAREA 1.0995 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.520 1.200 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.030 2.070 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.700 1.540 3.160 ;
        RECT  0.760 2.700 1.220 2.880 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.370 0.410 1.650 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.280 2.800 0.280 ;
        RECT  1.460 -0.280 2.140 0.340 ;
        RECT  0.410 -0.280 1.460 0.280 ;
        RECT  0.130 -0.280 0.410 0.460 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.420 3.320 2.800 3.880 ;
        RECT  2.140 3.200 2.420 3.880 ;
        RECT  0.410 3.320 2.140 3.880 ;
        RECT  0.130 2.800 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.040 1.580 2.260 1.870 ;
        RECT  1.970 0.660 2.190 1.250 ;
        RECT  1.520 1.580 2.040 1.740 ;
        RECT  1.220 0.660 1.970 0.820 ;
        RECT  1.360 1.170 1.520 2.400 ;
        RECT  1.170 1.170 1.360 1.330 ;
        RECT  0.860 2.240 1.360 2.400 ;
        RECT  0.930 0.540 1.220 0.820 ;
        RECT  0.890 1.010 1.170 1.330 ;
        RECT  0.580 2.210 0.860 2.490 ;
    END
END OAI2BB2XLTR

MACRO OAI2BB2X4TR
    CLASS CORE ;
    FOREIGN OAI2BB2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.000 0.960 6.240 3.160 ;
        RECT  5.000 0.960 6.000 1.200 ;
        RECT  5.920 1.840 6.000 3.160 ;
        RECT  5.680 1.840 5.920 2.830 ;
        RECT  4.880 2.590 5.680 2.830 ;
        RECT  4.760 0.960 5.000 1.520 ;
        RECT  4.600 2.590 4.880 2.890 ;
        RECT  4.160 1.280 4.760 1.520 ;
        RECT  3.840 2.590 4.600 2.830 ;
        RECT  4.000 1.090 4.160 1.520 ;
        RECT  3.840 1.090 4.000 1.370 ;
        RECT  3.560 2.590 3.840 2.890 ;
        RECT  2.520 2.590 3.560 2.830 ;
        RECT  2.240 2.590 2.520 3.160 ;
        END
        ANTENNADIFFAREA 8.312 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.760 1.680 4.880 1.840 ;
        RECT  4.600 1.680 4.760 2.110 ;
        RECT  3.120 1.950 4.600 2.110 ;
        RECT  3.000 1.720 3.120 2.110 ;
        RECT  2.840 1.460 3.000 2.110 ;
        RECT  1.920 1.460 2.840 1.620 ;
        RECT  1.680 1.460 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.460 1.360 5.640 1.520 ;
        RECT  5.300 1.360 5.460 2.430 ;
        RECT  2.680 2.270 5.300 2.430 ;
        RECT  2.520 1.800 2.680 2.430 ;
        RECT  2.320 1.800 2.520 1.960 ;
        RECT  2.080 1.800 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.640 1.520 2.360 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.680 1.920 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.160 -0.280 6.400 0.280 ;
        RECT  5.880 -0.280 6.160 0.800 ;
        RECT  5.120 -0.280 5.880 0.280 ;
        RECT  4.840 -0.280 5.120 0.400 ;
        RECT  3.120 -0.280 4.840 0.280 ;
        RECT  2.840 -0.280 3.120 0.400 ;
        RECT  1.720 -0.280 2.840 0.340 ;
        RECT  1.440 -0.280 1.720 0.670 ;
        RECT  0.580 -0.280 1.440 0.280 ;
        RECT  0.300 -0.280 0.580 1.080 ;
        RECT  0.000 -0.280 0.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.400 3.320 6.400 3.880 ;
        RECT  5.120 2.990 5.400 3.880 ;
        RECT  4.360 3.260 5.120 3.880 ;
        RECT  4.080 3.200 4.360 3.880 ;
        RECT  3.320 3.260 4.080 3.880 ;
        RECT  3.040 2.990 3.320 3.880 ;
        RECT  1.680 3.320 3.040 3.880 ;
        RECT  1.400 2.800 1.680 3.880 ;
        RECT  0.580 3.320 1.400 3.880 ;
        RECT  0.300 2.530 0.580 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.360 0.460 5.640 0.740 ;
        RECT  4.600 0.580 5.360 0.740 ;
        RECT  4.320 0.440 4.600 1.120 ;
        RECT  3.640 0.590 4.320 0.750 ;
        RECT  3.680 1.630 3.840 1.790 ;
        RECT  3.520 1.120 3.680 1.790 ;
        RECT  3.360 0.590 3.640 0.870 ;
        RECT  1.380 1.120 3.520 1.280 ;
        RECT  2.200 0.710 3.360 0.870 ;
        RECT  1.920 0.590 2.200 0.870 ;
        RECT  1.100 0.990 1.380 1.280 ;
        RECT  1.000 1.120 1.100 1.280 ;
        RECT  0.840 1.120 1.000 3.160 ;
    END
END OAI2BB2X4TR

MACRO OAI2BB2X2TR
    CLASS CORE ;
    FOREIGN OAI2BB2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.240 4.320 2.360 ;
        RECT  4.080 1.240 4.240 2.680 ;
        RECT  3.890 1.240 4.080 1.400 ;
        RECT  3.510 2.520 4.080 2.680 ;
        RECT  3.730 1.070 3.890 1.400 ;
        RECT  2.610 1.070 3.730 1.230 ;
        RECT  3.230 2.400 3.510 3.100 ;
        RECT  2.260 2.400 3.230 2.560 ;
        RECT  2.100 2.400 2.260 3.140 ;
        RECT  1.950 2.920 2.100 3.140 ;
        END
        ANTENNADIFFAREA 4.759 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 1.390 3.570 1.920 ;
        RECT  1.710 1.760 3.410 1.920 ;
        RECT  1.520 1.600 1.710 1.920 ;
        RECT  1.360 1.600 1.520 2.360 ;
        RECT  1.280 2.040 1.360 2.360 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 2.080 3.840 2.360 ;
        RECT  1.920 2.080 3.680 2.240 ;
        RECT  1.750 2.080 1.920 2.760 ;
        RECT  1.680 2.440 1.750 2.760 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.480 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.570 0.400 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.280 4.400 0.280 ;
        RECT  3.590 -0.280 3.870 0.400 ;
        RECT  1.950 -0.280 3.590 0.280 ;
        RECT  0.370 -0.280 1.950 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 3.320 4.400 3.880 ;
        RECT  2.750 2.910 3.030 3.880 ;
        RECT  1.430 3.320 2.750 3.880 ;
        RECT  1.150 2.890 1.430 3.880 ;
        RECT  0.370 3.260 1.150 3.880 ;
        RECT  0.090 2.780 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.050 0.650 4.270 1.080 ;
        RECT  3.310 0.650 4.050 0.810 ;
        RECT  3.030 0.480 3.310 0.810 ;
        RECT  2.030 1.420 3.190 1.580 ;
        RECT  2.350 0.650 3.030 0.810 ;
        RECT  2.070 0.650 2.350 0.930 ;
        RECT  1.430 0.650 2.070 0.810 ;
        RECT  1.870 1.160 2.030 1.580 ;
        RECT  1.090 1.160 1.870 1.320 ;
        RECT  1.150 0.530 1.430 0.810 ;
        RECT  0.810 1.030 1.090 1.320 ;
        RECT  0.720 2.120 0.890 2.400 ;
        RECT  0.720 1.160 0.810 1.320 ;
        RECT  0.560 1.160 0.720 2.400 ;
    END
END OAI2BB2X2TR

MACRO OAI2BB2X1TR
    CLASS CORE ;
    FOREIGN OAI2BB2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.030 3.120 2.360 ;
        RECT  2.500 2.120 2.840 2.360 ;
        RECT  2.220 2.120 2.500 2.400 ;
        END
        ANTENNADIFFAREA 2.312 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.840 1.560 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.200 2.360 1.640 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.480 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.680 0.400 1.980 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 -0.280 3.200 0.280 ;
        RECT  2.400 -0.280 2.680 0.340 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  1.940 -0.280 2.220 0.400 ;
        RECT  1.000 -0.280 1.940 0.280 ;
        RECT  0.720 -0.280 1.000 0.340 ;
        RECT  0.400 -0.280 0.720 0.280 ;
        RECT  0.120 -0.280 0.400 0.400 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.020 3.320 3.200 3.880 ;
        RECT  2.740 2.800 3.020 3.880 ;
        RECT  1.660 3.260 2.740 3.880 ;
        RECT  1.380 2.440 1.660 3.880 ;
        RECT  0.400 3.260 1.380 3.880 ;
        RECT  0.120 2.800 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.520 1.580 2.680 1.960 ;
        RECT  2.340 0.710 2.620 0.990 ;
        RECT  1.800 1.800 2.520 1.960 ;
        RECT  1.700 0.830 2.340 0.990 ;
        RECT  1.640 1.800 1.800 2.280 ;
        RECT  1.420 0.710 1.700 0.990 ;
        RECT  1.040 2.120 1.640 2.280 ;
        RECT  0.960 0.790 1.240 1.070 ;
        RECT  0.720 2.120 1.040 2.400 ;
        RECT  0.720 0.910 0.960 1.070 ;
        RECT  0.560 0.910 0.720 2.400 ;
    END
END OAI2BB2X1TR

MACRO OAI2BB1XLTR
    CLASS CORE ;
    FOREIGN OAI2BB1XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.840 2.320 2.910 ;
        RECT  2.080 0.840 2.160 1.960 ;
        RECT  1.760 2.750 2.160 2.910 ;
        RECT  2.040 0.840 2.080 1.180 ;
        RECT  1.920 0.900 2.040 1.180 ;
        RECT  1.480 2.750 1.760 3.030 ;
        END
        ANTENNADIFFAREA 1.952 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.840 1.560 1.650 ;
        RECT  1.240 0.840 1.280 1.160 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.440 0.760 0.870 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.640 1.120 1.970 ;
        RECT  0.800 1.570 1.060 1.970 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.280 2.400 0.280 ;
        RECT  1.040 -0.280 1.320 0.400 ;
        RECT  0.000 -0.280 1.040 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.320 2.400 3.880 ;
        RECT  1.940 3.200 2.220 3.880 ;
        RECT  1.300 3.320 1.940 3.880 ;
        RECT  1.020 2.800 1.300 3.880 ;
        RECT  0.380 3.260 1.020 3.880 ;
        RECT  0.090 2.500 0.380 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 1.690 1.920 2.290 ;
        RECT  0.840 2.130 1.720 2.290 ;
        RECT  0.560 2.130 0.840 2.890 ;
        RECT  0.450 2.130 0.560 2.290 ;
        RECT  0.290 1.030 0.450 2.290 ;
        RECT  0.170 1.030 0.290 1.310 ;
    END
END OAI2BB1XLTR

MACRO OAI2BB1X4TR
    CLASS CORE ;
    FOREIGN OAI2BB1X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 0.500 3.910 1.210 ;
        RECT  3.590 0.500 3.750 2.350 ;
        RECT  2.300 0.770 3.590 0.930 ;
        RECT  3.200 2.110 3.590 2.350 ;
        RECT  2.880 2.110 3.200 3.160 ;
        RECT  2.310 2.110 2.880 2.360 ;
        RECT  2.020 2.110 2.310 3.160 ;
        RECT  2.080 0.650 2.300 0.930 ;
        END
        ANTENNADIFFAREA 7.396 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.090 2.980 1.540 ;
        RECT  1.920 1.090 2.700 1.250 ;
        RECT  1.680 0.840 1.920 1.250 ;
        RECT  1.640 1.090 1.680 1.250 ;
        RECT  1.480 1.090 1.640 1.630 ;
        END
        ANTENNAGATEAREA 0.6024 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.570 0.400 1.860 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.228 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.200 1.300 1.630 ;
        END
        ANTENNAGATEAREA 0.228 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.100 -0.280 4.000 0.280 ;
        RECT  2.820 -0.280 3.100 0.610 ;
        RECT  1.500 -0.280 2.820 0.280 ;
        RECT  1.220 -0.280 1.500 0.900 ;
        RECT  0.400 -0.280 1.220 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.740 3.320 4.000 3.880 ;
        RECT  3.460 2.910 3.740 3.880 ;
        RECT  2.720 3.320 3.460 3.880 ;
        RECT  2.560 2.910 2.720 3.880 ;
        RECT  1.650 3.320 2.560 3.880 ;
        RECT  1.370 2.140 1.650 3.880 ;
        RECT  0.490 3.320 1.370 3.880 ;
        RECT  0.210 2.680 0.490 3.880 ;
        RECT  0.000 3.320 0.210 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 1.580 3.430 1.880 ;
        RECT  2.140 1.720 3.150 1.880 ;
        RECT  1.960 1.410 2.140 1.880 ;
        RECT  1.800 1.410 1.960 1.950 ;
        RECT  1.020 1.790 1.800 1.950 ;
        RECT  0.740 1.790 1.020 2.970 ;
        RECT  0.720 1.790 0.740 1.950 ;
        RECT  0.700 0.900 0.720 1.950 ;
        RECT  0.560 0.750 0.700 1.950 ;
        RECT  0.420 0.750 0.560 1.060 ;
    END
END OAI2BB1X4TR

MACRO OAI2BB1X2TR
    CLASS CORE ;
    FOREIGN OAI2BB1X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.960 0.840 3.120 2.200 ;
        RECT  2.260 0.840 2.960 1.000 ;
        RECT  2.360 2.040 2.960 2.200 ;
        RECT  2.320 2.040 2.360 2.360 ;
        RECT  2.040 2.040 2.320 3.160 ;
        RECT  1.980 0.720 2.260 1.000 ;
        END
        ANTENNADIFFAREA 3.75 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.660 1.240 2.800 1.860 ;
        RECT  2.580 1.160 2.660 1.860 ;
        RECT  2.440 1.160 2.580 1.560 ;
        RECT  1.380 1.160 2.440 1.440 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.720 1.770 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.600 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.100 -0.280 3.200 0.280 ;
        RECT  2.820 -0.280 3.100 0.680 ;
        RECT  1.450 -0.280 2.820 0.280 ;
        RECT  1.200 -0.280 1.450 1.000 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 3.320 3.200 3.880 ;
        RECT  2.560 2.360 2.840 3.880 ;
        RECT  1.740 3.320 2.560 3.880 ;
        RECT  1.460 2.460 1.740 3.880 ;
        RECT  0.650 3.260 1.460 3.880 ;
        RECT  0.370 1.950 0.650 3.880 ;
        RECT  0.000 3.320 0.370 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.880 1.600 2.060 1.880 ;
        RECT  1.720 1.600 1.880 2.280 ;
        RECT  1.170 2.120 1.720 2.280 ;
        RECT  1.040 2.120 1.170 2.400 ;
        RECT  0.880 0.920 1.040 2.400 ;
        RECT  0.650 0.920 0.880 1.080 ;
        RECT  0.370 0.800 0.650 1.080 ;
    END
END OAI2BB1X2TR

MACRO OAI2BB1X1TR
    CLASS CORE ;
    FOREIGN OAI2BB1X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.880 2.320 2.700 ;
        RECT  1.920 0.880 2.080 1.160 ;
        RECT  1.760 2.540 2.080 2.700 ;
        RECT  1.600 2.540 1.760 3.140 ;
        RECT  1.480 2.980 1.600 3.140 ;
        END
        ANTENNADIFFAREA 2.624 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.840 1.560 1.580 ;
        RECT  1.240 0.840 1.280 1.160 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.440 0.790 0.810 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.640 1.120 1.960 ;
        RECT  0.820 1.640 1.060 2.060 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.280 2.400 0.280 ;
        RECT  1.080 -0.280 1.360 0.400 ;
        RECT  0.000 -0.280 1.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.320 2.400 3.880 ;
        RECT  1.940 3.200 2.220 3.880 ;
        RECT  1.300 3.320 1.940 3.880 ;
        RECT  1.020 2.800 1.300 3.880 ;
        RECT  0.500 3.260 1.020 3.880 ;
        RECT  0.220 3.200 0.500 3.880 ;
        RECT  0.000 3.320 0.220 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 1.640 1.900 2.380 ;
        RECT  0.840 2.220 1.740 2.380 ;
        RECT  0.560 2.220 0.840 2.860 ;
        RECT  0.520 2.220 0.560 2.380 ;
        RECT  0.360 0.970 0.520 2.380 ;
        RECT  0.240 0.970 0.360 1.250 ;
    END
END OAI2BB1X1TR

MACRO OAI22XLTR
    CLASS CORE ;
    FOREIGN OAI22XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.150 2.320 2.680 ;
        RECT  1.830 1.150 2.080 1.310 ;
        RECT  1.350 2.520 2.080 2.680 ;
        RECT  1.550 0.910 1.830 1.310 ;
        RECT  1.070 2.120 1.350 2.680 ;
        END
        ANTENNADIFFAREA 0.72 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.560 0.540 1.880 ;
        RECT  0.320 1.240 0.330 1.880 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.360 1.020 1.640 ;
        RECT  0.700 1.360 0.860 2.360 ;
        RECT  0.480 2.040 0.700 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.480 1.920 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.540 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 -0.280 2.400 0.280 ;
        RECT  0.550 -0.280 0.830 0.400 ;
        RECT  0.000 -0.280 0.550 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.230 3.320 2.400 3.880 ;
        RECT  1.950 2.840 2.230 3.880 ;
        RECT  0.510 3.260 1.950 3.880 ;
        RECT  0.230 2.800 0.510 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.040 0.590 2.310 0.990 ;
        RECT  1.350 0.590 2.040 0.750 ;
        RECT  1.190 0.590 1.350 1.060 ;
        RECT  0.150 0.840 1.190 1.060 ;
    END
END OAI22XLTR

MACRO OAI22X4TR
    CLASS CORE ;
    FOREIGN OAI22X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 0.980 5.920 2.400 ;
        RECT  3.560 0.980 5.680 1.260 ;
        RECT  5.600 2.150 5.680 2.400 ;
        RECT  5.320 2.150 5.600 3.100 ;
        RECT  4.000 2.440 5.320 2.680 ;
        RECT  3.720 2.440 4.000 3.070 ;
        RECT  2.400 2.520 3.720 2.760 ;
        RECT  2.120 2.240 2.400 3.070 ;
        RECT  0.800 2.240 2.120 2.510 ;
        RECT  0.520 2.240 0.800 3.100 ;
        END
        ANTENNADIFFAREA 12.099 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 1.420 3.120 1.960 ;
        RECT  1.740 1.420 2.800 1.580 ;
        RECT  1.180 1.420 1.740 1.760 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.740 2.600 2.020 ;
        RECT  1.980 1.740 2.140 2.080 ;
        RECT  0.760 1.920 1.980 2.080 ;
        RECT  0.440 1.640 0.760 2.080 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.670 1.740 4.960 2.280 ;
        RECT  3.520 2.120 4.670 2.280 ;
        RECT  3.280 1.420 3.520 2.360 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.710 5.400 1.990 ;
        RECT  5.120 1.420 5.280 1.990 ;
        RECT  4.360 1.420 5.120 1.580 ;
        RECT  3.920 1.420 4.360 1.960 ;
        END
        ANTENNAGATEAREA 0.696 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.880 -0.280 6.400 0.280 ;
        RECT  2.600 -0.280 2.880 0.930 ;
        RECT  1.920 -0.280 2.600 0.340 ;
        RECT  1.640 -0.280 1.920 0.930 ;
        RECT  0.960 -0.280 1.640 0.280 ;
        RECT  0.680 -0.280 0.960 0.930 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.800 3.320 6.400 3.880 ;
        RECT  4.520 2.930 4.800 3.880 ;
        RECT  3.200 3.320 4.520 3.880 ;
        RECT  2.920 2.930 3.200 3.880 ;
        RECT  1.600 3.320 2.920 3.880 ;
        RECT  1.320 2.830 1.600 3.880 ;
        RECT  0.000 3.320 1.320 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.360 0.540 6.240 0.820 ;
        RECT  3.080 0.490 3.360 1.260 ;
        RECT  2.400 1.100 3.080 1.260 ;
        RECT  2.120 0.590 2.400 1.260 ;
        RECT  1.440 1.100 2.120 1.260 ;
        RECT  1.160 0.620 1.440 1.260 ;
        RECT  0.480 1.100 1.160 1.260 ;
        RECT  0.200 0.860 0.480 1.260 ;
    END
END OAI22X4TR

MACRO OAI22X2TR
    CLASS CORE ;
    FOREIGN OAI22X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.140 4.320 2.600 ;
        RECT  3.720 1.140 4.080 1.300 ;
        RECT  3.080 2.440 4.080 2.600 ;
        RECT  3.440 1.020 3.720 1.300 ;
        RECT  2.800 1.140 3.440 1.300 ;
        RECT  2.800 2.440 3.080 2.720 ;
        RECT  2.480 1.020 2.800 1.300 ;
        RECT  1.360 2.440 2.800 2.600 ;
        RECT  1.080 2.440 1.360 2.720 ;
        END
        ANTENNADIFFAREA 5.28 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.580 2.000 1.860 ;
        RECT  1.720 1.580 1.880 2.280 ;
        RECT  0.720 2.120 1.720 2.280 ;
        RECT  0.560 1.580 0.720 2.280 ;
        RECT  0.440 1.580 0.560 1.960 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.580 1.560 1.960 ;
        RECT  0.880 1.580 1.230 1.830 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.600 3.920 1.960 ;
        RECT  3.640 1.600 3.800 2.280 ;
        RECT  2.480 2.120 3.640 2.280 ;
        RECT  2.320 1.580 2.480 2.280 ;
        RECT  2.200 1.580 2.320 1.860 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.460 3.280 1.740 ;
        RECT  2.840 1.460 3.160 1.960 ;
        RECT  2.640 1.460 2.840 1.740 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.280 4.400 0.280 ;
        RECT  1.600 -0.280 1.880 0.390 ;
        RECT  0.880 -0.280 1.600 0.340 ;
        RECT  0.600 -0.280 0.880 0.980 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.920 3.320 4.400 3.880 ;
        RECT  3.640 2.800 3.920 3.880 ;
        RECT  2.240 3.320 3.640 3.880 ;
        RECT  1.960 2.760 2.240 3.880 ;
        RECT  0.560 3.320 1.960 3.880 ;
        RECT  0.280 2.470 0.560 3.880 ;
        RECT  0.000 3.320 0.280 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.920 0.700 4.200 0.980 ;
        RECT  3.240 0.700 3.920 0.860 ;
        RECT  2.960 0.700 3.240 0.980 ;
        RECT  2.280 0.700 2.960 0.860 ;
        RECT  2.000 0.700 2.280 1.300 ;
        RECT  1.360 1.140 2.000 1.300 ;
        RECT  1.080 0.700 1.360 1.300 ;
        RECT  0.400 1.140 1.080 1.300 ;
        RECT  0.120 1.020 0.400 1.300 ;
    END
END OAI22X2TR

MACRO OAI22X1TR
    CLASS CORE ;
    FOREIGN OAI22X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.150 2.320 2.370 ;
        RECT  2.080 1.150 2.240 2.680 ;
        RECT  1.830 1.150 2.080 1.310 ;
        RECT  1.350 2.520 2.080 2.680 ;
        RECT  1.550 1.030 1.830 1.310 ;
        RECT  1.070 2.120 1.350 2.870 ;
        END
        ANTENNADIFFAREA 2.592 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.560 0.540 1.880 ;
        RECT  0.320 1.240 0.330 1.880 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.360 1.020 1.640 ;
        RECT  0.700 1.360 0.860 2.360 ;
        RECT  0.480 2.040 0.700 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.480 1.920 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.540 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 -0.280 2.400 0.280 ;
        RECT  0.550 -0.280 0.830 0.400 ;
        RECT  0.000 -0.280 0.550 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.230 3.320 2.400 3.880 ;
        RECT  1.950 2.840 2.230 3.880 ;
        RECT  0.510 3.260 1.950 3.880 ;
        RECT  0.230 2.800 0.510 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.030 0.710 2.310 0.990 ;
        RECT  1.350 0.710 2.030 0.870 ;
        RECT  1.190 0.710 1.350 1.060 ;
        RECT  0.150 0.840 1.190 1.060 ;
    END
END OAI22X1TR

MACRO OAI222XLTR
    CLASS CORE ;
    FOREIGN OAI222XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.090 3.920 2.360 ;
        RECT  3.270 1.090 3.680 1.250 ;
        RECT  3.430 2.170 3.680 2.360 ;
        RECT  3.150 2.170 3.430 2.680 ;
        RECT  2.990 0.910 3.270 1.250 ;
        RECT  1.720 2.520 3.150 2.680 ;
        RECT  1.440 2.190 1.720 2.680 ;
        END
        ANTENNADIFFAREA 1.568 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.410 2.910 1.690 ;
        RECT  2.480 1.410 2.760 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.190 1.520 3.520 2.010 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.520 0.590 1.960 ;
        RECT  0.080 1.520 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.450 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.100 1.790 2.320 2.360 ;
        RECT  2.080 1.910 2.100 2.360 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.410 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.280 4.000 0.280 ;
        RECT  1.090 -0.280 1.370 0.800 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 3.320 4.000 3.880 ;
        RECT  2.280 2.840 2.560 3.880 ;
        RECT  0.880 3.320 2.280 3.880 ;
        RECT  0.600 2.320 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.470 0.570 3.750 0.930 ;
        RECT  2.790 0.570 3.470 0.730 ;
        RECT  2.510 0.570 2.790 0.930 ;
        RECT  1.830 0.570 2.510 0.730 ;
        RECT  2.030 0.910 2.310 1.250 ;
        RECT  0.850 1.090 2.030 1.250 ;
        RECT  1.550 0.570 1.830 0.930 ;
        RECT  0.570 0.830 0.850 1.250 ;
    END
END OAI222XLTR

MACRO OAI222X4TR
    CLASS CORE ;
    FOREIGN OAI222X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.580 0.840 4.720 2.070 ;
        RECT  4.360 0.440 4.580 3.160 ;
        RECT  4.300 0.440 4.360 1.340 ;
        RECT  4.300 1.880 4.360 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.640 2.400 2.360 ;
        RECT  2.080 2.040 2.240 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.640 3.350 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.150 0.890 1.560 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.640 2.070 1.880 ;
        RECT  1.680 1.640 1.920 2.070 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.800 1.520 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.060 -0.280 5.200 0.280 ;
        RECT  4.780 -0.280 5.060 0.670 ;
        RECT  4.060 -0.280 4.780 0.280 ;
        RECT  0.120 -0.280 4.060 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.060 3.320 5.200 3.880 ;
        RECT  4.780 2.230 5.060 3.880 ;
        RECT  4.100 3.320 4.780 3.880 ;
        RECT  3.820 2.440 4.100 3.880 ;
        RECT  2.250 3.260 3.820 3.880 ;
        RECT  1.970 3.200 2.250 3.880 ;
        RECT  0.610 3.260 1.970 3.880 ;
        RECT  0.330 2.610 0.610 3.880 ;
        RECT  0.000 3.320 0.330 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.080 1.470 4.180 1.750 ;
        RECT  3.920 1.000 4.080 2.280 ;
        RECT  3.620 1.000 3.920 1.160 ;
        RECT  3.620 2.120 3.920 2.280 ;
        RECT  3.540 1.320 3.760 1.660 ;
        RECT  3.340 0.880 3.620 1.160 ;
        RECT  3.340 2.120 3.620 3.100 ;
        RECT  2.760 1.320 3.540 1.480 ;
        RECT  2.810 2.520 3.090 2.800 ;
        RECT  2.720 2.520 2.810 2.680 ;
        RECT  2.720 1.200 2.760 1.480 ;
        RECT  2.560 1.200 2.720 2.680 ;
        RECT  2.480 1.200 2.560 1.480 ;
        RECT  1.410 2.520 2.560 2.680 ;
        RECT  2.000 1.170 2.280 1.450 ;
        RECT  1.360 1.290 2.000 1.450 ;
        RECT  1.480 0.700 1.760 0.980 ;
        RECT  0.830 0.820 1.480 0.980 ;
        RECT  1.130 2.520 1.410 2.800 ;
        RECT  1.070 1.290 1.360 1.570 ;
        RECT  0.610 0.700 0.830 0.980 ;
    END
END OAI222X4TR

MACRO OAI222X2TR
    CLASS CORE ;
    FOREIGN OAI222X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.880 1.030 6.040 2.680 ;
        RECT  5.680 1.030 5.880 1.560 ;
        RECT  5.120 2.520 5.880 2.680 ;
        RECT  5.500 1.030 5.680 1.330 ;
        RECT  4.860 1.170 5.500 1.330 ;
        RECT  4.840 2.520 5.120 2.810 ;
        RECT  4.580 1.050 4.860 1.330 ;
        RECT  3.440 2.520 4.840 2.680 ;
        RECT  3.160 2.520 3.440 2.800 ;
        RECT  1.720 2.520 3.160 2.680 ;
        RECT  1.440 2.520 1.720 2.800 ;
        END
        ANTENNADIFFAREA 7.164 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.600 1.820 5.720 2.100 ;
        RECT  5.440 1.820 5.600 2.360 ;
        RECT  4.720 2.200 5.440 2.360 ;
        RECT  4.480 1.510 4.720 2.360 ;
        RECT  4.300 1.510 4.480 1.790 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.640 5.280 1.960 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.730 2.320 2.010 ;
        RECT  2.040 1.730 2.200 2.330 ;
        RECT  1.120 2.170 2.040 2.330 ;
        RECT  0.920 1.640 1.120 2.330 ;
        RECT  0.480 1.640 0.920 1.980 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.640 1.760 2.010 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.020 1.710 4.140 1.990 ;
        RECT  3.860 1.710 4.020 2.360 ;
        RECT  3.680 2.040 3.860 2.360 ;
        RECT  2.800 2.120 3.680 2.280 ;
        RECT  2.640 1.730 2.800 2.280 ;
        RECT  2.520 1.730 2.640 2.010 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.590 3.520 1.960 ;
        RECT  2.960 1.590 3.280 1.870 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 -0.280 6.400 0.280 ;
        RECT  1.020 -0.280 2.160 0.340 ;
        RECT  0.380 -0.280 1.020 0.280 ;
        RECT  0.100 -0.280 0.380 0.340 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.960 3.320 6.400 3.880 ;
        RECT  5.680 2.930 5.960 3.880 ;
        RECT  4.280 3.320 5.680 3.880 ;
        RECT  4.000 2.840 4.280 3.880 ;
        RECT  2.560 3.260 4.000 3.880 ;
        RECT  2.280 2.840 2.560 3.880 ;
        RECT  0.880 3.260 2.280 3.880 ;
        RECT  0.600 2.700 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.040 0.630 6.300 0.870 ;
        RECT  5.340 0.710 6.040 0.870 ;
        RECT  5.060 0.710 5.340 1.010 ;
        RECT  3.660 0.730 3.940 1.370 ;
        RECT  3.020 0.730 3.660 0.890 ;
        RECT  2.740 0.730 3.020 1.430 ;
        RECT  1.720 0.770 2.740 0.930 ;
        RECT  1.440 0.650 1.720 0.930 ;
        RECT  0.800 0.770 1.440 0.930 ;
        RECT  0.520 0.650 0.800 0.930 ;
    END
END OAI222X2TR

MACRO OAI222X1TR
    CLASS CORE ;
    FOREIGN OAI222X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.090 3.920 2.360 ;
        RECT  3.270 1.090 3.680 1.250 ;
        RECT  3.430 2.170 3.680 2.360 ;
        RECT  3.150 2.170 3.430 2.960 ;
        RECT  2.990 0.970 3.270 1.250 ;
        RECT  1.720 2.520 3.150 2.680 ;
        RECT  1.440 2.520 1.720 2.800 ;
        END
        ANTENNADIFFAREA 4.044 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.410 2.850 1.960 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.640 3.520 2.010 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.520 0.590 1.800 ;
        RECT  0.080 1.520 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.450 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.790 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.410 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.280 4.000 0.280 ;
        RECT  1.090 -0.280 1.370 0.800 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.190 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 3.320 4.000 3.880 ;
        RECT  2.280 2.840 2.560 3.880 ;
        RECT  0.880 3.320 2.280 3.880 ;
        RECT  0.600 2.320 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.470 0.650 3.750 0.930 ;
        RECT  2.790 0.650 3.470 0.810 ;
        RECT  2.510 0.650 2.790 1.120 ;
        RECT  1.830 0.650 2.510 0.810 ;
        RECT  2.030 0.970 2.310 1.250 ;
        RECT  0.850 1.090 2.030 1.250 ;
        RECT  1.550 0.650 1.830 0.930 ;
        RECT  0.570 0.770 0.850 1.250 ;
    END
END OAI222X1TR

MACRO OAI221XLTR
    CLASS CORE ;
    FOREIGN OAI221XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.890 0.810 3.120 2.940 ;
        RECT  2.880 0.810 2.890 1.960 ;
        RECT  2.810 2.660 2.890 2.940 ;
        RECT  1.620 2.660 2.810 2.820 ;
        RECT  1.340 2.410 1.620 2.820 ;
        END
        ANTENNADIFFAREA 2.694 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 2.040 2.720 2.500 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.610 0.500 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 1.120 1.560 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.600 2.490 1.820 ;
        RECT  2.080 1.600 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.640 1.920 2.070 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.200 -0.280 3.200 0.280 ;
        RECT  0.920 -0.280 1.200 0.400 ;
        RECT  0.400 -0.280 0.920 0.280 ;
        RECT  0.120 -0.280 0.400 0.410 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.570 3.320 3.200 3.880 ;
        RECT  2.290 3.200 2.570 3.880 ;
        RECT  0.670 3.260 2.290 3.880 ;
        RECT  0.390 2.250 0.670 3.880 ;
        RECT  0.000 3.320 0.390 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.360 0.920 2.630 1.370 ;
        RECT  1.660 1.200 2.360 1.370 ;
        RECT  1.870 0.640 2.150 1.040 ;
        RECT  0.800 0.640 1.870 0.800 ;
        RECT  1.390 1.020 1.660 1.370 ;
        RECT  0.520 0.640 0.800 0.970 ;
    END
END OAI221XLTR

MACRO OAI221X4TR
    CLASS CORE ;
    FOREIGN OAI221X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.320 1.020 4.720 2.360 ;
        RECT  4.280 1.020 4.320 2.610 ;
        RECT  4.220 1.020 4.280 1.310 ;
        RECT  4.200 1.840 4.280 2.610 ;
        RECT  3.940 0.440 4.220 1.310 ;
        RECT  3.940 1.840 4.200 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.340 2.400 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.640 0.520 1.920 ;
        RECT  0.080 1.640 0.360 2.760 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.750 ;
        RECT  0.720 1.410 1.280 1.750 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.770 1.920 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.040 1.430 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.280 4.800 0.280 ;
        RECT  4.420 -0.280 4.700 0.670 ;
        RECT  3.740 -0.280 4.420 0.280 ;
        RECT  3.460 -0.280 3.740 1.130 ;
        RECT  1.200 -0.280 3.460 0.280 ;
        RECT  0.120 -0.280 1.200 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.480 2.520 4.700 3.880 ;
        RECT  3.700 3.320 4.480 3.880 ;
        RECT  3.420 3.200 3.700 3.880 ;
        RECT  2.900 3.320 3.420 3.880 ;
        RECT  2.620 3.200 2.900 3.880 ;
        RECT  1.920 3.260 2.620 3.880 ;
        RECT  1.640 3.200 1.920 3.880 ;
        RECT  0.400 3.260 1.640 3.880 ;
        RECT  0.120 3.200 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.780 1.470 4.120 1.680 ;
        RECT  3.620 1.470 3.780 2.750 ;
        RECT  3.260 1.470 3.620 1.630 ;
        RECT  3.020 2.470 3.620 2.750 ;
        RECT  2.810 2.030 3.460 2.310 ;
        RECT  3.100 0.440 3.260 1.630 ;
        RECT  2.980 0.440 3.100 1.130 ;
        RECT  2.810 1.470 2.920 1.750 ;
        RECT  2.650 1.470 2.810 2.730 ;
        RECT  2.440 2.570 2.650 2.730 ;
        RECT  2.160 2.570 2.440 2.890 ;
        RECT  0.900 2.610 2.160 2.890 ;
        RECT  1.780 0.850 2.060 1.130 ;
        RECT  0.790 0.850 1.780 1.010 ;
        RECT  0.520 0.850 0.790 1.130 ;
    END
END OAI221X4TR

MACRO OAI221X2TR
    CLASS CORE ;
    FOREIGN OAI221X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.220 1.150 4.320 2.760 ;
        RECT  4.120 1.030 4.220 2.850 ;
        RECT  3.940 1.030 4.120 1.310 ;
        RECT  3.940 2.440 4.120 2.850 ;
        RECT  2.900 2.540 3.940 2.760 ;
        RECT  2.620 2.540 2.900 3.160 ;
        RECT  1.210 2.540 2.620 2.700 ;
        RECT  0.930 2.470 1.210 2.750 ;
        END
        ANTENNADIFFAREA 5.22 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.600 3.960 1.960 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 1.580 1.860 1.880 ;
        RECT  0.720 1.720 1.590 1.880 ;
        RECT  0.350 1.240 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.420 1.560 ;
        END
        ANTENNAGATEAREA 0.3768 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 2.040 3.520 2.360 ;
        RECT  3.280 1.720 3.440 2.360 ;
        RECT  2.300 1.720 3.280 1.880 ;
        RECT  2.020 1.720 2.300 2.310 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 2.040 3.020 2.380 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.280 4.800 0.280 ;
        RECT  2.100 -0.280 2.380 0.400 ;
        RECT  1.380 -0.280 2.100 0.280 ;
        RECT  1.100 -0.280 1.380 0.720 ;
        RECT  0.410 -0.280 1.100 0.280 ;
        RECT  0.130 -0.280 0.410 1.080 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.420 2.920 4.700 3.880 ;
        RECT  3.700 3.320 4.420 3.880 ;
        RECT  3.420 2.990 3.700 3.880 ;
        RECT  2.100 3.320 3.420 3.880 ;
        RECT  1.820 2.930 2.100 3.880 ;
        RECT  0.370 3.260 1.820 3.880 ;
        RECT  0.090 2.340 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.420 0.650 4.700 0.930 ;
        RECT  3.730 0.650 4.420 0.810 ;
        RECT  3.610 0.650 3.730 1.310 ;
        RECT  3.450 0.500 3.610 1.310 ;
        RECT  2.770 0.500 3.450 0.660 ;
        RECT  2.970 0.820 3.250 1.560 ;
        RECT  1.860 1.260 2.970 1.420 ;
        RECT  2.610 0.500 2.770 1.100 ;
        RECT  2.490 0.820 2.610 1.100 ;
        RECT  1.700 0.440 1.860 1.420 ;
        RECT  1.580 0.440 1.700 1.060 ;
        RECT  0.900 0.900 1.580 1.060 ;
        RECT  0.620 0.440 0.900 1.060 ;
    END
END OAI221X2TR

MACRO OAI221X1TR
    CLASS CORE ;
    FOREIGN OAI221X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 1.640 3.520 2.760 ;
        RECT  3.280 0.710 3.440 2.760 ;
        RECT  3.000 0.710 3.280 1.250 ;
        RECT  3.020 2.200 3.280 2.680 ;
        RECT  1.640 2.520 3.020 2.680 ;
        END
        ANTENNADIFFAREA 3.662 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.780 1.530 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.240 0.660 1.490 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.240 1.230 1.560 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.220 1.480 2.460 2.360 ;
        RECT  2.080 2.040 2.220 2.360 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.520 2.060 1.800 ;
        RECT  1.610 1.520 1.790 2.360 ;
        RECT  1.280 2.040 1.610 2.360 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.380 -0.280 3.600 0.280 ;
        RECT  1.100 -0.280 1.380 0.340 ;
        RECT  0.380 -0.280 1.100 0.280 ;
        RECT  0.100 -0.280 0.380 1.080 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.780 3.320 3.600 3.880 ;
        RECT  2.440 2.840 2.780 3.880 ;
        RECT  1.080 3.320 2.440 3.880 ;
        RECT  0.800 1.940 1.080 3.880 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.580 0.650 2.740 1.310 ;
        RECT  1.780 1.150 2.580 1.310 ;
        RECT  2.100 0.500 2.260 0.930 ;
        RECT  0.800 0.500 2.100 0.660 ;
        RECT  1.620 1.030 1.780 1.310 ;
        RECT  0.640 0.500 0.800 1.080 ;
    END
END OAI221X1TR

MACRO OAI21XLTR
    CLASS CORE ;
    FOREIGN OAI21XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.240 1.920 2.360 ;
        RECT  1.680 0.730 1.840 2.360 ;
        RECT  1.560 0.730 1.680 1.040 ;
        RECT  0.960 2.180 1.680 2.360 ;
        END
        ANTENNADIFFAREA 1.066 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.800 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.620 0.600 1.910 ;
        RECT  0.330 1.240 0.340 1.910 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.640 1.120 1.960 ;
        RECT  0.760 1.600 0.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.280 2.000 0.280 ;
        RECT  0.600 -0.280 0.880 0.760 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 3.320 2.000 3.880 ;
        RECT  1.520 2.520 1.800 3.880 ;
        RECT  0.400 3.320 1.520 3.880 ;
        RECT  0.120 2.720 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 0.610 1.360 1.080 ;
        RECT  0.400 0.920 1.080 1.080 ;
        RECT  0.120 0.620 0.400 1.080 ;
    END
END OAI21XLTR

MACRO OAI21X4TR
    CLASS CORE ;
    FOREIGN OAI21X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.430 0.840 4.670 2.080 ;
        RECT  3.370 0.840 4.430 1.080 ;
        RECT  4.320 1.840 4.430 2.080 ;
        RECT  4.120 1.840 4.320 2.560 ;
        RECT  3.850 1.840 4.120 2.760 ;
        RECT  3.250 1.840 3.850 2.080 ;
        RECT  3.010 1.840 3.250 2.420 ;
        RECT  1.570 2.180 3.010 2.420 ;
        RECT  1.290 2.180 1.570 3.020 ;
        END
        ANTENNADIFFAREA 8.294 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.240 4.270 1.600 ;
        END
        ANTENNAGATEAREA 0.6024 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.240 2.530 1.660 ;
        RECT  0.690 1.240 1.890 1.400 ;
        RECT  0.320 1.240 0.690 1.900 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.672 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.360 2.970 1.640 ;
        RECT  2.690 1.360 2.850 1.980 ;
        RECT  1.480 1.820 2.690 1.980 ;
        RECT  0.880 1.640 1.480 1.980 ;
        END
        ANTENNAGATEAREA 0.672 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.770 -0.280 4.800 0.280 ;
        RECT  1.570 -0.280 2.770 0.340 ;
        RECT  0.930 -0.280 1.570 0.280 ;
        RECT  0.650 -0.280 0.930 0.340 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.670 3.320 4.800 3.880 ;
        RECT  4.390 2.720 4.670 3.880 ;
        RECT  3.650 3.260 4.390 3.880 ;
        RECT  3.430 2.480 3.650 3.880 ;
        RECT  2.370 3.320 3.430 3.880 ;
        RECT  2.090 2.630 2.370 3.880 ;
        RECT  0.770 3.320 2.090 3.880 ;
        RECT  0.490 2.190 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.850 0.480 4.130 0.670 ;
        RECT  3.170 0.480 3.850 0.640 ;
        RECT  3.010 0.480 3.170 1.080 ;
        RECT  2.890 0.810 3.010 1.080 ;
        RECT  2.260 0.910 2.890 1.080 ;
        RECT  1.970 0.800 2.260 1.080 ;
        RECT  1.330 0.920 1.970 1.080 ;
        RECT  1.050 0.800 1.330 1.080 ;
        RECT  0.410 0.920 1.050 1.080 ;
        RECT  0.130 0.440 0.410 1.080 ;
    END
END OAI21X4TR

MACRO OAI21X2TR
    CLASS CORE ;
    FOREIGN OAI21X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.240 3.160 1.560 ;
        RECT  2.960 1.030 3.040 2.280 ;
        RECT  2.880 1.030 2.960 2.400 ;
        RECT  2.720 1.030 2.880 1.310 ;
        RECT  2.680 2.120 2.880 2.400 ;
        RECT  1.480 2.120 2.680 2.280 ;
        RECT  1.200 2.120 1.480 2.740 ;
        END
        ANTENNADIFFAREA 3.762 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.490 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.240 2.160 1.640 ;
        RECT  0.720 1.240 1.890 1.400 ;
        RECT  0.390 1.240 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.580 1.680 1.960 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.280 3.600 0.280 ;
        RECT  1.720 -0.280 2.000 0.760 ;
        RECT  0.950 -0.280 1.720 0.280 ;
        RECT  0.680 -0.280 0.950 0.760 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.480 3.320 3.600 3.880 ;
        RECT  3.200 1.910 3.480 3.880 ;
        RECT  2.360 3.320 3.200 3.880 ;
        RECT  2.080 2.460 2.360 3.880 ;
        RECT  0.690 3.320 2.080 3.880 ;
        RECT  0.410 1.910 0.690 3.880 ;
        RECT  0.000 3.320 0.410 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.200 0.710 3.480 0.990 ;
        RECT  2.520 0.710 3.200 0.870 ;
        RECT  2.240 0.710 2.520 1.080 ;
        RECT  1.480 0.920 2.240 1.080 ;
        RECT  1.200 0.800 1.480 1.080 ;
        RECT  0.440 0.920 1.200 1.080 ;
        RECT  0.160 0.800 0.440 1.080 ;
    END
END OAI21X2TR

MACRO OAI21X1TR
    CLASS CORE ;
    FOREIGN OAI21X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.640 1.920 2.760 ;
        RECT  1.680 1.030 1.840 2.760 ;
        RECT  1.560 1.030 1.680 1.310 ;
        RECT  1.240 2.520 1.680 2.680 ;
        RECT  0.960 2.520 1.240 2.810 ;
        END
        ANTENNADIFFAREA 2.56 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.520 1.520 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.640 0.600 1.960 ;
        RECT  0.080 1.640 0.380 2.760 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.640 1.120 1.960 ;
        RECT  0.760 1.600 0.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.280 2.000 0.280 ;
        RECT  0.600 -0.280 0.880 0.990 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 3.320 2.000 3.880 ;
        RECT  1.520 2.930 1.800 3.880 ;
        RECT  0.400 3.320 1.520 3.880 ;
        RECT  0.130 2.920 0.400 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 1.030 1.360 1.310 ;
        RECT  0.400 1.150 1.080 1.310 ;
        RECT  0.120 1.030 0.400 1.310 ;
    END
END OAI21X1TR

MACRO OAI211XLTR
    CLASS CORE ;
    FOREIGN OAI211XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.440 2.320 1.560 ;
        RECT  2.120 0.440 2.310 2.330 ;
        RECT  2.080 0.440 2.120 1.560 ;
        RECT  2.080 2.080 2.120 2.330 ;
        RECT  1.120 2.120 2.080 2.280 ;
        RECT  0.960 2.120 1.120 2.470 ;
        END
        ANTENNADIFFAREA 2.549 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 1.920 1.960 ;
        RECT  1.340 1.640 1.680 1.880 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.600 2.120 2.780 ;
        RECT  1.280 2.440 1.520 2.780 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.520 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.880 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.280 2.400 0.280 ;
        RECT  0.640 -0.280 0.920 0.520 ;
        RECT  0.000 -0.280 0.640 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 3.320 2.400 3.880 ;
        RECT  0.390 3.260 1.760 3.880 ;
        RECT  0.110 2.250 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.370 0.920 1.540 1.080 ;
        RECT  0.090 0.920 0.370 1.200 ;
    END
END OAI211XLTR

MACRO OAI211X4TR
    CLASS CORE ;
    FOREIGN OAI211X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.040 3.520 2.070 ;
        RECT  3.280 0.440 3.430 3.160 ;
        RECT  3.150 0.440 3.280 1.310 ;
        RECT  3.150 1.910 3.280 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.200 1.520 1.560 ;
        RECT  1.280 1.200 1.500 1.670 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 1.990 2.030 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.370 0.570 1.630 ;
        RECT  0.340 1.240 0.350 1.630 ;
        RECT  0.080 1.240 0.340 2.370 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.360 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 -0.280 4.000 0.280 ;
        RECT  3.630 -0.280 3.910 0.670 ;
        RECT  2.950 -0.280 3.630 0.280 ;
        RECT  2.670 -0.280 2.950 0.840 ;
        RECT  0.850 -0.280 2.670 0.340 ;
        RECT  0.570 -0.280 0.850 1.130 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 3.320 4.000 3.880 ;
        RECT  3.630 2.230 3.910 3.880 ;
        RECT  2.950 3.320 3.630 3.880 ;
        RECT  2.670 2.910 2.950 3.880 ;
        RECT  1.730 3.260 2.670 3.880 ;
        RECT  1.450 2.800 1.730 3.880 ;
        RECT  0.390 3.260 1.450 3.880 ;
        RECT  0.110 2.800 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.990 1.470 3.120 1.750 ;
        RECT  2.830 1.000 2.990 2.670 ;
        RECT  2.470 1.000 2.830 1.160 ;
        RECT  2.430 2.510 2.830 2.670 ;
        RECT  2.450 1.320 2.610 2.350 ;
        RECT  2.310 0.560 2.470 1.160 ;
        RECT  2.100 1.320 2.450 1.480 ;
        RECT  2.090 2.190 2.450 2.350 ;
        RECT  2.270 2.510 2.430 2.930 ;
        RECT  2.190 0.560 2.310 0.850 ;
        RECT  2.150 2.650 2.270 2.930 ;
        RECT  1.820 1.030 2.100 1.480 ;
        RECT  1.810 2.190 2.090 2.470 ;
        RECT  1.290 2.190 1.810 2.350 ;
        RECT  1.130 2.190 1.290 2.900 ;
        RECT  0.950 2.620 1.130 2.900 ;
    END
END OAI211X4TR

MACRO OAI211X2TR
    CLASS CORE ;
    FOREIGN OAI211X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.000 3.920 2.440 ;
        RECT  3.560 1.000 3.760 1.160 ;
        RECT  3.160 2.280 3.760 2.440 ;
        RECT  3.280 0.840 3.560 1.160 ;
        RECT  3.080 0.840 3.280 1.080 ;
        RECT  2.880 2.280 3.160 3.100 ;
        RECT  2.800 0.800 3.080 1.080 ;
        RECT  2.200 2.280 2.880 2.440 ;
        RECT  1.920 2.260 2.200 2.890 ;
        RECT  0.560 2.260 1.920 2.420 ;
        RECT  0.280 2.260 0.560 2.890 ;
        END
        ANTENNADIFFAREA 6.442 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.840 3.600 2.120 ;
        RECT  2.720 1.960 3.320 2.120 ;
        RECT  2.440 1.490 2.720 2.120 ;
        RECT  2.200 1.490 2.440 1.770 ;
        END
        ANTENNAGATEAREA 0.2928 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.120 1.800 ;
        END
        ANTENNAGATEAREA 0.2928 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.500 1.560 1.780 ;
        RECT  0.880 1.240 1.160 1.780 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.500 2.000 1.770 ;
        RECT  1.720 1.500 1.880 2.100 ;
        RECT  0.720 1.940 1.720 2.100 ;
        RECT  0.440 1.640 0.720 2.100 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.280 4.000 0.280 ;
        RECT  1.480 -0.280 1.760 0.400 ;
        RECT  0.960 -0.280 1.480 0.280 ;
        RECT  0.680 -0.280 0.960 0.400 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 3.320 4.000 3.880 ;
        RECT  2.400 2.600 2.680 3.880 ;
        RECT  1.360 3.320 2.400 3.880 ;
        RECT  1.080 2.610 1.360 3.880 ;
        RECT  0.000 3.320 1.080 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.800 2.280 1.080 ;
        RECT  1.360 0.920 2.000 1.080 ;
        RECT  1.080 0.800 1.360 1.080 ;
        RECT  0.440 0.920 1.080 1.080 ;
        RECT  0.160 0.800 0.440 1.080 ;
    END
END OAI211X2TR

MACRO OAI211X1TR
    CLASS CORE ;
    FOREIGN OAI211X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.440 2.320 1.560 ;
        RECT  2.120 0.440 2.280 2.400 ;
        RECT  2.080 0.440 2.120 1.560 ;
        RECT  2.070 2.080 2.120 2.400 ;
        RECT  2.060 2.120 2.070 2.400 ;
        RECT  1.120 2.120 2.060 2.280 ;
        RECT  0.960 2.120 1.120 2.900 ;
        END
        ANTENNADIFFAREA 4.112 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 1.920 1.960 ;
        RECT  1.340 1.640 1.680 1.920 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.820 2.120 3.000 ;
        RECT  1.280 2.440 1.520 3.000 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.590 0.540 1.900 ;
        RECT  0.340 1.240 0.360 1.900 ;
        RECT  0.080 1.240 0.340 2.360 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.880 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.280 2.400 0.280 ;
        RECT  0.630 -0.280 0.930 0.760 ;
        RECT  0.000 -0.280 0.630 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.830 3.320 2.400 3.880 ;
        RECT  0.390 3.260 1.830 3.880 ;
        RECT  0.110 2.570 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.370 0.920 1.500 1.080 ;
        RECT  0.090 0.600 0.370 1.080 ;
    END
END OAI211X1TR

MACRO OA22XLTR
    CLASS CORE ;
    FOREIGN OA22XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.680 2.720 1.960 ;
        RECT  2.470 0.680 2.630 3.160 ;
        RECT  2.250 0.680 2.470 0.940 ;
        RECT  2.270 2.880 2.470 3.160 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.040 1.920 2.360 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.050 1.520 1.630 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.170 0.430 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 2.040 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.280 2.800 0.280 ;
        RECT  1.650 -0.280 2.000 0.560 ;
        RECT  0.000 -0.280 1.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 3.320 2.800 3.880 ;
        RECT  1.790 2.880 2.070 3.880 ;
        RECT  0.350 3.320 1.790 3.880 ;
        RECT  0.090 2.520 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.140 2.110 2.300 2.720 ;
        RECT  1.170 2.560 2.140 2.720 ;
        RECT  1.970 1.630 2.030 1.870 ;
        RECT  1.810 0.720 1.970 1.870 ;
        RECT  1.370 0.720 1.810 0.880 ;
        RECT  1.760 1.630 1.810 1.870 ;
        RECT  1.090 0.520 1.370 0.880 ;
        RECT  0.890 2.560 1.170 2.840 ;
        RECT  0.370 0.520 1.090 0.680 ;
        RECT  0.670 2.560 0.890 2.720 ;
        RECT  0.670 0.990 0.750 1.880 ;
        RECT  0.590 0.990 0.670 2.720 ;
        RECT  0.510 1.720 0.590 2.720 ;
        RECT  0.090 0.480 0.370 0.680 ;
    END
END OA22XLTR

MACRO OA22X4TR
    CLASS CORE ;
    FOREIGN OA22X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.210 3.520 2.680 ;
        RECT  3.360 0.440 3.430 2.680 ;
        RECT  3.280 0.440 3.360 3.160 ;
        RECT  3.150 0.440 3.280 1.450 ;
        RECT  3.080 2.440 3.280 3.160 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.760 1.920 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.640 2.320 1.960 ;
        RECT  2.080 1.600 2.190 1.960 ;
        RECT  1.910 1.600 2.080 1.880 ;
        END
        ANTENNAGATEAREA 0.2376 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.570 0.760 1.970 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.040 1.920 2.360 ;
        RECT  1.590 1.460 1.750 2.360 ;
        RECT  1.470 1.460 1.590 1.740 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 -0.280 4.000 0.280 ;
        RECT  3.630 -0.280 3.910 1.050 ;
        RECT  2.950 -0.280 3.630 0.280 ;
        RECT  2.670 -0.280 2.950 1.070 ;
        RECT  1.990 -0.280 2.670 0.280 ;
        RECT  1.710 -0.280 1.990 0.800 ;
        RECT  0.000 -0.280 1.710 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 3.320 4.000 3.880 ;
        RECT  3.560 2.930 3.840 3.880 ;
        RECT  2.860 3.320 3.560 3.880 ;
        RECT  2.540 2.440 2.860 3.880 ;
        RECT  1.110 3.320 2.540 3.880 ;
        RECT  0.830 2.220 1.110 3.880 ;
        RECT  0.000 3.320 0.830 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.080 1.620 3.100 1.970 ;
        RECT  2.920 1.620 3.080 2.280 ;
        RECT  2.240 2.120 2.920 2.280 ;
        RECT  2.320 0.520 2.470 0.920 ;
        RECT  2.160 0.520 2.320 1.300 ;
        RECT  2.080 2.120 2.240 2.680 ;
        RECT  1.520 1.140 2.160 1.300 ;
        RECT  1.950 2.520 2.080 2.680 ;
        RECT  1.670 2.520 1.950 3.080 ;
        RECT  1.430 2.520 1.670 2.680 ;
        RECT  1.240 0.500 1.520 1.300 ;
        RECT  1.270 1.900 1.430 2.680 ;
        RECT  1.080 1.900 1.270 2.060 ;
        RECT  0.550 0.500 1.240 0.660 ;
        RECT  0.920 0.930 1.080 2.060 ;
        RECT  0.750 0.930 0.920 1.250 ;
        RECT  0.270 0.500 0.550 1.280 ;
    END
END OA22X4TR

MACRO OA22X2TR
    CLASS CORE ;
    FOREIGN OA22X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 0.500 3.120 3.160 ;
        RECT  2.830 0.500 2.920 1.260 ;
        RECT  2.880 2.040 2.920 3.160 ;
        RECT  2.720 2.440 2.880 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.440 2.360 1.960 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.680 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.240 0.420 1.610 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.790 1.520 2.360 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.280 3.200 0.280 ;
        RECT  1.510 -0.280 2.530 0.520 ;
        RECT  0.000 -0.280 1.510 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 3.320 3.200 3.880 ;
        RECT  2.080 2.490 2.370 3.880 ;
        RECT  0.420 3.320 2.080 3.880 ;
        RECT  0.140 2.520 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.680 1.470 2.750 1.800 ;
        RECT  2.520 1.470 2.680 2.280 ;
        RECT  1.840 2.120 2.520 2.280 ;
        RECT  1.280 0.920 2.220 1.080 ;
        RECT  1.680 2.120 1.840 2.680 ;
        RECT  1.340 2.520 1.680 2.680 ;
        RECT  1.060 2.520 1.340 2.800 ;
        RECT  1.270 0.920 1.280 1.350 ;
        RECT  1.110 0.710 1.270 1.350 ;
        RECT  0.370 0.710 1.110 0.870 ;
        RECT  0.740 2.520 1.060 2.680 ;
        RECT  0.740 1.030 0.850 1.310 ;
        RECT  0.580 1.030 0.740 2.680 ;
        RECT  0.090 0.710 0.370 1.050 ;
    END
END OA22X2TR

MACRO OA22X1TR
    CLASS CORE ;
    FOREIGN OA22X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.680 2.720 1.960 ;
        RECT  2.470 0.680 2.630 3.160 ;
        RECT  2.250 0.680 2.470 0.940 ;
        RECT  2.270 2.880 2.470 3.160 ;
        END
        ANTENNADIFFAREA 1.783 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.040 1.920 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.050 1.520 1.630 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.170 0.430 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 2.040 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.280 2.800 0.280 ;
        RECT  1.650 -0.280 2.000 0.560 ;
        RECT  0.000 -0.280 1.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 3.320 2.800 3.880 ;
        RECT  1.790 2.880 2.070 3.880 ;
        RECT  0.350 3.320 1.790 3.880 ;
        RECT  0.090 2.460 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.140 2.110 2.300 2.720 ;
        RECT  1.170 2.560 2.140 2.720 ;
        RECT  1.970 1.630 2.040 1.870 ;
        RECT  1.810 0.720 1.970 1.870 ;
        RECT  1.370 0.720 1.810 0.880 ;
        RECT  1.760 1.630 1.810 1.870 ;
        RECT  1.090 0.520 1.370 0.880 ;
        RECT  0.890 2.560 1.170 2.840 ;
        RECT  0.370 0.520 1.090 0.680 ;
        RECT  0.670 2.560 0.890 2.720 ;
        RECT  0.670 0.990 0.750 1.880 ;
        RECT  0.590 0.990 0.670 2.720 ;
        RECT  0.510 1.720 0.590 2.720 ;
        RECT  0.090 0.440 0.370 0.680 ;
    END
END OA22X1TR

MACRO OA21XLTR
    CLASS CORE ;
    FOREIGN OA21XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.440 2.320 2.760 ;
        RECT  1.940 0.440 2.160 0.720 ;
        RECT  2.080 1.640 2.160 2.760 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.470 1.420 1.750 ;
        RECT  1.120 0.840 1.280 1.750 ;
        RECT  0.880 0.840 1.120 1.160 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.400 0.910 1.650 ;
        RECT  0.480 1.240 0.720 1.650 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.660 -0.280 2.400 0.280 ;
        RECT  1.380 -0.280 1.660 0.610 ;
        RECT  0.650 -0.280 1.380 0.280 ;
        RECT  0.370 -0.280 0.650 1.080 ;
        RECT  0.000 -0.280 0.370 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 3.320 2.400 3.880 ;
        RECT  1.510 2.230 1.790 3.880 ;
        RECT  0.370 3.320 1.510 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.820 1.390 1.920 1.710 ;
        RECT  1.810 1.030 1.820 1.710 ;
        RECT  1.650 1.030 1.810 2.070 ;
        RECT  1.440 1.030 1.650 1.310 ;
        RECT  1.160 1.910 1.650 2.070 ;
        RECT  1.000 1.910 1.160 2.300 ;
    END
END OA21XLTR

MACRO OA21X4TR
    CLASS CORE ;
    FOREIGN OA21X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.840 3.300 2.760 ;
        RECT  2.980 1.510 3.210 2.760 ;
        RECT  2.820 1.510 2.980 1.750 ;
        RECT  2.540 0.520 2.820 1.750 ;
        RECT  2.380 1.510 2.540 1.750 ;
        RECT  2.140 1.510 2.380 2.760 ;
        RECT  2.060 1.840 2.140 2.760 ;
        END
        ANTENNADIFFAREA 4.868 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.540 1.540 1.960 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.720 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.340 -0.280 3.600 0.280 ;
        RECT  3.060 -0.280 3.340 1.310 ;
        RECT  2.340 -0.280 3.060 0.280 ;
        RECT  2.060 -0.280 2.340 1.260 ;
        RECT  0.900 -0.280 2.060 0.280 ;
        RECT  0.620 -0.280 0.900 0.670 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.820 3.320 3.600 3.880 ;
        RECT  2.540 1.910 2.820 3.880 ;
        RECT  1.780 3.320 2.540 3.880 ;
        RECT  1.500 2.480 1.780 3.880 ;
        RECT  0.420 3.320 1.500 3.880 ;
        RECT  0.140 2.120 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 1.460 1.980 1.680 ;
        RECT  1.720 0.690 1.900 2.280 ;
        RECT  1.580 0.690 1.720 1.310 ;
        RECT  1.300 2.120 1.720 2.280 ;
        RECT  1.100 0.500 1.380 1.080 ;
        RECT  1.020 2.120 1.300 2.930 ;
        RECT  0.420 0.920 1.100 1.080 ;
        RECT  0.140 0.440 0.420 1.080 ;
    END
END OA21X4TR

MACRO OA21X2TR
    CLASS CORE ;
    FOREIGN OA21X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.440 2.720 2.170 ;
        RECT  2.160 0.840 2.480 1.090 ;
        RECT  2.180 2.010 2.480 2.170 ;
        RECT  2.020 2.010 2.180 2.810 ;
        RECT  1.890 0.440 2.160 1.090 ;
        RECT  1.860 2.530 2.020 2.810 ;
        END
        ANTENNADIFFAREA 2.561 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 0.840 1.620 1.160 ;
        RECT  1.380 1.770 1.500 2.050 ;
        RECT  1.220 0.840 1.380 2.050 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.320 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.560 1.020 1.960 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 -0.280 2.800 0.280 ;
        RECT  0.540 -0.280 0.820 1.090 ;
        RECT  0.000 -0.280 0.540 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 3.320 2.800 3.880 ;
        RECT  2.340 2.420 2.620 3.880 ;
        RECT  1.620 3.260 2.340 3.880 ;
        RECT  1.340 3.200 1.620 3.880 ;
        RECT  0.420 3.260 1.340 3.880 ;
        RECT  0.140 3.200 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.820 1.560 2.160 1.850 ;
        RECT  1.660 1.330 1.820 2.370 ;
        RECT  1.540 1.330 1.660 1.610 ;
        RECT  1.220 2.210 1.660 2.370 ;
        RECT  0.940 2.210 1.220 2.580 ;
    END
END OA21X2TR

MACRO OA21X1TR
    CLASS CORE ;
    FOREIGN OA21X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.240 2.720 2.390 ;
        RECT  2.310 0.770 2.470 2.390 ;
        RECT  2.230 0.770 2.310 0.930 ;
        RECT  2.160 1.870 2.310 2.390 ;
        RECT  1.950 0.570 2.230 0.930 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.360 1.630 1.640 ;
        RECT  1.350 0.840 1.560 1.640 ;
        RECT  1.240 0.840 1.350 1.160 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.440 0.370 1.640 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.510 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.280 2.800 0.280 ;
        RECT  2.430 -0.280 2.710 0.610 ;
        RECT  0.870 -0.280 2.430 0.280 ;
        RECT  0.590 -0.280 0.870 1.310 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.920 3.320 2.800 3.880 ;
        RECT  1.640 2.250 1.920 3.880 ;
        RECT  0.510 3.320 1.640 3.880 ;
        RECT  0.230 2.070 0.510 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.070 1.430 2.150 1.710 ;
        RECT  1.950 1.090 2.070 1.710 ;
        RECT  1.790 1.090 1.950 1.960 ;
        RECT  1.480 1.800 1.790 1.960 ;
        RECT  1.320 1.800 1.480 2.290 ;
        RECT  1.030 2.130 1.320 2.290 ;
    END
END OA21X1TR

MACRO NOR4BBXLTR
    CLASS CORE ;
    FOREIGN NOR4BBXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.710 3.520 2.760 ;
        RECT  2.430 0.710 3.360 0.870 ;
        RECT  2.760 2.600 3.360 2.760 ;
        RECT  2.310 2.440 2.760 2.760 ;
        RECT  2.150 0.510 2.430 0.870 ;
        RECT  1.430 0.710 2.150 0.870 ;
        RECT  1.150 0.710 1.430 1.080 ;
        END
        ANTENNADIFFAREA 2.384 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.720 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.430 1.670 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.560 3.200 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.460 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.280 3.600 0.280 ;
        RECT  2.840 -0.280 3.140 0.540 ;
        RECT  1.870 -0.280 2.840 0.280 ;
        RECT  1.590 -0.280 1.870 0.400 ;
        RECT  0.870 -0.280 1.590 0.340 ;
        RECT  0.590 -0.280 0.870 0.810 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.200 3.320 3.600 3.880 ;
        RECT  2.920 2.930 3.200 3.880 ;
        RECT  1.150 3.260 2.920 3.880 ;
        RECT  0.870 2.440 1.150 3.880 ;
        RECT  0.000 3.320 0.870 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 1.030 3.200 1.400 ;
        RECT  2.920 2.120 3.200 2.400 ;
        RECT  2.720 1.240 2.920 1.400 ;
        RECT  2.720 2.120 2.920 2.280 ;
        RECT  2.560 1.240 2.720 2.280 ;
        RECT  2.190 1.240 2.560 1.400 ;
        RECT  2.110 1.770 2.390 2.280 ;
        RECT  1.910 1.240 2.190 1.520 ;
        RECT  0.480 2.120 2.110 2.280 ;
        RECT  0.310 2.120 0.480 2.400 ;
        RECT  0.310 1.030 0.370 1.310 ;
        RECT  0.150 1.030 0.310 2.400 ;
        RECT  0.090 1.030 0.150 1.310 ;
    END
END NOR4BBXLTR

MACRO NOR4BBX4TR
    CLASS CORE ;
    FOREIGN NOR4BBX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.420 0.500 8.660 3.060 ;
        RECT  1.050 0.500 8.420 0.740 ;
        RECT  7.920 2.820 8.420 3.060 ;
        RECT  7.680 1.840 7.920 3.060 ;
        RECT  6.120 2.820 7.680 3.060 ;
        RECT  5.840 2.820 6.120 3.100 ;
        RECT  2.400 2.820 5.840 3.060 ;
        RECT  2.120 2.820 2.400 3.100 ;
        END
        ANTENNADIFFAREA 9.771 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.860 7.500 2.660 ;
        RECT  4.390 2.500 7.340 2.660 ;
        RECT  4.110 2.140 4.390 2.660 ;
        RECT  1.560 2.440 4.110 2.660 ;
        RECT  1.480 2.440 1.560 2.760 ;
        RECT  1.240 2.140 1.480 2.760 ;
        RECT  1.160 2.140 1.240 2.300 ;
        RECT  1.000 1.670 1.160 2.300 ;
        RECT  0.880 1.670 1.000 1.910 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.940 1.840 7.100 2.340 ;
        RECT  5.200 2.180 6.940 2.340 ;
        RECT  5.040 1.580 5.200 2.340 ;
        RECT  4.840 1.580 5.040 1.980 ;
        RECT  3.320 1.820 4.840 1.980 ;
        RECT  3.040 1.700 3.320 1.980 ;
        RECT  1.480 1.820 3.040 1.980 ;
        RECT  1.320 1.220 1.480 1.980 ;
        RECT  1.150 1.220 1.320 1.380 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.260 1.240 7.520 1.700 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.380 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.110 -0.280 8.800 0.280 ;
        RECT  1.570 -0.280 7.110 0.340 ;
        RECT  0.850 -0.280 1.570 0.280 ;
        RECT  0.570 -0.280 0.850 0.660 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 3.320 8.800 3.880 ;
        RECT  7.520 3.220 7.800 3.880 ;
        RECT  3.960 3.320 7.520 3.880 ;
        RECT  3.680 3.220 3.960 3.880 ;
        RECT  0.890 3.320 3.680 3.880 ;
        RECT  0.610 2.460 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.100 0.910 8.260 2.620 ;
        RECT  7.100 0.910 8.100 1.080 ;
        RECT  6.940 0.910 7.100 1.600 ;
        RECT  6.730 1.440 6.940 1.600 ;
        RECT  6.570 1.440 6.730 1.960 ;
        RECT  6.510 0.900 6.670 1.280 ;
        RECT  5.970 1.800 6.570 1.960 ;
        RECT  2.450 0.900 6.510 1.060 ;
        RECT  5.790 1.260 5.970 1.960 ;
        RECT  2.880 1.260 5.790 1.420 ;
        RECT  2.650 1.260 2.880 1.660 ;
        RECT  1.920 1.500 2.650 1.660 ;
        RECT  2.210 0.900 2.450 1.280 ;
        RECT  0.380 0.900 2.210 1.060 ;
        RECT  1.640 1.300 1.920 1.660 ;
        RECT  0.370 0.500 0.380 1.060 ;
        RECT  0.270 0.500 0.370 1.200 ;
        RECT  0.270 2.190 0.360 3.080 ;
        RECT  0.110 0.500 0.270 3.080 ;
    END
END NOR4BBX4TR

MACRO NOR4BBX2TR
    CLASS CORE ;
    FOREIGN NOR4BBX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 0.520 6.320 3.080 ;
        RECT  4.580 0.520 6.080 0.720 ;
        RECT  3.240 2.920 6.080 3.080 ;
        RECT  4.300 0.440 4.580 0.720 ;
        RECT  3.240 0.560 4.300 0.720 ;
        RECT  2.960 0.440 3.240 0.720 ;
        RECT  2.960 2.840 3.240 3.080 ;
        RECT  2.200 0.560 2.960 0.720 ;
        RECT  1.920 0.440 2.200 0.720 ;
        END
        ANTENNADIFFAREA 5.128 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.140 1.520 4.430 1.740 ;
        RECT  2.720 1.580 4.140 1.740 ;
        RECT  2.620 1.580 2.720 1.960 ;
        RECT  2.480 1.530 2.620 1.960 ;
        RECT  1.720 1.530 2.480 1.690 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.910 2.040 5.120 2.360 ;
        RECT  4.880 1.520 4.910 2.360 ;
        RECT  4.630 1.520 4.880 2.280 ;
        RECT  4.160 2.120 4.630 2.280 ;
        RECT  3.850 1.900 4.160 2.280 ;
        RECT  2.300 2.120 3.850 2.280 ;
        RECT  2.040 1.880 2.300 2.280 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.640 0.760 1.960 ;
        RECT  0.400 1.600 0.560 1.960 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.640 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.180 -0.280 6.400 0.280 ;
        RECT  5.900 -0.280 6.180 0.300 ;
        RECT  5.100 -0.280 5.900 0.280 ;
        RECT  4.820 -0.280 5.100 0.360 ;
        RECT  3.930 -0.280 4.820 0.280 ;
        RECT  3.650 -0.280 3.930 0.360 ;
        RECT  2.720 -0.280 3.650 0.280 ;
        RECT  2.440 -0.280 2.720 0.360 ;
        RECT  1.680 -0.280 2.440 0.280 ;
        RECT  1.400 -0.280 1.680 0.360 ;
        RECT  0.860 -0.280 1.400 0.340 ;
        RECT  0.580 -0.280 0.860 0.930 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 3.320 6.400 3.880 ;
        RECT  4.490 3.240 4.830 3.880 ;
        RECT  1.800 3.320 4.490 3.880 ;
        RECT  1.360 3.150 1.800 3.880 ;
        RECT  0.860 3.260 1.360 3.880 ;
        RECT  0.580 2.120 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.640 0.880 5.800 2.680 ;
        RECT  3.440 0.880 5.640 1.040 ;
        RECT  1.390 2.520 5.640 2.680 ;
        RECT  3.840 1.200 5.420 1.360 ;
        RECT  3.620 1.200 3.840 1.420 ;
        RECT  2.960 1.260 3.620 1.420 ;
        RECT  3.160 0.880 3.440 1.100 ;
        RECT  1.340 0.880 3.160 1.040 ;
        RECT  2.820 1.200 2.960 1.420 ;
        RECT  0.380 1.200 2.820 1.360 ;
        RECT  1.340 2.120 1.390 2.680 ;
        RECT  1.060 0.760 1.340 1.040 ;
        RECT  1.060 2.120 1.340 2.900 ;
        RECT  0.240 0.930 0.380 1.360 ;
        RECT  0.240 2.120 0.380 2.900 ;
        RECT  0.080 0.930 0.240 2.900 ;
    END
END NOR4BBX2TR

MACRO NOR4BBX1TR
    CLASS CORE ;
    FOREIGN NOR4BBX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.330 0.710 3.490 2.760 ;
        RECT  2.210 0.710 3.330 0.870 ;
        RECT  2.480 2.600 3.330 2.760 ;
        RECT  2.040 2.440 2.480 3.110 ;
        RECT  1.930 0.590 2.210 0.870 ;
        RECT  1.290 0.710 1.930 0.870 ;
        RECT  1.010 0.710 1.290 0.990 ;
        END
        ANTENNADIFFAREA 3.576 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.520 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.160 1.560 1.600 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.640 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 -0.280 3.600 0.280 ;
        RECT  2.480 -0.280 2.760 0.400 ;
        RECT  1.690 -0.280 2.480 0.280 ;
        RECT  0.770 -0.280 1.690 0.340 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 3.320 3.600 3.880 ;
        RECT  2.890 3.080 3.170 3.880 ;
        RECT  1.040 3.320 2.890 3.880 ;
        RECT  0.760 2.840 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.890 2.120 3.170 2.440 ;
        RECT  2.880 1.030 3.160 1.310 ;
        RECT  2.600 2.120 2.890 2.280 ;
        RECT  2.600 1.140 2.880 1.310 ;
        RECT  2.440 1.140 2.600 2.280 ;
        RECT  2.020 1.140 2.440 1.300 ;
        RECT  2.000 1.580 2.280 1.860 ;
        RECT  1.740 1.140 2.020 1.420 ;
        RECT  1.880 1.700 2.000 1.860 ;
        RECT  1.720 1.700 1.880 2.680 ;
        RECT  0.680 2.490 1.720 2.680 ;
        RECT  0.520 0.920 0.680 2.680 ;
        RECT  0.370 0.920 0.520 1.080 ;
        RECT  0.210 2.520 0.520 2.680 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END NOR4BBX1TR

MACRO NOR4BXLTR
    CLASS CORE ;
    FOREIGN NOR4BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.640 2.720 2.760 ;
        RECT  2.480 0.920 2.640 2.760 ;
        RECT  2.250 0.920 2.480 1.080 ;
        RECT  2.200 2.470 2.480 2.760 ;
        RECT  1.970 0.540 2.250 1.080 ;
        RECT  1.320 0.920 1.970 1.080 ;
        RECT  1.040 0.540 1.320 1.080 ;
        END
        ANTENNADIFFAREA 3.04 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.640 1.120 1.990 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.760 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.420 1.960 1.600 ;
        RECT  1.680 1.420 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.280 2.800 0.280 ;
        RECT  2.430 -0.280 2.710 0.680 ;
        RECT  1.790 -0.280 2.430 0.280 ;
        RECT  1.510 -0.280 1.790 0.680 ;
        RECT  0.860 -0.280 1.510 0.280 ;
        RECT  0.580 -0.280 0.860 0.760 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 3.320 2.800 3.880 ;
        RECT  0.800 2.470 1.040 3.880 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.080 1.760 2.320 2.310 ;
        RECT  0.640 2.150 2.080 2.310 ;
        RECT  0.480 0.920 0.640 2.690 ;
        RECT  0.370 0.920 0.480 1.080 ;
        RECT  0.210 2.530 0.480 2.690 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END NOR4BXLTR

MACRO NOR4BX4TR
    CLASS CORE ;
    FOREIGN NOR4BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.580 0.440 7.820 3.060 ;
        RECT  7.280 0.440 7.580 1.360 ;
        RECT  6.120 2.820 7.580 3.060 ;
        RECT  1.050 0.460 7.280 0.700 ;
        RECT  5.840 2.820 6.120 3.100 ;
        RECT  2.400 2.820 5.840 3.060 ;
        RECT  2.120 2.820 2.400 3.100 ;
        END
        ANTENNADIFFAREA 9.771 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.200 1.760 7.420 2.660 ;
        RECT  4.390 2.500 7.200 2.660 ;
        RECT  4.110 2.140 4.390 2.660 ;
        RECT  1.560 2.440 4.110 2.660 ;
        RECT  1.480 2.440 1.560 2.760 ;
        RECT  1.240 2.140 1.480 2.760 ;
        RECT  1.160 2.140 1.240 2.300 ;
        RECT  1.000 1.560 1.160 2.300 ;
        RECT  0.880 1.560 1.000 1.800 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 1.280 7.120 1.560 ;
        RECT  6.880 1.280 7.040 2.340 ;
        RECT  5.200 2.180 6.880 2.340 ;
        RECT  5.040 1.520 5.200 2.340 ;
        RECT  4.840 1.520 5.040 1.980 ;
        RECT  3.320 1.820 4.840 1.980 ;
        RECT  3.040 1.700 3.320 1.980 ;
        RECT  1.480 1.820 3.040 1.980 ;
        RECT  1.320 1.180 1.480 1.980 ;
        RECT  1.190 1.180 1.320 1.400 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 1.740 6.720 2.020 ;
        RECT  5.880 1.740 6.440 1.900 ;
        RECT  5.760 1.520 5.880 1.900 ;
        RECT  5.600 1.200 5.760 1.900 ;
        RECT  2.880 1.200 5.600 1.360 ;
        RECT  2.650 1.200 2.880 1.660 ;
        RECT  1.960 1.500 2.650 1.660 ;
        RECT  1.640 1.240 1.960 1.660 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.380 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.050 -0.280 8.000 0.280 ;
        RECT  6.770 -0.280 7.050 0.300 ;
        RECT  6.010 -0.280 6.770 0.280 ;
        RECT  5.730 -0.280 6.010 0.300 ;
        RECT  4.970 -0.280 5.730 0.280 ;
        RECT  4.690 -0.280 4.970 0.300 ;
        RECT  3.930 -0.280 4.690 0.280 ;
        RECT  3.650 -0.280 3.930 0.300 ;
        RECT  2.890 -0.280 3.650 0.280 ;
        RECT  2.610 -0.280 2.890 0.300 ;
        RECT  1.850 -0.280 2.610 0.280 ;
        RECT  1.570 -0.280 1.850 0.300 ;
        RECT  0.850 -0.280 1.570 0.280 ;
        RECT  0.570 -0.280 0.850 0.660 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.720 3.320 8.000 3.880 ;
        RECT  7.440 3.220 7.720 3.880 ;
        RECT  3.960 3.320 7.440 3.880 ;
        RECT  3.680 3.220 3.960 3.880 ;
        RECT  0.850 3.320 3.680 3.880 ;
        RECT  0.570 2.460 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.480 1.300 6.650 1.580 ;
        RECT  6.320 0.860 6.480 1.580 ;
        RECT  2.490 0.860 6.320 1.020 ;
        RECT  2.210 0.860 2.490 1.280 ;
        RECT  0.370 0.860 2.210 1.020 ;
        RECT  0.240 0.500 0.370 1.220 ;
        RECT  0.240 2.190 0.370 3.080 ;
        RECT  0.080 0.500 0.240 3.080 ;
    END
END NOR4BX4TR

MACRO NOR4BX2TR
    CLASS CORE ;
    FOREIGN NOR4BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.600 0.820 4.720 2.760 ;
        RECT  4.560 0.820 4.600 3.040 ;
        RECT  4.240 0.820 4.560 0.980 ;
        RECT  4.440 1.640 4.560 3.040 ;
        RECT  2.520 2.880 4.440 3.040 ;
        RECT  3.960 0.700 4.240 0.980 ;
        RECT  3.320 0.700 3.960 0.860 ;
        RECT  3.040 0.700 3.320 0.980 ;
        RECT  2.380 0.700 3.040 0.930 ;
        RECT  2.240 2.880 2.520 3.160 ;
        RECT  1.060 0.650 2.380 0.930 ;
        END
        ANTENNADIFFAREA 5.328 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.240 3.960 1.920 ;
        RECT  3.680 1.240 3.840 2.400 ;
        RECT  1.280 2.240 3.680 2.400 ;
        RECT  1.120 1.750 1.280 2.400 ;
        RECT  1.000 1.750 1.120 2.030 ;
        END
        ANTENNAGATEAREA 0.3792 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.320 3.520 2.080 ;
        RECT  1.600 1.920 3.280 2.080 ;
        RECT  1.440 1.410 1.600 2.080 ;
        RECT  1.320 1.410 1.440 1.590 ;
        END
        ANTENNAGATEAREA 0.3792 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.240 3.120 1.760 ;
        RECT  2.100 1.600 2.760 1.760 ;
        RECT  1.820 1.410 2.100 1.760 ;
        END
        ANTENNAGATEAREA 0.3792 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.540 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.640 -0.280 4.800 0.280 ;
        RECT  4.360 -0.280 4.640 0.390 ;
        RECT  3.720 -0.280 4.360 0.280 ;
        RECT  3.440 -0.280 3.720 0.390 ;
        RECT  2.900 -0.280 3.440 0.280 ;
        RECT  2.620 -0.280 2.900 0.390 ;
        RECT  1.860 -0.280 2.620 0.280 ;
        RECT  1.580 -0.280 1.860 0.400 ;
        RECT  0.820 -0.280 1.580 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        RECT  0.000 -0.280 0.540 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.000 3.320 4.800 3.880 ;
        RECT  3.720 3.200 4.000 3.880 ;
        RECT  1.080 3.320 3.720 3.880 ;
        RECT  0.800 2.930 1.080 3.880 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.280 1.210 4.400 1.480 ;
        RECT  4.120 1.210 4.280 2.720 ;
        RECT  0.540 2.560 4.120 2.720 ;
        RECT  2.300 1.090 2.580 1.440 ;
        RECT  0.420 1.090 2.300 1.250 ;
        RECT  0.300 2.120 0.540 2.800 ;
        RECT  0.300 0.970 0.420 1.250 ;
        RECT  0.140 0.970 0.300 2.800 ;
    END
END NOR4BX2TR

MACRO NOR4BX1TR
    CLASS CORE ;
    FOREIGN NOR4BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.640 2.720 2.920 ;
        RECT  2.480 1.260 2.640 2.920 ;
        RECT  2.280 1.260 2.480 1.420 ;
        RECT  2.260 2.640 2.480 2.920 ;
        RECT  2.120 0.590 2.280 1.420 ;
        RECT  1.930 0.590 2.120 0.870 ;
        RECT  1.290 0.710 1.930 0.870 ;
        RECT  1.010 0.710 1.290 0.990 ;
        END
        ANTENNADIFFAREA 3.576 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.520 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.160 1.520 1.760 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.200 1.960 1.420 ;
        RECT  1.740 1.200 1.920 1.960 ;
        RECT  1.680 1.640 1.740 1.960 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.690 -0.280 2.800 0.280 ;
        RECT  2.440 -0.280 2.690 0.960 ;
        RECT  0.770 -0.280 2.440 0.280 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 3.320 2.800 3.880 ;
        RECT  0.760 2.840 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.080 1.580 2.300 2.280 ;
        RECT  1.880 2.120 2.080 2.280 ;
        RECT  1.720 2.120 1.880 2.680 ;
        RECT  0.680 2.490 1.720 2.680 ;
        RECT  0.520 0.920 0.680 2.680 ;
        RECT  0.370 0.920 0.520 1.080 ;
        RECT  0.210 2.520 0.520 2.680 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END NOR4BX1TR

MACRO NOR4XLTR
    CLASS CORE ;
    FOREIGN NOR4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 2.120 2.120 2.400 ;
        RECT  1.640 0.800 1.920 1.080 ;
        RECT  0.680 2.120 1.840 2.280 ;
        RECT  0.720 0.920 1.640 1.080 ;
        RECT  0.680 0.440 0.720 1.080 ;
        RECT  0.520 0.440 0.680 2.280 ;
        RECT  0.480 0.440 0.520 1.210 ;
        END
        ANTENNADIFFAREA 2.96 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.120 1.680 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.240 1.920 1.560 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.840 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 3.320 2.400 3.880 ;
        RECT  0.320 2.800 0.600 3.880 ;
        RECT  0.000 3.320 0.320 3.880 ;
        END
    END VDD
END NOR4XLTR

MACRO NOR4X8TR
    CLASS CORE ;
    FOREIGN NOR4X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.430 1.830 16.520 2.560 ;
        RECT  16.340 0.550 16.430 2.560 ;
        RECT  15.950 0.550 16.340 3.040 ;
        RECT  0.900 0.550 15.950 0.940 ;
        RECT  15.840 1.830 15.950 3.040 ;
        RECT  4.330 2.650 15.840 3.040 ;
        RECT  1.800 2.690 4.330 3.040 ;
        RECT  0.610 0.550 0.900 1.060 ;
        END
        ANTENNADIFFAREA 23.988 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.600 1.130 15.790 1.410 ;
        RECT  15.460 1.240 15.600 1.410 ;
        RECT  15.300 1.240 15.460 2.490 ;
        RECT  12.490 2.330 15.300 2.490 ;
        RECT  12.210 2.200 12.490 2.490 ;
        RECT  4.130 2.330 12.210 2.490 ;
        RECT  3.910 2.330 4.130 2.530 ;
        RECT  0.600 2.370 3.910 2.530 ;
        RECT  0.350 1.790 0.600 2.530 ;
        RECT  0.320 1.240 0.350 2.530 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 1.4016 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.960 1.120 15.140 2.010 ;
        RECT  14.800 1.120 14.960 1.360 ;
        RECT  13.520 1.850 14.960 2.010 ;
        RECT  13.180 1.850 13.520 2.070 ;
        RECT  11.460 1.850 13.180 2.010 ;
        RECT  11.440 1.850 11.460 2.100 ;
        RECT  11.190 1.790 11.440 2.100 ;
        RECT  9.330 1.940 11.190 2.100 ;
        RECT  9.050 1.790 9.330 2.100 ;
        RECT  7.330 1.940 9.050 2.100 ;
        RECT  7.040 1.780 7.330 2.100 ;
        RECT  5.210 1.940 7.040 2.100 ;
        RECT  4.930 1.790 5.210 2.100 ;
        RECT  3.130 1.940 4.930 2.100 ;
        RECT  3.090 1.790 3.130 2.100 ;
        RECT  2.890 1.790 3.090 2.210 ;
        RECT  1.120 2.050 2.890 2.210 ;
        RECT  0.930 1.440 1.120 2.210 ;
        RECT  0.810 1.440 0.930 1.960 ;
        END
        ANTENNAGATEAREA 1.4016 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.040 1.530 14.780 1.690 ;
        RECT  13.420 1.460 14.040 1.690 ;
        RECT  10.200 1.460 13.420 1.630 ;
        RECT  9.920 1.460 10.200 1.750 ;
        RECT  6.880 1.460 9.920 1.620 ;
        RECT  6.660 1.460 6.880 1.750 ;
        RECT  5.720 1.460 6.660 1.620 ;
        RECT  5.440 1.460 5.720 1.740 ;
        RECT  2.680 1.460 5.440 1.620 ;
        RECT  2.520 1.460 2.680 1.890 ;
        RECT  1.540 1.730 2.520 1.890 ;
        RECT  1.380 1.240 1.540 1.890 ;
        RECT  1.280 1.240 1.380 1.560 ;
        END
        ANTENNAGATEAREA 1.4016 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.330 1.110 14.390 1.270 ;
        RECT  14.110 1.100 14.330 1.270 ;
        RECT  2.320 1.100 14.110 1.260 ;
        RECT  2.080 1.100 2.320 1.560 ;
        RECT  1.870 1.100 2.080 1.370 ;
        END
        ANTENNAGATEAREA 1.4016 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.950 -0.280 16.800 0.280 ;
        RECT  15.670 -0.280 15.950 0.380 ;
        RECT  14.810 -0.280 15.670 0.280 ;
        RECT  14.530 -0.280 14.810 0.390 ;
        RECT  13.690 -0.280 14.530 0.280 ;
        RECT  13.410 -0.280 13.690 0.380 ;
        RECT  12.570 -0.280 13.410 0.280 ;
        RECT  12.290 -0.280 12.570 0.380 ;
        RECT  11.450 -0.280 12.290 0.280 ;
        RECT  11.170 -0.280 11.450 0.380 ;
        RECT  10.300 -0.280 11.170 0.280 ;
        RECT  10.020 -0.280 10.300 0.380 ;
        RECT  9.180 -0.280 10.020 0.280 ;
        RECT  8.900 -0.280 9.180 0.380 ;
        RECT  8.060 -0.280 8.900 0.280 ;
        RECT  7.780 -0.280 8.060 0.380 ;
        RECT  6.940 -0.280 7.780 0.280 ;
        RECT  6.660 -0.280 6.940 0.380 ;
        RECT  5.820 -0.280 6.660 0.280 ;
        RECT  5.540 -0.280 5.820 0.380 ;
        RECT  4.700 -0.280 5.540 0.280 ;
        RECT  4.420 -0.280 4.700 0.380 ;
        RECT  3.580 -0.280 4.420 0.280 ;
        RECT  3.300 -0.280 3.580 0.380 ;
        RECT  2.460 -0.280 3.300 0.280 ;
        RECT  2.180 -0.280 2.460 0.380 ;
        RECT  1.340 -0.280 2.180 0.280 ;
        RECT  1.060 -0.280 1.340 0.330 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 1.060 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.090 3.320 16.800 3.880 ;
        RECT  15.810 3.200 16.090 3.880 ;
        RECT  12.170 3.320 15.810 3.880 ;
        RECT  11.890 3.200 12.170 3.880 ;
        RECT  7.990 3.320 11.890 3.880 ;
        RECT  7.730 3.200 7.990 3.880 ;
        RECT  3.840 3.320 7.730 3.880 ;
        RECT  3.560 3.200 3.840 3.880 ;
        RECT  0.580 3.320 3.560 3.880 ;
        RECT  0.300 2.810 0.580 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
END NOR4X8TR

MACRO NOR4X6TR
    CLASS CORE ;
    FOREIGN NOR4X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.180 0.460 11.520 2.940 ;
        RECT  10.680 0.460 11.180 1.360 ;
        RECT  9.840 2.580 11.180 2.940 ;
        RECT  2.480 0.460 10.680 0.820 ;
        RECT  9.560 2.580 9.840 3.140 ;
        RECT  6.120 2.580 9.560 2.940 ;
        RECT  5.840 2.580 6.120 3.140 ;
        RECT  2.290 2.580 5.840 2.940 ;
        RECT  0.840 0.460 2.480 0.680 ;
        RECT  1.980 2.580 2.290 3.140 ;
        RECT  0.590 0.460 0.840 1.140 ;
        END
        ANTENNADIFFAREA 15.032 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.860 1.860 11.020 2.420 ;
        RECT  8.070 2.250 10.860 2.420 ;
        RECT  7.690 2.140 8.070 2.420 ;
        RECT  4.160 2.250 7.690 2.420 ;
        RECT  3.880 2.140 4.160 2.420 ;
        RECT  0.720 2.260 3.880 2.420 ;
        RECT  0.480 1.840 0.720 2.420 ;
        END
        ANTENNAGATEAREA 1.0488 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.640 1.540 10.760 1.700 ;
        RECT  10.480 1.540 10.640 1.980 ;
        RECT  8.920 1.820 10.480 1.980 ;
        RECT  8.640 1.700 8.920 1.980 ;
        RECT  7.040 1.820 8.640 1.980 ;
        RECT  6.760 1.700 7.040 1.980 ;
        RECT  5.200 1.820 6.760 1.980 ;
        RECT  4.920 1.700 5.200 1.980 ;
        RECT  3.240 1.820 4.920 1.980 ;
        RECT  3.120 1.700 3.240 1.980 ;
        RECT  2.960 1.700 3.120 2.100 ;
        RECT  1.120 1.940 2.960 2.100 ;
        RECT  0.880 1.330 1.120 2.100 ;
        END
        ANTENNAGATEAREA 1.0488 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.160 1.000 10.320 1.540 ;
        RECT  9.600 1.380 10.160 1.540 ;
        RECT  9.320 1.380 9.600 1.660 ;
        RECT  6.600 1.380 9.320 1.540 ;
        RECT  6.320 1.380 6.600 1.660 ;
        RECT  5.640 1.380 6.320 1.540 ;
        RECT  5.360 1.380 5.640 1.660 ;
        RECT  2.800 1.380 5.360 1.540 ;
        RECT  2.520 1.380 2.800 1.780 ;
        RECT  1.620 1.620 2.520 1.780 ;
        RECT  1.280 1.240 1.620 1.780 ;
        END
        ANTENNAGATEAREA 1.0488 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.640 1.000 9.920 1.220 ;
        RECT  6.240 1.060 9.640 1.220 ;
        RECT  2.320 1.000 6.240 1.220 ;
        RECT  2.160 0.840 2.320 1.220 ;
        RECT  1.880 0.840 2.160 1.460 ;
        END
        ANTENNAGATEAREA 1.0488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.720 -0.280 11.600 0.280 ;
        RECT  10.440 -0.280 10.720 0.300 ;
        RECT  9.680 -0.280 10.440 0.280 ;
        RECT  9.400 -0.280 9.680 0.300 ;
        RECT  8.640 -0.280 9.400 0.280 ;
        RECT  8.360 -0.280 8.640 0.300 ;
        RECT  7.600 -0.280 8.360 0.280 ;
        RECT  7.320 -0.280 7.600 0.300 ;
        RECT  6.560 -0.280 7.320 0.280 ;
        RECT  6.280 -0.280 6.560 0.300 ;
        RECT  5.520 -0.280 6.280 0.280 ;
        RECT  5.240 -0.280 5.520 0.300 ;
        RECT  4.480 -0.280 5.240 0.280 ;
        RECT  4.200 -0.280 4.480 0.300 ;
        RECT  3.440 -0.280 4.200 0.280 ;
        RECT  3.160 -0.280 3.440 0.300 ;
        RECT  2.400 -0.280 3.160 0.280 ;
        RECT  2.120 -0.280 2.400 0.300 ;
        RECT  0.380 -0.280 2.120 0.280 ;
        RECT  0.090 -0.280 0.380 1.090 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.320 3.320 11.600 3.880 ;
        RECT  11.040 3.200 11.320 3.880 ;
        RECT  7.680 3.320 11.040 3.880 ;
        RECT  7.400 3.200 7.680 3.880 ;
        RECT  3.880 3.320 7.400 3.880 ;
        RECT  3.600 3.200 3.880 3.880 ;
        RECT  0.720 3.320 3.600 3.880 ;
        RECT  0.440 2.800 0.720 3.880 ;
        RECT  0.000 3.320 0.440 3.880 ;
        END
    END VDD
END NOR4X6TR

MACRO NOR4X4TR
    CLASS CORE ;
    FOREIGN NOR4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.320 1.020 7.520 3.070 ;
        RECT  7.120 1.020 7.320 1.360 ;
        RECT  1.810 2.830 7.320 3.070 ;
        RECT  6.880 0.520 7.120 1.360 ;
        RECT  6.000 0.520 6.880 0.760 ;
        RECT  5.720 0.480 6.000 0.760 ;
        RECT  4.960 0.520 5.720 0.760 ;
        RECT  4.680 0.480 4.960 0.760 ;
        RECT  3.920 0.520 4.680 0.760 ;
        RECT  3.640 0.480 3.920 0.760 ;
        RECT  1.720 0.510 3.640 0.760 ;
        RECT  1.440 0.480 1.720 0.760 ;
        RECT  0.800 0.520 1.440 0.760 ;
        RECT  0.520 0.520 0.800 0.930 ;
        END
        ANTENNADIFFAREA 11.298 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.820 7.160 2.670 ;
        RECT  4.120 2.510 7.000 2.670 ;
        RECT  3.840 2.000 4.120 2.670 ;
        RECT  0.720 2.460 3.840 2.620 ;
        RECT  0.650 2.000 0.720 2.620 ;
        RECT  0.530 1.720 0.650 2.620 ;
        RECT  0.480 1.720 0.530 2.360 ;
        RECT  0.330 1.720 0.480 1.980 ;
        END
        ANTENNAGATEAREA 0.72 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.720 1.530 6.840 2.350 ;
        RECT  6.680 1.360 6.720 2.350 ;
        RECT  6.560 1.360 6.680 1.690 ;
        RECT  4.980 2.190 6.680 2.350 ;
        RECT  4.820 1.560 4.980 2.350 ;
        RECT  4.700 1.560 4.820 1.840 ;
        RECT  3.120 1.680 4.700 1.840 ;
        RECT  2.960 1.680 3.120 2.300 ;
        RECT  1.120 2.140 2.960 2.300 ;
        RECT  0.930 1.240 1.120 2.300 ;
        RECT  0.850 1.240 0.930 1.660 ;
        END
        ANTENNAGATEAREA 0.72 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.210 1.810 6.440 2.030 ;
        RECT  5.420 1.870 6.210 2.030 ;
        RECT  5.260 1.240 5.420 2.030 ;
        RECT  2.740 1.240 5.260 1.400 ;
        RECT  2.570 1.240 2.740 1.980 ;
        RECT  1.520 1.820 2.570 1.980 ;
        RECT  1.280 1.300 1.520 1.980 ;
        END
        ANTENNAGATEAREA 0.72 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.070 6.200 1.350 ;
        RECT  5.920 0.920 6.080 1.350 ;
        RECT  2.320 0.920 5.920 1.080 ;
        RECT  2.080 0.920 2.320 1.660 ;
        RECT  1.730 1.380 2.080 1.660 ;
        END
        ANTENNAGATEAREA 0.72 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.520 -0.280 7.600 0.280 ;
        RECT  6.240 -0.280 6.520 0.360 ;
        RECT  5.480 -0.280 6.240 0.280 ;
        RECT  5.200 -0.280 5.480 0.360 ;
        RECT  4.440 -0.280 5.200 0.280 ;
        RECT  4.160 -0.280 4.440 0.360 ;
        RECT  3.400 -0.280 4.160 0.280 ;
        RECT  3.120 -0.280 3.400 0.340 ;
        RECT  2.240 -0.280 3.120 0.280 ;
        RECT  1.960 -0.280 2.240 0.340 ;
        RECT  0.000 -0.280 1.960 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.500 3.320 7.600 3.880 ;
        RECT  7.220 3.230 7.500 3.880 ;
        RECT  3.880 3.260 7.220 3.880 ;
        RECT  3.600 3.230 3.880 3.880 ;
        RECT  0.530 3.320 3.600 3.880 ;
        RECT  0.250 2.780 0.530 3.880 ;
        RECT  0.000 3.320 0.250 3.880 ;
        END
    END VDD
END NOR4X4TR

MACRO NOR4X2TR
    CLASS CORE ;
    FOREIGN NOR4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 0.720 3.760 1.000 ;
        RECT  2.800 0.840 3.480 1.000 ;
        RECT  2.520 0.720 2.800 1.000 ;
        RECT  1.760 0.840 2.520 1.000 ;
        RECT  0.240 2.680 2.260 2.960 ;
        RECT  1.480 0.720 1.760 1.000 ;
        RECT  0.840 0.840 1.480 1.000 ;
        RECT  0.240 0.840 0.840 1.160 ;
        RECT  0.080 0.840 0.240 2.960 ;
        END
        ANTENNADIFFAREA 6.432 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.640 3.960 1.960 ;
        RECT  3.680 1.640 3.840 2.520 ;
        RECT  0.680 2.360 3.680 2.520 ;
        RECT  0.400 1.640 0.680 2.520 ;
        END
        ANTENNAGATEAREA 0.3984 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 1.240 3.520 1.640 ;
        RECT  3.200 1.240 3.360 2.200 ;
        RECT  1.120 2.040 3.200 2.200 ;
        RECT  0.960 1.320 1.120 2.200 ;
        RECT  0.840 1.320 0.960 1.600 ;
        END
        ANTENNAGATEAREA 0.3984 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.600 2.840 1.880 ;
        RECT  1.560 1.720 2.560 1.880 ;
        RECT  1.400 1.240 1.560 1.880 ;
        RECT  1.280 1.240 1.400 1.560 ;
        END
        ANTENNAGATEAREA 0.3984 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.240 2.380 1.560 ;
        END
        ANTENNAGATEAREA 0.3984 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 -0.280 4.400 0.280 ;
        RECT  3.950 -0.280 4.240 1.060 ;
        RECT  3.320 -0.280 3.950 0.280 ;
        RECT  3.040 -0.280 3.320 0.400 ;
        RECT  2.280 -0.280 3.040 0.280 ;
        RECT  2.000 -0.280 2.280 0.400 ;
        RECT  0.160 -0.280 2.000 0.340 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.800 3.320 4.400 3.880 ;
        RECT  3.520 2.800 3.800 3.880 ;
        RECT  0.600 3.320 3.520 3.880 ;
        RECT  0.320 3.200 0.600 3.880 ;
        RECT  0.000 3.320 0.320 3.880 ;
        END
    END VDD
END NOR4X2TR

MACRO NOR4X1TR
    CLASS CORE ;
    FOREIGN NOR4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.840 2.720 2.080 ;
        RECT  2.180 0.840 2.480 1.000 ;
        RECT  2.370 1.920 2.480 2.080 ;
        RECT  2.090 1.920 2.370 3.080 ;
        RECT  1.900 0.720 2.180 1.000 ;
        RECT  1.140 0.840 1.900 1.000 ;
        RECT  0.860 0.720 1.140 1.000 ;
        END
        ANTENNADIFFAREA 3.576 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.240 0.720 1.950 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.160 1.390 1.480 ;
        RECT  0.880 1.160 1.130 1.970 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.160 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.760 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 -0.280 2.800 0.280 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  1.660 -0.280 2.420 0.280 ;
        RECT  1.380 -0.280 1.660 0.400 ;
        RECT  0.660 -0.280 1.380 0.280 ;
        RECT  0.380 -0.280 0.660 0.930 ;
        RECT  0.000 -0.280 0.380 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.890 3.320 2.800 3.880 ;
        RECT  0.610 2.420 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
END NOR4X1TR

MACRO NOR3BXLTR
    CLASS CORE ;
    FOREIGN NOR3BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.440 2.320 1.560 ;
        RECT  2.080 0.440 2.210 2.350 ;
        RECT  1.930 0.520 2.080 2.350 ;
        RECT  1.130 0.520 1.930 0.760 ;
        END
        ANTENNADIFFAREA 2.4295 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.360 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.600 1.680 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.280 2.400 0.280 ;
        RECT  0.670 -0.280 0.940 0.750 ;
        RECT  0.000 -0.280 0.670 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 3.320 2.400 3.880 ;
        RECT  0.770 2.840 1.050 3.880 ;
        RECT  0.000 3.320 0.770 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.370 2.660 2.010 2.940 ;
        RECT  1.210 2.520 1.370 2.940 ;
        RECT  0.640 2.520 1.210 2.680 ;
        RECT  0.480 0.920 0.640 2.680 ;
        RECT  0.090 0.920 0.480 1.080 ;
        RECT  0.370 2.520 0.480 2.680 ;
        RECT  0.090 2.520 0.370 2.800 ;
    END
END NOR3BXLTR

MACRO NOR3BX4TR
    CLASS CORE ;
    FOREIGN NOR3BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.310 0.640 5.550 2.760 ;
        RECT  5.280 0.640 5.310 1.360 ;
        RECT  4.290 2.520 5.310 2.760 ;
        RECT  4.250 0.970 5.280 1.210 ;
        RECT  4.010 2.440 4.290 3.040 ;
        RECT  3.970 0.440 4.250 1.210 ;
        RECT  2.050 2.440 4.010 2.680 ;
        RECT  3.170 0.560 3.970 0.800 ;
        RECT  2.890 0.440 3.170 0.800 ;
        RECT  2.130 0.560 2.890 0.800 ;
        RECT  1.850 0.560 2.130 0.840 ;
        RECT  1.770 2.440 2.050 3.040 ;
        END
        ANTENNADIFFAREA 8.47 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.710 5.150 2.360 ;
        RECT  4.880 2.040 4.990 2.360 ;
        RECT  3.170 2.120 4.880 2.280 ;
        RECT  2.890 1.700 3.170 2.280 ;
        RECT  1.250 2.120 2.890 2.280 ;
        RECT  0.850 2.060 1.250 2.280 ;
        END
        ANTENNAGATEAREA 0.6432 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.370 5.100 1.530 ;
        RECT  3.810 1.370 3.930 1.640 ;
        RECT  3.650 1.060 3.810 1.640 ;
        RECT  2.410 1.060 3.650 1.220 ;
        RECT  2.250 1.060 2.410 1.640 ;
        RECT  2.130 1.200 2.250 1.640 ;
        RECT  1.520 1.200 2.130 1.360 ;
        RECT  1.170 0.840 1.520 1.360 ;
        END
        ANTENNAGATEAREA 0.6432 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.800 1.580 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.770 -0.280 6.000 0.280 ;
        RECT  4.490 -0.280 4.770 0.810 ;
        RECT  3.690 -0.280 4.490 0.280 ;
        RECT  3.410 -0.280 3.690 0.400 ;
        RECT  2.650 -0.280 3.410 0.280 ;
        RECT  2.370 -0.280 2.650 0.400 ;
        RECT  1.650 -0.280 2.370 0.280 ;
        RECT  0.930 -0.280 1.650 0.680 ;
        RECT  0.650 -0.280 0.930 1.080 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 3.320 6.000 3.880 ;
        RECT  5.340 2.920 5.620 3.880 ;
        RECT  3.170 3.320 5.340 3.880 ;
        RECT  2.890 2.840 3.170 3.880 ;
        RECT  0.930 3.320 2.890 3.880 ;
        RECT  0.650 2.530 0.930 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.170 1.690 4.450 1.960 ;
        RECT  3.490 1.800 4.170 1.960 ;
        RECT  3.330 1.380 3.490 1.960 ;
        RECT  2.730 1.380 3.330 1.540 ;
        RECT  2.570 1.380 2.730 1.960 ;
        RECT  1.850 1.800 2.570 1.960 ;
        RECT  1.570 1.740 1.850 1.960 ;
        RECT  0.320 1.740 1.570 1.900 ;
        RECT  0.320 0.800 0.490 1.080 ;
        RECT  0.320 2.170 0.450 2.970 ;
        RECT  0.160 0.800 0.320 2.970 ;
    END
END NOR3BX4TR

MACRO NOR3BX2TR
    CLASS CORE ;
    FOREIGN NOR3BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 0.440 1.810 1.060 ;
        RECT  0.850 0.900 1.520 1.060 ;
        RECT  1.280 2.670 1.520 3.160 ;
        RECT  0.240 2.670 1.280 2.830 ;
        RECT  0.570 0.440 0.850 1.060 ;
        RECT  0.240 0.900 0.570 1.060 ;
        RECT  0.080 0.900 0.240 2.830 ;
        END
        ANTENNADIFFAREA 5 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.580 2.460 1.860 ;
        RECT  2.180 1.580 2.340 2.510 ;
        RECT  0.720 2.350 2.180 2.510 ;
        RECT  0.560 2.040 0.720 2.510 ;
        RECT  0.400 1.840 0.560 2.510 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.590 1.930 1.750 ;
        RECT  1.650 1.590 1.810 2.180 ;
        RECT  1.040 2.020 1.650 2.180 ;
        RECT  1.040 1.240 1.120 1.580 ;
        RECT  0.880 1.240 1.040 2.180 ;
        RECT  0.690 1.240 0.880 1.580 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.440 2.760 0.760 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 -0.280 3.200 0.280 ;
        RECT  2.160 -0.280 2.320 0.820 ;
        RECT  1.330 -0.280 2.160 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.870 3.320 3.200 3.880 ;
        RECT  2.590 2.920 2.870 3.880 ;
        RECT  0.370 3.320 2.590 3.880 ;
        RECT  0.090 2.990 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.830 0.920 3.110 2.380 ;
        RECT  1.440 1.260 2.830 1.420 ;
        RECT  1.280 1.260 1.440 1.640 ;
    END
END NOR3BX2TR

MACRO NOR3BX1TR
    CLASS CORE ;
    FOREIGN NOR3BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.440 2.320 2.720 ;
        RECT  2.080 0.440 2.160 1.560 ;
        RECT  1.760 2.440 2.160 2.720 ;
        RECT  1.390 0.900 2.080 1.060 ;
        RECT  1.110 0.780 1.390 1.060 ;
        END
        ANTENNADIFFAREA 3.196 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.220 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.220 1.560 1.570 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.240 0.720 1.560 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 -0.280 2.400 0.280 ;
        RECT  0.590 -0.280 1.790 0.340 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 3.320 2.400 3.880 ;
        RECT  0.600 2.800 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.880 1.580 1.920 1.860 ;
        RECT  1.720 1.580 1.880 2.280 ;
        RECT  0.370 2.120 1.720 2.280 ;
        RECT  0.240 0.800 0.370 1.080 ;
        RECT  0.240 1.920 0.370 2.280 ;
        RECT  0.080 0.800 0.240 2.280 ;
    END
END NOR3BX1TR

MACRO NOR3XLTR
    CLASS CORE ;
    FOREIGN NOR3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.910 1.920 2.360 ;
        RECT  1.680 0.910 1.740 2.680 ;
        RECT  0.900 0.910 1.680 1.070 ;
        RECT  1.460 2.040 1.680 2.680 ;
        RECT  0.590 0.910 0.900 1.260 ;
        END
        ANTENNADIFFAREA 2.048 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.540 0.660 1.790 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.520 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.230 1.520 1.800 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.090 -0.280 1.360 0.550 ;
        RECT  0.410 -0.280 1.090 0.280 ;
        RECT  0.130 -0.280 0.410 0.670 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 3.320 2.000 3.880 ;
        RECT  0.300 2.190 0.590 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
END NOR3XLTR

MACRO NOR3X8TR
    CLASS CORE ;
    FOREIGN NOR3X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.230 0.440 8.710 2.860 ;
        RECT  6.090 0.440 8.230 0.850 ;
        RECT  7.880 1.830 8.230 2.860 ;
        RECT  6.210 2.380 7.880 2.860 ;
        RECT  5.930 2.380 6.210 3.160 ;
        RECT  1.090 0.450 6.090 0.670 ;
        RECT  3.890 2.380 5.930 2.860 ;
        RECT  3.610 2.380 3.890 3.160 ;
        RECT  1.570 2.380 3.610 2.860 ;
        RECT  1.290 2.380 1.570 3.160 ;
        RECT  0.810 0.450 1.090 1.150 ;
        END
        ANTENNADIFFAREA 18.1165 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.970 1.650 7.240 2.220 ;
        RECT  5.130 2.060 6.970 2.220 ;
        RECT  4.850 1.590 5.130 2.220 ;
        RECT  2.490 2.030 4.850 2.220 ;
        RECT  2.210 1.590 2.490 2.220 ;
        RECT  0.530 2.050 2.210 2.220 ;
        RECT  0.320 1.590 0.530 2.220 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 1.3632 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.330 7.690 1.490 ;
        RECT  6.650 1.330 6.810 1.900 ;
        RECT  6.530 1.590 6.650 1.900 ;
        RECT  5.470 1.740 6.530 1.900 ;
        RECT  5.310 1.150 5.470 1.900 ;
        RECT  4.410 1.150 5.310 1.430 ;
        RECT  4.250 1.150 4.410 1.610 ;
        RECT  3.130 1.450 4.250 1.610 ;
        RECT  2.970 1.150 3.130 1.610 ;
        RECT  1.960 1.150 2.970 1.430 ;
        RECT  1.640 1.150 1.960 1.870 ;
        RECT  0.970 1.710 1.640 1.870 ;
        RECT  0.690 1.590 0.970 1.870 ;
        END
        ANTENNAGATEAREA 1.3632 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.910 1.010 8.070 1.640 ;
        RECT  6.170 1.010 7.910 1.170 ;
        RECT  5.920 1.010 6.170 1.580 ;
        RECT  5.890 0.830 5.920 1.580 ;
        RECT  5.680 0.830 5.890 1.170 ;
        RECT  4.090 0.830 5.680 0.990 ;
        RECT  3.410 0.830 4.090 1.290 ;
        RECT  1.410 0.830 3.410 0.990 ;
        RECT  1.250 0.830 1.410 1.550 ;
        RECT  1.130 1.330 1.250 1.550 ;
        END
        ANTENNAGATEAREA 1.3632 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.930 -0.280 8.800 0.280 ;
        RECT  5.650 -0.280 5.930 0.290 ;
        RECT  4.890 -0.280 5.650 0.280 ;
        RECT  4.610 -0.280 4.890 0.290 ;
        RECT  3.850 -0.280 4.610 0.280 ;
        RECT  3.570 -0.280 3.850 0.290 ;
        RECT  1.610 -0.280 3.570 0.280 ;
        RECT  1.330 -0.280 1.610 0.290 ;
        RECT  0.610 -0.280 1.330 0.280 ;
        RECT  0.330 -0.280 0.610 0.800 ;
        RECT  0.000 -0.280 0.330 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.450 3.320 8.800 3.880 ;
        RECT  7.170 3.180 7.450 3.880 ;
        RECT  5.050 3.320 7.170 3.880 ;
        RECT  4.770 3.180 5.050 3.880 ;
        RECT  2.730 3.320 4.770 3.880 ;
        RECT  2.450 3.180 2.730 3.880 ;
        RECT  0.370 3.320 2.450 3.880 ;
        RECT  0.090 2.590 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END NOR3X8TR

MACRO NOR3X6TR
    CLASS CORE ;
    FOREIGN NOR3X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 0.440 7.120 2.960 ;
        RECT  6.300 0.440 6.760 0.930 ;
        RECT  6.260 2.240 6.760 2.960 ;
        RECT  1.200 0.440 6.300 0.760 ;
        RECT  5.980 2.240 6.260 3.100 ;
        RECT  4.020 2.240 5.980 2.600 ;
        RECT  3.740 2.240 4.020 3.160 ;
        RECT  1.700 2.400 3.740 2.760 ;
        RECT  1.420 2.400 1.700 3.160 ;
        RECT  0.920 0.440 1.200 0.980 ;
        END
        ANTENNADIFFAREA 14.002 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.260 1.850 6.590 2.080 ;
        RECT  5.330 1.920 6.260 2.080 ;
        RECT  4.660 1.640 5.330 2.080 ;
        RECT  2.620 1.920 4.660 2.080 ;
        RECT  2.500 1.640 2.620 2.080 ;
        RECT  2.340 1.640 2.500 2.240 ;
        RECT  0.720 2.080 2.340 2.240 ;
        RECT  0.560 1.240 0.720 2.240 ;
        RECT  0.420 1.240 0.560 1.600 ;
        END
        ANTENNAGATEAREA 1.0752 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.140 1.260 5.740 1.420 ;
        RECT  3.980 1.260 4.140 1.760 ;
        RECT  3.260 1.600 3.980 1.760 ;
        RECT  3.100 1.240 3.260 1.760 ;
        RECT  1.920 1.240 3.100 1.460 ;
        RECT  1.680 1.240 1.920 1.920 ;
        RECT  1.040 1.760 1.680 1.920 ;
        RECT  0.880 1.640 1.040 1.920 ;
        END
        ANTENNAGATEAREA 1.0752 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.140 1.240 6.320 1.580 ;
        RECT  5.980 0.920 6.140 1.580 ;
        RECT  3.820 0.920 5.980 1.080 ;
        RECT  3.540 0.920 3.820 1.440 ;
        RECT  1.520 0.920 3.540 1.080 ;
        RECT  1.360 0.920 1.520 1.600 ;
        RECT  1.220 1.320 1.360 1.600 ;
        END
        ANTENNAGATEAREA 1.0752 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.280 7.200 0.280 ;
        RECT  0.440 -0.280 0.720 0.870 ;
        RECT  0.000 -0.280 0.440 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.140 3.320 7.200 3.880 ;
        RECT  4.860 2.930 5.140 3.880 ;
        RECT  2.820 3.320 4.860 3.880 ;
        RECT  2.540 2.930 2.820 3.880 ;
        RECT  0.500 3.320 2.540 3.880 ;
        RECT  0.220 2.400 0.500 3.880 ;
        RECT  0.000 3.320 0.220 3.880 ;
        END
    END VDD
END NOR3X6TR

MACRO NOR3X4TR
    CLASS CORE ;
    FOREIGN NOR3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.130 5.120 2.760 ;
        RECT  4.720 1.130 4.880 1.370 ;
        RECT  3.860 2.520 4.880 2.760 ;
        RECT  4.480 0.600 4.720 1.370 ;
        RECT  3.780 0.600 4.480 0.840 ;
        RECT  3.580 2.440 3.860 2.760 ;
        RECT  3.770 0.440 3.780 0.840 ;
        RECT  3.520 0.440 3.770 1.060 ;
        RECT  1.620 2.440 3.580 2.660 ;
        RECT  3.500 0.440 3.520 0.840 ;
        RECT  1.400 0.560 3.500 0.840 ;
        RECT  1.340 2.440 1.620 2.720 ;
        END
        ANTENNADIFFAREA 8.496 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.560 1.720 4.720 2.280 ;
        RECT  4.320 2.120 4.560 2.280 ;
        RECT  4.080 2.040 4.320 2.360 ;
        RECT  2.720 2.120 4.080 2.280 ;
        RECT  2.440 1.720 2.720 2.280 ;
        RECT  0.740 2.120 2.440 2.280 ;
        RECT  0.580 1.680 0.740 2.280 ;
        RECT  0.340 1.680 0.580 1.850 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.220 4.320 1.700 ;
        RECT  3.480 1.220 4.160 1.400 ;
        RECT  3.360 1.220 3.480 1.640 ;
        RECT  3.200 1.080 3.360 1.640 ;
        RECT  1.960 1.080 3.200 1.240 ;
        RECT  1.680 1.080 1.960 1.640 ;
        RECT  0.890 1.080 1.680 1.240 ;
        RECT  0.600 0.840 0.890 1.460 ;
        RECT  0.480 0.840 0.600 1.160 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.640 3.920 1.960 ;
        RECT  3.040 1.800 3.680 1.960 ;
        RECT  2.880 1.400 3.040 1.960 ;
        RECT  2.280 1.400 2.880 1.560 ;
        RECT  2.120 1.400 2.280 1.960 ;
        RECT  1.420 1.800 2.120 1.960 ;
        RECT  1.140 1.680 1.420 1.960 ;
        END
        ANTENNAGATEAREA 0.6912 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.320 -0.280 5.200 0.280 ;
        RECT  4.040 -0.280 4.320 0.400 ;
        RECT  3.260 -0.280 4.040 0.280 ;
        RECT  2.980 -0.280 3.260 0.400 ;
        RECT  2.200 -0.280 2.980 0.280 ;
        RECT  1.920 -0.280 2.200 0.400 ;
        RECT  1.200 -0.280 1.920 0.280 ;
        RECT  0.920 -0.280 1.200 0.670 ;
        RECT  0.000 -0.280 0.920 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.020 3.320 5.200 3.880 ;
        RECT  4.740 3.010 5.020 3.880 ;
        RECT  2.740 3.320 4.740 3.880 ;
        RECT  2.460 2.820 2.740 3.880 ;
        RECT  0.420 3.260 2.460 3.880 ;
        RECT  0.140 2.120 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
END NOR3X4TR

MACRO NOR3X2TR
    CLASS CORE ;
    FOREIGN NOR3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.840 2.360 1.160 ;
        RECT  1.890 0.840 1.970 2.280 ;
        RECT  1.810 0.800 1.890 2.280 ;
        RECT  1.610 0.800 1.810 1.080 ;
        RECT  1.490 2.120 1.810 2.280 ;
        RECT  0.850 0.920 1.610 1.080 ;
        RECT  1.210 2.120 1.490 2.400 ;
        RECT  0.570 0.440 0.850 1.080 ;
        END
        ANTENNADIFFAREA 4.548 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.620 2.410 1.900 ;
        RECT  2.130 1.620 2.290 2.720 ;
        RECT  0.690 2.560 2.130 2.720 ;
        RECT  0.690 1.240 0.720 1.560 ;
        RECT  0.530 1.240 0.690 2.720 ;
        RECT  0.350 1.240 0.530 1.560 ;
        END
        ANTENNAGATEAREA 0.3264 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.280 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.3264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.640 1.820 ;
        END
        ANTENNAGATEAREA 0.3264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.280 2.800 0.280 ;
        RECT  1.090 -0.280 1.370 0.400 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.450 2.110 2.710 3.880 ;
        RECT  0.370 3.260 2.450 3.880 ;
        RECT  0.090 1.970 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END NOR3X2TR

MACRO NOR3X1TR
    CLASS CORE ;
    FOREIGN NOR3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.910 1.920 2.360 ;
        RECT  1.680 0.910 1.740 2.980 ;
        RECT  0.950 0.910 1.680 1.070 ;
        RECT  1.460 2.040 1.680 2.980 ;
        RECT  0.660 0.910 0.950 1.260 ;
        END
        ANTENNADIFFAREA 3.196 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.540 0.660 1.790 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.520 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.230 1.520 1.800 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.090 -0.280 1.360 0.550 ;
        RECT  0.410 -0.280 1.090 0.280 ;
        RECT  0.130 -0.280 0.410 0.680 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 3.320 2.000 3.880 ;
        RECT  0.300 2.190 0.590 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
END NOR3X1TR

MACRO NOR2BXLTR
    CLASS CORE ;
    FOREIGN NOR2BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.790 1.920 3.160 ;
        RECT  1.220 0.790 1.760 1.090 ;
        RECT  1.600 1.940 1.760 3.160 ;
        END
        ANTENNADIFFAREA 1.492 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.610 1.120 2.070 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.240 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.280 2.000 0.280 ;
        RECT  0.720 -0.280 1.880 0.340 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 3.320 2.000 3.880 ;
        RECT  0.680 2.560 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.360 1.600 1.640 ;
        RECT  1.280 1.290 1.440 2.400 ;
        RECT  1.040 1.290 1.280 1.450 ;
        RECT  0.380 2.240 1.280 2.400 ;
        RECT  0.880 0.910 1.040 1.450 ;
        RECT  0.370 0.910 0.880 1.080 ;
        RECT  0.090 1.940 0.380 2.400 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END NOR2BXLTR

MACRO NOR2BX4TR
    CLASS CORE ;
    FOREIGN NOR2BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.060 3.440 3.010 ;
        RECT  2.320 1.060 3.200 1.220 ;
        RECT  3.090 1.840 3.200 3.010 ;
        RECT  2.880 1.840 3.090 2.560 ;
        RECT  1.760 2.140 2.880 2.300 ;
        RECT  2.070 0.440 2.320 1.220 ;
        RECT  2.040 0.440 2.070 1.100 ;
        RECT  1.360 0.940 2.040 1.100 ;
        RECT  1.480 2.140 1.760 2.950 ;
        RECT  1.080 0.440 1.360 1.100 ;
        END
        ANTENNADIFFAREA 6.981 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.700 2.400 1.980 ;
        RECT  1.520 1.820 2.120 1.980 ;
        RECT  1.130 1.640 1.520 1.980 ;
        RECT  0.880 1.580 1.130 1.980 ;
        END
        ANTENNAGATEAREA 0.5952 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2472 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.020 -0.280 3.600 0.280 ;
        RECT  3.020 0.570 3.240 0.840 ;
        RECT  2.740 -0.280 3.020 0.840 ;
        RECT  1.840 -0.280 2.740 0.280 ;
        RECT  2.560 0.570 2.740 0.840 ;
        RECT  1.560 -0.280 1.840 0.670 ;
        RECT  0.880 -0.280 1.560 0.280 ;
        RECT  0.600 -0.280 0.880 1.100 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 3.320 3.600 3.880 ;
        RECT  2.280 2.460 2.560 3.880 ;
        RECT  0.960 3.260 2.280 3.880 ;
        RECT  0.680 2.140 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.760 1.380 3.040 1.660 ;
        RECT  1.900 1.380 2.760 1.540 ;
        RECT  1.890 1.260 1.900 1.540 ;
        RECT  1.730 1.260 1.890 1.660 ;
        RECT  0.400 1.260 1.730 1.420 ;
        RECT  0.240 2.120 0.480 2.920 ;
        RECT  0.240 0.500 0.400 1.420 ;
        RECT  0.200 0.500 0.240 2.920 ;
        RECT  0.080 0.500 0.200 2.280 ;
    END
END NOR2BX4TR

MACRO NOR2BX2TR
    CLASS CORE ;
    FOREIGN NOR2BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.110 2.400 2.030 ;
        RECT  1.880 1.110 2.240 1.270 ;
        RECT  1.920 1.870 2.240 2.030 ;
        RECT  1.760 1.870 1.920 2.720 ;
        RECT  1.600 0.440 1.880 1.270 ;
        RECT  1.720 2.440 1.760 2.720 ;
        RECT  1.240 2.440 1.720 2.760 ;
        END
        ANTENNADIFFAREA 3.168 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.430 2.080 1.710 ;
        RECT  1.160 1.430 1.800 1.590 ;
        RECT  1.000 1.430 1.160 1.960 ;
        RECT  0.840 1.640 1.000 1.960 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.440 0.320 1.640 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.280 2.800 0.280 ;
        RECT  2.120 -0.280 2.400 0.950 ;
        RECT  1.360 -0.280 2.120 0.280 ;
        RECT  1.080 -0.280 1.360 1.270 ;
        RECT  0.000 -0.280 1.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 3.320 2.800 3.880 ;
        RECT  2.240 2.190 2.520 3.880 ;
        RECT  0.920 3.320 2.240 3.880 ;
        RECT  0.640 2.440 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.320 1.750 1.600 2.280 ;
        RECT  0.680 2.120 1.320 2.280 ;
        RECT  0.680 1.010 0.840 1.290 ;
        RECT  0.520 1.010 0.680 2.280 ;
        RECT  0.440 2.120 0.520 2.280 ;
        RECT  0.160 2.120 0.440 2.400 ;
    END
END NOR2BX2TR

MACRO NOR2BX1TR
    CLASS CORE ;
    FOREIGN NOR2BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.850 1.920 3.160 ;
        RECT  1.200 0.850 1.760 1.130 ;
        RECT  1.600 1.940 1.760 3.160 ;
        END
        ANTENNADIFFAREA 2.508 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.610 1.120 2.070 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.240 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.280 2.000 0.280 ;
        RECT  0.800 -0.280 1.880 0.340 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 3.320 2.000 3.880 ;
        RECT  0.680 2.560 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.360 1.600 1.640 ;
        RECT  1.280 1.290 1.440 2.400 ;
        RECT  1.040 1.290 1.280 1.450 ;
        RECT  0.350 2.240 1.280 2.400 ;
        RECT  0.880 0.910 1.040 1.450 ;
        RECT  0.370 0.910 0.880 1.080 ;
        RECT  0.090 0.800 0.370 1.080 ;
        RECT  0.090 1.940 0.350 2.400 ;
    END
END NOR2BX1TR

MACRO NOR2XLTR
    CLASS CORE ;
    FOREIGN NOR2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.920 1.520 2.760 ;
        RECT  0.960 0.920 1.360 1.080 ;
        RECT  1.280 1.640 1.360 2.760 ;
        RECT  1.040 1.980 1.280 2.260 ;
        RECT  0.660 0.740 0.960 1.080 ;
        END
        ANTENNADIFFAREA 1.316 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.360 0.680 1.640 ;
        RECT  0.080 0.440 0.320 1.640 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.120 1.640 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.510 -0.280 1.600 0.280 ;
        RECT  1.230 -0.280 1.510 0.760 ;
        RECT  0.000 -0.280 1.230 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 3.320 1.600 3.880 ;
        RECT  0.240 1.980 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
END NOR2XLTR

MACRO NOR2X8TR
    CLASS CORE ;
    FOREIGN NOR2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.740 0.600 5.120 2.960 ;
        RECT  4.520 0.600 4.740 1.080 ;
        RECT  4.520 2.060 4.740 2.960 ;
        RECT  4.240 0.440 4.520 1.080 ;
        RECT  4.240 2.060 4.520 3.080 ;
        RECT  3.480 0.600 4.240 1.080 ;
        RECT  2.920 2.060 4.240 2.540 ;
        RECT  3.200 0.440 3.480 1.080 ;
        RECT  2.440 0.600 3.200 1.080 ;
        RECT  2.640 2.060 2.920 3.160 ;
        RECT  1.320 2.060 2.640 2.530 ;
        RECT  2.160 0.440 2.440 1.080 ;
        RECT  1.400 0.600 2.160 1.080 ;
        RECT  1.120 0.440 1.400 1.080 ;
        RECT  1.040 2.060 1.320 3.160 ;
        END
        ANTENNADIFFAREA 12.874 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 1.560 3.760 1.900 ;
        RECT  2.280 1.740 3.480 1.900 ;
        RECT  1.640 1.560 2.280 1.900 ;
        RECT  0.760 1.740 1.640 1.900 ;
        RECT  0.440 1.240 0.760 1.900 ;
        END
        ANTENNAGATEAREA 1.1928 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.320 1.500 4.580 1.840 ;
        RECT  4.080 1.240 4.320 1.840 ;
        RECT  3.120 1.240 4.080 1.400 ;
        RECT  2.440 1.240 3.120 1.580 ;
        RECT  1.200 1.240 2.440 1.400 ;
        RECT  0.920 1.240 1.200 1.580 ;
        END
        ANTENNAGATEAREA 1.1928 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.040 -0.280 5.200 0.280 ;
        RECT  4.760 -0.280 5.040 0.400 ;
        RECT  4.000 -0.280 4.760 0.280 ;
        RECT  3.720 -0.280 4.000 0.400 ;
        RECT  2.960 -0.280 3.720 0.280 ;
        RECT  2.680 -0.280 2.960 0.400 ;
        RECT  1.920 -0.280 2.680 0.280 ;
        RECT  1.640 -0.280 1.920 0.400 ;
        RECT  0.880 -0.280 1.640 0.280 ;
        RECT  0.600 -0.280 0.880 1.040 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 3.320 5.200 3.880 ;
        RECT  3.440 2.930 3.720 3.880 ;
        RECT  2.120 3.320 3.440 3.880 ;
        RECT  1.840 2.930 2.120 3.880 ;
        RECT  0.520 3.320 1.840 3.880 ;
        RECT  0.240 2.060 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
END NOR2X8TR

MACRO NOR2X6TR
    CLASS CORE ;
    FOREIGN NOR2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.500 0.740 3.860 3.100 ;
        RECT  2.780 0.740 3.500 1.100 ;
        RECT  3.080 1.840 3.500 2.560 ;
        RECT  2.200 2.120 3.080 2.480 ;
        RECT  2.500 0.440 2.780 1.100 ;
        RECT  1.820 0.770 2.500 1.100 ;
        RECT  1.920 2.120 2.200 3.160 ;
        RECT  0.540 2.120 1.920 2.480 ;
        RECT  1.540 0.440 1.820 1.100 ;
        RECT  0.860 0.770 1.540 1.100 ;
        RECT  0.580 0.440 0.860 1.100 ;
        RECT  0.260 2.120 0.540 2.970 ;
        END
        ANTENNADIFFAREA 10.884 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.660 1.680 2.880 1.960 ;
        RECT  1.560 1.800 2.660 1.960 ;
        RECT  0.880 1.580 1.560 1.960 ;
        END
        ANTENNAGATEAREA 0.888 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.260 3.340 1.640 ;
        RECT  2.400 1.260 3.180 1.420 ;
        RECT  1.720 1.260 2.400 1.640 ;
        RECT  0.720 1.260 1.720 1.420 ;
        RECT  0.560 1.260 0.720 1.960 ;
        RECT  0.440 1.560 0.560 1.960 ;
        RECT  0.300 1.560 0.440 1.840 ;
        END
        ANTENNAGATEAREA 0.888 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.300 -0.280 4.000 0.280 ;
        RECT  3.020 -0.280 3.300 0.400 ;
        RECT  2.300 -0.280 3.020 0.280 ;
        RECT  2.020 -0.280 2.300 0.610 ;
        RECT  1.340 -0.280 2.020 0.280 ;
        RECT  1.060 -0.280 1.340 0.610 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 1.310 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 3.320 4.000 3.880 ;
        RECT  2.720 2.930 3.000 3.880 ;
        RECT  1.360 3.320 2.720 3.880 ;
        RECT  1.080 2.690 1.360 3.880 ;
        RECT  0.000 3.320 1.080 3.880 ;
        END
    END VDD
END NOR2X6TR

MACRO NOR2X4TR
    CLASS CORE ;
    FOREIGN NOR2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.960 3.120 2.760 ;
        RECT  2.850 0.960 2.970 3.160 ;
        RECT  2.000 0.960 2.850 1.200 ;
        RECT  2.480 2.030 2.850 3.160 ;
        RECT  1.370 2.120 2.480 2.360 ;
        RECT  1.720 0.440 2.000 1.200 ;
        RECT  0.960 0.830 1.720 1.080 ;
        RECT  1.090 2.120 1.370 2.970 ;
        RECT  0.680 0.440 0.960 1.080 ;
        END
        ANTENNADIFFAREA 7.207 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.680 2.200 1.960 ;
        RECT  0.760 1.800 1.920 1.960 ;
        RECT  0.480 1.580 0.760 1.960 ;
        RECT  0.440 1.640 0.480 1.960 ;
        END
        ANTENNAGATEAREA 0.6168 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.360 2.690 1.640 ;
        RECT  1.570 1.360 2.410 1.520 ;
        RECT  1.560 1.360 1.570 1.640 ;
        RECT  1.240 1.240 1.560 1.640 ;
        RECT  0.920 1.360 1.240 1.640 ;
        END
        ANTENNAGATEAREA 0.6168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 -0.280 3.200 0.280 ;
        RECT  2.520 0.500 2.920 0.770 ;
        RECT  2.240 -0.280 2.520 0.770 ;
        RECT  1.480 -0.280 2.240 0.280 ;
        RECT  1.200 -0.280 1.480 0.400 ;
        RECT  0.440 -0.280 1.200 0.280 ;
        RECT  0.160 -0.280 0.440 1.310 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 3.320 3.200 3.880 ;
        RECT  1.890 2.530 2.170 3.880 ;
        RECT  0.570 3.320 1.890 3.880 ;
        RECT  0.250 2.120 0.570 3.880 ;
        RECT  0.000 3.320 0.250 3.880 ;
        END
    END VDD
END NOR2X4TR

MACRO NOR2X2TR
    CLASS CORE ;
    FOREIGN NOR2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.240 1.920 2.360 ;
        RECT  1.680 0.920 1.760 2.360 ;
        RECT  1.600 0.920 1.680 2.300 ;
        RECT  1.300 0.920 1.600 1.080 ;
        RECT  1.190 2.120 1.600 2.300 ;
        RECT  1.020 0.440 1.300 1.080 ;
        RECT  0.910 2.120 1.190 2.870 ;
        END
        ANTENNADIFFAREA 3.168 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.440 1.640 ;
        RECT  0.720 1.240 1.280 1.400 ;
        RECT  0.540 1.240 0.720 1.560 ;
        RECT  0.310 1.240 0.540 1.870 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.120 1.960 ;
        RECT  0.800 1.740 0.880 1.960 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.820 -0.280 2.000 0.280 ;
        RECT  1.540 -0.280 1.820 0.760 ;
        RECT  0.830 -0.280 1.540 0.280 ;
        RECT  0.530 -0.280 0.830 1.080 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 3.320 2.000 3.880 ;
        RECT  1.640 3.220 1.880 3.880 ;
        RECT  0.410 3.320 1.640 3.880 ;
        RECT  0.110 2.150 0.410 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
END NOR2X2TR

MACRO NOR2X1TR
    CLASS CORE ;
    FOREIGN NOR2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.920 1.520 3.160 ;
        RECT  0.920 0.920 1.360 1.080 ;
        RECT  1.280 1.910 1.360 3.160 ;
        RECT  1.040 1.910 1.280 2.750 ;
        RECT  0.640 0.800 0.920 1.080 ;
        END
        ANTENNADIFFAREA 2.172 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.430 0.680 1.710 ;
        RECT  0.320 1.240 0.360 1.710 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.160 1.700 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 -0.280 1.600 0.280 ;
        RECT  1.160 -0.280 1.470 0.760 ;
        RECT  0.450 -0.280 1.160 0.280 ;
        RECT  0.150 -0.280 0.450 1.080 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 3.320 1.600 3.880 ;
        RECT  0.240 2.530 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
END NOR2X1TR

MACRO NAND4BBXLTR
    CLASS CORE ;
    FOREIGN NAND4BBXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.690 2.490 0.990 ;
        RECT  2.240 1.910 2.360 2.600 ;
        RECT  2.240 0.440 2.330 0.990 ;
        RECT  2.080 0.440 2.240 2.600 ;
        RECT  1.090 2.440 2.080 2.600 ;
        END
        ANTENNADIFFAREA 0.832 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.270 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.540 1.790 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.240 0.720 1.680 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.440 3.520 1.750 ;
        RECT  2.970 1.470 3.240 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.280 3.600 0.280 ;
        RECT  0.690 -0.280 0.970 0.760 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 3.320 3.600 3.880 ;
        RECT  2.560 2.270 2.840 3.880 ;
        RECT  1.770 3.260 2.560 3.880 ;
        RECT  1.490 3.200 1.770 3.880 ;
        RECT  0.890 3.260 1.490 3.880 ;
        RECT  0.610 2.440 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.070 1.910 3.360 2.370 ;
        RECT  2.810 1.910 3.070 2.070 ;
        RECT  2.810 1.030 2.950 1.310 ;
        RECT  2.650 1.030 2.810 2.070 ;
        RECT  2.400 1.430 2.650 1.710 ;
        RECT  1.700 0.920 1.920 2.280 ;
        RECT  0.410 0.920 1.700 1.080 ;
        RECT  0.360 2.120 1.700 2.280 ;
        RECT  0.130 0.780 0.410 1.080 ;
        RECT  0.090 2.120 0.360 2.530 ;
    END
END NAND4BBXLTR

MACRO NAND4BBX4TR
    CLASS CORE ;
    FOREIGN NAND4BBX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.520 8.320 3.050 ;
        RECT  5.560 0.520 8.080 0.760 ;
        RECT  7.520 2.810 8.080 3.050 ;
        RECT  7.280 2.240 7.520 3.050 ;
        RECT  1.060 2.810 7.280 3.050 ;
        RECT  5.280 0.440 5.560 1.070 ;
        RECT  2.680 0.830 5.280 1.070 ;
        RECT  2.400 0.440 2.680 1.070 ;
        END
        ANTENNADIFFAREA 11.88 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.000 1.240 7.120 1.630 ;
        RECT  6.840 1.240 7.000 2.650 ;
        RECT  1.120 2.490 6.840 2.650 ;
        RECT  0.960 1.610 1.120 2.650 ;
        END
        ANTENNAGATEAREA 0.6696 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.520 1.610 6.640 1.890 ;
        RECT  6.360 1.610 6.520 2.270 ;
        RECT  1.580 2.050 6.360 2.270 ;
        RECT  1.420 1.610 1.580 2.270 ;
        RECT  1.280 1.610 1.420 1.960 ;
        END
        ANTENNAGATEAREA 0.6696 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.240 7.920 1.760 ;
        RECT  7.600 1.490 7.680 1.760 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.640 0.790 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.160 -0.280 8.400 0.280 ;
        RECT  6.880 -0.280 7.160 0.340 ;
        RECT  4.120 -0.280 6.880 0.280 ;
        RECT  3.840 -0.280 4.120 0.670 ;
        RECT  1.080 -0.280 3.840 0.280 ;
        RECT  0.770 -0.280 1.080 1.010 ;
        RECT  0.000 -0.280 0.770 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.440 3.320 8.400 3.880 ;
        RECT  7.160 3.210 7.440 3.880 ;
        RECT  6.400 3.320 7.160 3.880 ;
        RECT  6.120 3.210 6.400 3.880 ;
        RECT  5.360 3.320 6.120 3.880 ;
        RECT  5.080 3.210 5.360 3.880 ;
        RECT  2.900 3.260 5.080 3.880 ;
        RECT  2.620 3.210 2.900 3.880 ;
        RECT  1.860 3.320 2.620 3.880 ;
        RECT  1.580 3.210 1.860 3.880 ;
        RECT  0.800 3.320 1.580 3.880 ;
        RECT  0.580 2.120 0.800 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.680 1.920 7.900 2.310 ;
        RECT  7.440 0.920 7.880 1.080 ;
        RECT  7.440 1.920 7.680 2.080 ;
        RECT  7.280 0.920 7.440 2.080 ;
        RECT  6.080 0.920 7.280 1.080 ;
        RECT  5.920 0.920 6.080 1.890 ;
        RECT  4.760 1.610 5.920 1.890 ;
        RECT  0.420 1.270 5.760 1.430 ;
        RECT  3.200 1.610 4.760 1.770 ;
        RECT  2.920 1.610 3.200 1.890 ;
        RECT  2.100 1.610 2.920 1.770 ;
        RECT  1.820 1.610 2.100 1.890 ;
        RECT  0.240 0.540 0.420 1.430 ;
        RECT  0.240 2.160 0.380 3.140 ;
        RECT  0.080 0.540 0.240 3.140 ;
    END
END NAND4BBX4TR

MACRO NAND4BBX2TR
    CLASS CORE ;
    FOREIGN NAND4BBX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.500 0.520 2.780 1.130 ;
        RECT  2.340 2.840 2.620 3.120 ;
        RECT  0.320 0.640 2.500 0.800 ;
        RECT  1.580 2.840 2.340 3.000 ;
        RECT  1.300 2.840 1.580 3.120 ;
        RECT  0.260 2.840 1.300 3.000 ;
        RECT  0.260 0.440 0.320 1.560 ;
        RECT  0.100 0.440 0.260 3.000 ;
        RECT  0.080 0.440 0.100 1.560 ;
        END
        ANTENNADIFFAREA 5.904 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 2.390 3.740 2.760 ;
        RECT  1.420 2.520 3.240 2.680 ;
        RECT  1.200 1.510 1.420 2.680 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.580 1.630 3.700 1.910 ;
        RECT  3.420 1.630 3.580 2.230 ;
        RECT  1.960 2.070 3.420 2.230 ;
        RECT  1.860 2.040 1.960 2.360 ;
        RECT  1.640 1.670 1.860 2.360 ;
        RECT  1.580 1.670 1.640 1.950 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.640 4.360 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.480 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.220 -0.280 4.800 0.280 ;
        RECT  3.940 -0.280 4.220 1.040 ;
        RECT  1.300 -0.280 3.940 0.280 ;
        RECT  1.020 -0.280 1.300 0.400 ;
        RECT  0.000 -0.280 1.020 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.180 3.320 4.800 3.880 ;
        RECT  3.900 2.440 4.180 3.880 ;
        RECT  3.140 3.260 3.900 3.880 ;
        RECT  2.860 3.200 3.140 3.880 ;
        RECT  2.100 3.320 2.860 3.880 ;
        RECT  1.820 3.200 2.100 3.880 ;
        RECT  1.060 3.320 1.820 3.880 ;
        RECT  0.780 3.200 1.060 3.880 ;
        RECT  0.000 3.320 0.780 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.540 0.960 4.700 2.930 ;
        RECT  4.420 0.960 4.540 1.470 ;
        RECT  4.420 2.340 4.540 2.930 ;
        RECT  3.260 1.310 4.420 1.470 ;
        RECT  3.100 1.310 3.260 1.910 ;
        RECT  2.980 1.630 3.100 1.910 ;
        RECT  2.060 1.690 2.980 1.850 ;
        RECT  1.740 1.350 2.820 1.510 ;
        RECT  1.580 1.160 1.740 1.510 ;
        RECT  1.040 1.160 1.580 1.320 ;
        RECT  0.880 1.160 1.040 2.280 ;
        RECT  0.780 1.160 0.880 1.320 ;
        RECT  0.700 2.120 0.880 2.280 ;
        RECT  0.500 0.960 0.780 1.320 ;
        RECT  0.420 2.120 0.700 2.400 ;
    END
END NAND4BBX2TR

MACRO NAND4BBX1TR
    CLASS CORE ;
    FOREIGN NAND4BBX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.440 2.490 1.190 ;
        RECT  2.240 1.910 2.360 2.600 ;
        RECT  2.080 0.440 2.240 2.600 ;
        RECT  1.090 2.440 2.080 2.600 ;
        END
        ANTENNADIFFAREA 3.776 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.270 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.540 1.790 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.240 0.720 1.680 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.440 3.520 1.750 ;
        RECT  2.970 1.470 3.240 1.750 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.280 3.600 0.280 ;
        RECT  0.690 -0.280 0.970 0.640 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 3.320 3.600 3.880 ;
        RECT  2.560 2.270 2.840 3.880 ;
        RECT  1.770 3.260 2.560 3.880 ;
        RECT  1.490 3.200 1.770 3.880 ;
        RECT  0.890 3.260 1.490 3.880 ;
        RECT  0.610 2.440 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.170 1.910 3.450 2.190 ;
        RECT  2.810 1.910 3.170 2.070 ;
        RECT  2.810 1.030 2.950 1.310 ;
        RECT  2.650 1.030 2.810 2.070 ;
        RECT  2.400 1.430 2.650 1.710 ;
        RECT  1.700 0.920 1.920 2.280 ;
        RECT  0.410 0.920 1.700 1.080 ;
        RECT  0.090 2.120 1.700 2.280 ;
        RECT  0.130 0.800 0.410 1.080 ;
    END
END NAND4BBX1TR

MACRO NAND4BXLTR
    CLASS CORE ;
    FOREIGN NAND4BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.600 2.720 2.290 ;
        RECT  2.500 0.600 2.560 0.760 ;
        RECT  2.320 2.120 2.560 2.290 ;
        RECT  2.040 0.440 2.500 0.760 ;
        RECT  2.030 2.120 2.320 2.360 ;
        RECT  1.370 2.120 2.030 2.290 ;
        RECT  1.080 2.120 1.370 2.360 ;
        END
        ANTENNADIFFAREA 0.832 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.240 1.120 1.740 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.450 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.840 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.380 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.280 2.800 0.280 ;
        RECT  0.750 -0.280 1.050 0.760 ;
        RECT  0.000 -0.280 0.750 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.430 3.190 2.710 3.880 ;
        RECT  1.710 3.320 2.430 3.880 ;
        RECT  0.700 3.030 1.710 3.880 ;
        RECT  0.000 3.320 0.700 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.920 2.400 1.520 ;
        RECT  0.700 0.920 2.120 1.080 ;
        RECT  0.540 0.920 0.700 2.710 ;
        RECT  0.400 0.920 0.540 1.080 ;
        RECT  0.160 2.550 0.540 2.710 ;
        RECT  0.120 0.800 0.400 1.080 ;
    END
END NAND4BXLTR

MACRO NAND4BX4TR
    CLASS CORE ;
    FOREIGN NAND4BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.880 1.120 7.120 3.070 ;
        RECT  6.720 1.120 6.880 1.360 ;
        RECT  6.620 2.830 6.880 3.070 ;
        RECT  6.480 0.610 6.720 1.360 ;
        RECT  6.260 2.830 6.620 3.160 ;
        RECT  5.350 0.830 6.480 1.070 ;
        RECT  5.580 2.830 6.260 3.070 ;
        RECT  5.220 2.830 5.580 3.160 ;
        RECT  5.060 0.440 5.350 1.070 ;
        RECT  2.380 2.830 5.220 3.070 ;
        RECT  2.460 0.830 5.060 1.070 ;
        RECT  2.160 0.440 2.460 1.070 ;
        RECT  2.100 2.830 2.380 3.160 ;
        RECT  1.360 2.830 2.100 3.070 ;
        RECT  1.050 2.830 1.360 3.160 ;
        END
        ANTENNADIFFAREA 11.808 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.610 6.720 1.890 ;
        RECT  6.500 1.610 6.670 2.660 ;
        RECT  1.120 2.500 6.500 2.660 ;
        RECT  0.920 1.610 1.120 2.660 ;
        RECT  0.880 1.610 0.920 1.970 ;
        END
        ANTENNAGATEAREA 0.66 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.610 6.320 2.340 ;
        RECT  1.520 2.120 6.050 2.340 ;
        RECT  1.280 1.610 1.520 2.340 ;
        END
        ANTENNAGATEAREA 0.66 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.610 5.790 1.890 ;
        RECT  2.980 1.730 4.540 1.890 ;
        RECT  2.700 1.610 2.980 1.890 ;
        RECT  1.920 1.610 2.700 1.770 ;
        RECT  1.680 1.610 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.66 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.590 0.720 2.410 ;
        RECT  0.440 1.590 0.480 1.860 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.100 -0.280 7.200 0.280 ;
        RECT  6.880 -0.280 7.100 0.750 ;
        RECT  3.900 -0.280 6.880 0.280 ;
        RECT  3.620 -0.280 3.900 0.670 ;
        RECT  0.900 -0.280 3.620 0.280 ;
        RECT  0.620 -0.280 0.900 1.060 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.100 3.320 7.200 3.880 ;
        RECT  6.820 3.230 7.100 3.880 ;
        RECT  6.060 3.320 6.820 3.880 ;
        RECT  5.780 3.230 6.060 3.880 ;
        RECT  5.030 3.320 5.780 3.880 ;
        RECT  4.750 3.230 5.030 3.880 ;
        RECT  2.900 3.260 4.750 3.880 ;
        RECT  2.620 3.230 2.900 3.880 ;
        RECT  1.860 3.320 2.620 3.880 ;
        RECT  1.580 3.230 1.860 3.880 ;
        RECT  0.860 3.320 1.580 3.880 ;
        RECT  0.580 2.930 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.380 1.230 5.540 1.430 ;
        RECT  0.260 0.500 0.380 1.430 ;
        RECT  0.260 2.120 0.320 3.160 ;
        RECT  0.100 0.500 0.260 3.160 ;
    END
END NAND4BX4TR

MACRO NAND4BX2TR
    CLASS CORE ;
    FOREIGN NAND4BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 3.920 3.100 ;
        RECT  3.680 1.240 3.760 2.360 ;
        RECT  2.290 2.940 3.760 3.100 ;
        RECT  2.810 1.240 3.680 1.440 ;
        RECT  2.650 0.990 2.810 1.440 ;
        RECT  2.440 0.990 2.650 1.150 ;
        RECT  2.160 0.870 2.440 1.150 ;
        RECT  2.010 2.940 2.290 3.160 ;
        RECT  1.250 2.940 2.010 3.100 ;
        RECT  0.970 2.940 1.250 3.160 ;
        END
        ANTENNADIFFAREA 5.889 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 2.620 3.520 2.780 ;
        RECT  0.880 1.660 1.120 2.780 ;
        END
        ANTENNAGATEAREA 0.3384 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.600 3.520 2.460 ;
        RECT  1.520 2.300 3.260 2.460 ;
        RECT  1.280 1.700 1.520 2.460 ;
        END
        ANTENNAGATEAREA 0.3384 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.920 3.040 2.140 ;
        RECT  1.680 1.640 1.960 2.140 ;
        END
        ANTENNAGATEAREA 0.3384 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.630 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.880 -0.280 4.000 0.280 ;
        RECT  3.600 -0.280 3.880 0.730 ;
        RECT  0.890 -0.280 3.600 0.280 ;
        RECT  0.610 -0.280 0.890 1.150 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.810 3.320 4.000 3.880 ;
        RECT  2.530 3.260 2.810 3.880 ;
        RECT  1.770 3.320 2.530 3.880 ;
        RECT  1.490 3.260 1.770 3.880 ;
        RECT  0.730 3.320 1.490 3.880 ;
        RECT  0.450 3.200 0.730 3.880 ;
        RECT  0.000 3.320 0.450 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.210 1.310 2.490 1.620 ;
        RECT  0.370 1.310 2.210 1.470 ;
        RECT  0.240 0.990 0.370 1.470 ;
        RECT  0.240 2.120 0.310 2.650 ;
        RECT  0.080 0.990 0.240 2.650 ;
    END
END NAND4BX2TR

MACRO NAND4BX1TR
    CLASS CORE ;
    FOREIGN NAND4BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.600 2.720 2.290 ;
        RECT  2.500 0.600 2.560 0.760 ;
        RECT  2.320 2.130 2.560 2.290 ;
        RECT  2.040 0.440 2.500 0.760 ;
        RECT  2.080 2.130 2.320 2.760 ;
        RECT  1.370 2.130 2.080 2.290 ;
        RECT  1.080 2.130 1.370 2.440 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.240 1.120 1.740 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.450 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.960 1.780 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.580 0.380 1.860 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.280 2.800 0.280 ;
        RECT  0.750 -0.280 1.050 0.700 ;
        RECT  0.000 -0.280 0.750 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.430 3.190 2.710 3.880 ;
        RECT  1.790 3.320 2.430 3.880 ;
        RECT  0.680 3.030 1.790 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.920 2.400 1.520 ;
        RECT  0.700 0.920 2.120 1.080 ;
        RECT  0.540 0.920 0.700 2.750 ;
        RECT  0.400 0.920 0.540 1.080 ;
        RECT  0.400 2.590 0.540 2.750 ;
        RECT  0.120 0.800 0.400 1.080 ;
        RECT  0.120 2.590 0.400 2.870 ;
    END
END NAND4BX1TR

MACRO NAND4XLTR
    CLASS CORE ;
    FOREIGN NAND4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.440 2.140 0.610 ;
        RECT  1.870 0.440 1.920 0.760 ;
        RECT  1.810 0.440 1.870 2.160 ;
        RECT  1.710 0.440 1.810 2.510 ;
        RECT  1.680 0.440 1.710 0.760 ;
        RECT  1.530 2.000 1.710 2.510 ;
        RECT  0.850 2.000 1.530 2.160 ;
        RECT  0.570 2.000 0.850 2.500 ;
        END
        ANTENNADIFFAREA 0.832 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.590 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.840 1.120 1.840 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.550 1.840 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.840 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.680 -0.280 2.400 0.280 ;
        RECT  0.360 -0.280 0.680 0.680 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 3.320 2.400 3.880 ;
        RECT  2.000 2.290 2.290 3.880 ;
        RECT  1.340 3.320 2.000 3.880 ;
        RECT  1.040 2.320 1.340 3.880 ;
        RECT  0.400 3.320 1.040 3.880 ;
        RECT  0.120 2.970 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND4XLTR

MACRO NAND4X8TR
    CLASS CORE ;
    FOREIGN NAND4X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.830 0.770 12.320 3.160 ;
        RECT  11.720 0.770 11.830 1.360 ;
        RECT  9.200 2.700 11.830 3.160 ;
        RECT  11.080 0.640 11.720 1.360 ;
        RECT  10.780 0.640 11.080 1.160 ;
        RECT  10.560 0.440 10.780 1.160 ;
        RECT  10.500 0.440 10.560 0.940 ;
        RECT  7.060 0.500 10.500 0.940 ;
        RECT  2.140 2.740 9.200 3.160 ;
        RECT  6.740 0.500 7.060 1.200 ;
        RECT  4.240 0.770 6.740 1.200 ;
        RECT  3.960 0.440 4.240 1.200 ;
        RECT  1.720 2.120 2.140 3.160 ;
        RECT  0.920 2.120 1.720 2.610 ;
        RECT  0.640 2.120 0.920 3.160 ;
        RECT  0.580 0.500 0.860 1.160 ;
        RECT  0.400 2.120 0.640 2.610 ;
        RECT  0.400 0.730 0.580 1.160 ;
        RECT  0.090 0.730 0.400 2.610 ;
        END
        ANTENNADIFFAREA 23.244 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 2.380 11.590 2.540 ;
        RECT  8.680 2.090 8.960 2.580 ;
        RECT  2.730 2.420 8.680 2.580 ;
        RECT  2.570 1.560 2.730 2.580 ;
        RECT  2.480 1.560 2.570 2.360 ;
        RECT  2.080 1.560 2.480 1.780 ;
        END
        ANTENNAGATEAREA 1.2888 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.420 1.870 11.670 2.200 ;
        RECT  9.760 2.040 11.420 2.200 ;
        RECT  9.600 1.740 9.760 2.200 ;
        RECT  8.020 1.740 9.600 1.900 ;
        RECT  7.860 1.740 8.020 2.260 ;
        RECT  3.160 2.100 7.860 2.260 ;
        RECT  3.000 1.240 3.160 2.260 ;
        RECT  1.920 1.240 3.000 1.400 ;
        RECT  1.680 1.240 1.920 1.900 ;
        RECT  1.660 1.620 1.680 1.900 ;
        END
        ANTENNAGATEAREA 1.2888 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.200 1.520 11.380 1.680 ;
        RECT  11.040 1.520 11.200 1.880 ;
        RECT  10.080 1.720 11.040 1.880 ;
        RECT  9.920 1.420 10.080 1.880 ;
        RECT  7.700 1.420 9.920 1.580 ;
        RECT  7.540 1.420 7.700 1.900 ;
        RECT  3.480 1.740 7.540 1.900 ;
        RECT  3.320 0.920 3.480 1.900 ;
        RECT  1.500 0.920 3.320 1.080 ;
        RECT  1.340 0.920 1.500 1.920 ;
        RECT  1.120 1.640 1.340 1.920 ;
        RECT  0.880 1.640 1.120 1.960 ;
        END
        ANTENNAGATEAREA 1.2888 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.400 1.360 10.880 1.520 ;
        RECT  10.240 1.100 10.400 1.520 ;
        RECT  7.380 1.100 10.240 1.260 ;
        RECT  7.220 1.100 7.380 1.520 ;
        RECT  3.800 1.360 7.220 1.520 ;
        RECT  3.640 0.600 3.800 1.520 ;
        RECT  3.160 0.600 3.640 0.760 ;
        RECT  2.880 0.440 3.160 0.760 ;
        RECT  1.180 0.600 2.880 0.760 ;
        RECT  1.020 0.600 1.180 1.480 ;
        RECT  0.720 1.320 1.020 1.480 ;
        RECT  0.560 1.320 0.720 1.600 ;
        END
        ANTENNAGATEAREA 1.2888 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.300 -0.280 12.400 0.280 ;
        RECT  12.020 -0.280 12.300 0.610 ;
        RECT  9.080 -0.280 12.020 0.280 ;
        RECT  8.400 -0.280 9.080 0.340 ;
        RECT  5.680 -0.280 8.400 0.280 ;
        RECT  5.400 -0.280 5.680 0.610 ;
        RECT  2.700 -0.280 5.400 0.280 ;
        RECT  2.070 -0.280 2.700 0.400 ;
        RECT  0.000 -0.280 2.070 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 3.320 12.400 3.880 ;
        RECT  1.200 2.800 1.480 3.880 ;
        RECT  0.400 3.320 1.200 3.880 ;
        RECT  0.120 2.790 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND4X8TR

MACRO NAND4X6TR
    CLASS CORE ;
    FOREIGN NAND4X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.580 0.640 8.940 3.100 ;
        RECT  8.280 0.640 8.580 1.360 ;
        RECT  1.960 2.730 8.580 3.100 ;
        RECT  7.100 0.810 8.280 1.170 ;
        RECT  6.820 0.440 7.100 1.170 ;
        RECT  4.220 0.810 6.820 1.170 ;
        RECT  3.940 0.440 4.220 1.170 ;
        RECT  1.680 2.120 1.960 3.100 ;
        RECT  0.920 2.120 1.680 2.480 ;
        RECT  0.640 2.120 0.920 3.160 ;
        RECT  0.320 0.790 0.740 1.080 ;
        RECT  0.320 2.120 0.640 2.480 ;
        RECT  0.090 0.790 0.320 2.480 ;
        END
        ANTENNADIFFAREA 17.398 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.240 1.650 8.400 2.570 ;
        RECT  2.760 2.410 8.240 2.570 ;
        RECT  2.600 1.640 2.760 2.570 ;
        RECT  2.100 1.640 2.600 1.960 ;
        END
        ANTENNAGATEAREA 0.9336 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.900 1.650 8.020 1.930 ;
        RECT  7.740 1.650 7.900 2.250 ;
        RECT  3.140 2.090 7.740 2.250 ;
        RECT  2.980 1.320 3.140 2.250 ;
        RECT  1.920 1.320 2.980 1.480 ;
        RECT  1.760 1.320 1.920 1.960 ;
        RECT  1.540 1.640 1.760 1.960 ;
        END
        ANTENNAGATEAREA 0.9336 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.300 1.630 7.580 1.930 ;
        RECT  3.460 1.710 7.300 1.930 ;
        RECT  3.300 1.000 3.460 1.930 ;
        RECT  1.380 1.000 3.300 1.160 ;
        RECT  1.220 1.000 1.380 1.960 ;
        RECT  0.880 1.640 1.220 1.960 ;
        END
        ANTENNAGATEAREA 0.9336 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.780 1.330 6.980 1.490 ;
        RECT  3.620 0.680 3.780 1.490 ;
        RECT  1.060 0.680 3.620 0.840 ;
        RECT  0.900 0.680 1.060 1.480 ;
        RECT  0.720 1.240 0.900 1.480 ;
        RECT  0.480 1.240 0.720 1.740 ;
        END
        ANTENNAGATEAREA 0.9336 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.580 -0.280 9.200 0.280 ;
        RECT  8.300 -0.280 8.580 0.400 ;
        RECT  5.660 -0.280 8.300 0.280 ;
        RECT  5.380 -0.280 5.660 0.650 ;
        RECT  2.480 -0.280 5.380 0.280 ;
        RECT  2.200 -0.280 2.480 0.400 ;
        RECT  0.000 -0.280 2.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.740 3.320 9.200 3.880 ;
        RECT  8.460 3.260 8.740 3.880 ;
        RECT  7.700 3.320 8.460 3.880 ;
        RECT  7.420 3.260 7.700 3.880 ;
        RECT  6.660 3.320 7.420 3.880 ;
        RECT  4.280 3.260 6.660 3.880 ;
        RECT  3.520 3.320 4.280 3.880 ;
        RECT  3.240 3.260 3.520 3.880 ;
        RECT  2.480 3.320 3.240 3.880 ;
        RECT  2.200 3.260 2.480 3.880 ;
        RECT  1.440 3.320 2.200 3.880 ;
        RECT  1.160 2.780 1.440 3.880 ;
        RECT  0.400 3.320 1.160 3.880 ;
        RECT  0.120 2.740 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND4X6TR

MACRO NAND4X4TR
    CLASS CORE ;
    FOREIGN NAND4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.730 0.840 6.960 3.020 ;
        RECT  6.720 0.640 6.730 3.020 ;
        RECT  6.480 0.640 6.720 1.360 ;
        RECT  6.370 2.800 6.720 3.020 ;
        RECT  5.010 0.840 6.480 1.080 ;
        RECT  6.090 2.800 6.370 3.140 ;
        RECT  5.330 2.800 6.090 3.020 ;
        RECT  5.050 2.800 5.330 3.140 ;
        RECT  2.040 2.800 5.050 3.040 ;
        RECT  4.730 0.730 5.010 1.080 ;
        RECT  2.130 0.860 4.730 1.080 ;
        RECT  1.850 0.750 2.130 1.080 ;
        RECT  1.760 2.800 2.040 3.140 ;
        RECT  1.000 2.800 1.760 3.040 ;
        RECT  0.720 2.800 1.000 3.140 ;
        END
        ANTENNADIFFAREA 11.592 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.660 6.510 2.640 ;
        RECT  0.720 2.480 6.350 2.640 ;
        RECT  0.560 1.640 0.720 2.640 ;
        RECT  0.440 1.640 0.560 1.960 ;
        END
        ANTENNAGATEAREA 0.6672 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.650 5.970 1.930 ;
        RECT  5.690 1.650 5.850 2.320 ;
        RECT  1.140 2.100 5.690 2.320 ;
        RECT  1.120 1.710 1.140 2.320 ;
        RECT  0.880 1.240 1.120 2.320 ;
        END
        ANTENNAGATEAREA 0.6672 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 1.660 5.530 1.940 ;
        RECT  4.490 1.780 5.250 1.940 ;
        RECT  4.210 1.720 4.490 1.940 ;
        RECT  2.650 1.780 4.210 1.940 ;
        RECT  2.370 1.720 2.650 1.940 ;
        RECT  1.640 1.780 2.370 1.940 ;
        RECT  1.520 1.650 1.640 1.940 ;
        RECT  1.320 0.840 1.520 1.940 ;
        RECT  1.280 0.840 1.320 1.160 ;
        END
        ANTENNAGATEAREA 0.6672 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.770 1.330 5.050 1.610 ;
        RECT  2.360 1.400 4.770 1.560 ;
        RECT  2.260 1.240 2.360 1.560 ;
        RECT  1.960 1.240 2.260 1.590 ;
        END
        ANTENNAGATEAREA 0.6672 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 -0.280 7.200 0.280 ;
        RECT  6.250 -0.280 6.530 0.480 ;
        RECT  3.570 -0.280 6.250 0.280 ;
        RECT  3.290 -0.280 3.570 0.700 ;
        RECT  0.680 -0.280 3.290 0.280 ;
        RECT  0.400 -0.280 0.680 1.260 ;
        RECT  0.000 -0.280 0.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.890 3.320 7.200 3.880 ;
        RECT  6.610 3.200 6.890 3.880 ;
        RECT  5.850 3.320 6.610 3.880 ;
        RECT  5.570 3.200 5.850 3.880 ;
        RECT  4.810 3.320 5.570 3.880 ;
        RECT  4.530 3.200 4.810 3.880 ;
        RECT  2.560 3.260 4.530 3.880 ;
        RECT  2.280 3.200 2.560 3.880 ;
        RECT  1.520 3.320 2.280 3.880 ;
        RECT  1.240 3.200 1.520 3.880 ;
        RECT  0.400 3.320 1.240 3.880 ;
        RECT  0.120 2.190 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND4X4TR

MACRO NAND4X2TR
    CLASS CORE ;
    FOREIGN NAND4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.030 3.470 2.940 ;
        RECT  2.760 1.030 3.310 1.190 ;
        RECT  1.890 2.780 3.310 2.940 ;
        RECT  2.480 0.800 2.760 1.190 ;
        RECT  1.970 0.800 2.480 0.960 ;
        RECT  1.690 0.800 1.970 1.080 ;
        RECT  1.610 2.780 1.890 3.060 ;
        RECT  0.850 2.780 1.610 2.940 ;
        RECT  0.570 2.780 0.850 3.060 ;
        END
        ANTENNADIFFAREA 5.652 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.990 1.460 3.150 2.620 ;
        RECT  0.670 2.460 2.990 2.620 ;
        RECT  0.670 1.240 0.720 1.560 ;
        RECT  0.510 1.240 0.670 2.620 ;
        RECT  0.290 1.240 0.510 1.680 ;
        END
        ANTENNAGATEAREA 0.3288 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 2.140 2.810 2.300 ;
        RECT  0.960 1.640 1.120 2.300 ;
        RECT  0.880 1.640 0.960 1.980 ;
        RECT  0.830 1.720 0.880 1.980 ;
        END
        ANTENNAGATEAREA 0.3288 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.760 2.490 1.920 ;
        RECT  1.280 1.240 1.560 1.920 ;
        END
        ANTENNAGATEAREA 0.3288 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.240 2.320 1.600 ;
        END
        ANTENNAGATEAREA 0.3288 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.410 -0.280 3.600 0.280 ;
        RECT  3.130 -0.280 3.410 0.870 ;
        RECT  0.480 -0.280 3.130 0.280 ;
        RECT  0.200 -0.280 0.480 0.990 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 3.320 3.600 3.880 ;
        RECT  2.130 3.200 2.410 3.880 ;
        RECT  1.370 3.320 2.130 3.880 ;
        RECT  1.090 3.200 1.370 3.880 ;
        RECT  0.350 3.320 1.090 3.880 ;
        RECT  0.090 2.050 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END NAND4X2TR

MACRO NAND4X1TR
    CLASS CORE ;
    FOREIGN NAND4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.440 2.140 0.610 ;
        RECT  1.870 0.440 1.920 0.760 ;
        RECT  1.810 0.440 1.870 2.160 ;
        RECT  1.710 0.440 1.810 2.510 ;
        RECT  1.680 0.440 1.710 0.760 ;
        RECT  1.530 2.000 1.710 2.510 ;
        RECT  0.850 2.000 1.530 2.160 ;
        RECT  0.570 2.000 0.850 2.500 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.590 1.520 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.840 1.120 1.840 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.550 1.840 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.840 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.680 -0.280 2.400 0.280 ;
        RECT  0.360 -0.280 0.680 0.680 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 3.320 2.400 3.880 ;
        RECT  2.000 2.290 2.280 3.880 ;
        RECT  1.320 3.320 2.000 3.880 ;
        RECT  1.040 2.320 1.320 3.880 ;
        RECT  0.360 3.320 1.040 3.880 ;
        RECT  0.080 2.120 0.360 3.880 ;
        RECT  0.000 3.320 0.080 3.880 ;
        END
    END VDD
END NAND4X1TR

MACRO NAND3BXLTR
    CLASS CORE ;
    FOREIGN NAND3BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.440 2.320 2.720 ;
        RECT  2.080 0.440 2.150 1.560 ;
        RECT  1.090 2.440 2.150 2.720 ;
        RECT  1.850 0.840 2.080 1.160 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.910 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.510 1.590 1.960 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.550 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.280 2.400 0.280 ;
        RECT  0.690 -0.280 0.970 1.080 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 3.320 2.400 3.880 ;
        RECT  1.480 3.090 1.780 3.880 ;
        RECT  0.890 3.260 1.480 3.880 ;
        RECT  0.610 2.460 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.830 1.760 1.990 2.280 ;
        RECT  0.370 2.120 1.830 2.280 ;
        RECT  0.250 1.030 0.410 1.350 ;
        RECT  0.250 2.120 0.370 2.620 ;
        RECT  0.090 1.030 0.250 2.620 ;
    END
END NAND3BXLTR

MACRO NAND3BX4TR
    CLASS CORE ;
    FOREIGN NAND3BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 0.750 4.720 2.340 ;
        RECT  4.480 0.440 4.570 2.340 ;
        RECT  4.290 0.440 4.480 1.180 ;
        RECT  4.320 2.040 4.480 2.340 ;
        RECT  4.080 2.040 4.320 3.160 ;
        RECT  2.330 0.770 4.290 0.990 ;
        RECT  3.850 2.100 4.080 3.160 ;
        RECT  1.490 2.440 3.850 2.720 ;
        RECT  2.050 0.710 2.330 0.990 ;
        RECT  1.210 2.440 1.490 3.160 ;
        END
        ANTENNADIFFAREA 12.81 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.790 3.290 2.030 ;
        RECT  3.010 1.790 3.170 2.280 ;
        RECT  1.290 2.120 3.010 2.280 ;
        RECT  1.130 1.630 1.290 2.280 ;
        RECT  0.880 1.630 1.130 1.960 ;
        END
        ANTENNAGATEAREA 0.5904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.810 1.720 3.930 1.880 ;
        RECT  3.650 1.470 3.810 1.880 ;
        RECT  2.850 1.470 3.650 1.630 ;
        RECT  2.690 1.470 2.850 1.960 ;
        RECT  2.570 1.660 2.690 1.960 ;
        RECT  1.960 1.800 2.570 1.960 ;
        RECT  1.450 1.640 1.960 1.960 ;
        END
        ANTENNAGATEAREA 0.5904 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.720 1.680 ;
        END
        ANTENNAGATEAREA 0.2472 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.280 4.800 0.280 ;
        RECT  3.170 -0.280 3.450 0.610 ;
        RECT  1.170 -0.280 3.170 0.280 ;
        RECT  0.090 -0.280 1.170 0.290 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.650 3.320 4.800 3.880 ;
        RECT  3.370 2.930 3.650 3.880 ;
        RECT  1.970 3.260 3.370 3.880 ;
        RECT  1.690 2.930 1.970 3.880 ;
        RECT  0.960 3.320 1.690 3.880 ;
        RECT  0.680 2.120 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.130 1.340 4.310 1.620 ;
        RECT  4.090 1.150 4.130 1.620 ;
        RECT  3.970 1.150 4.090 1.560 ;
        RECT  2.400 1.150 3.970 1.310 ;
        RECT  2.120 1.150 2.400 1.620 ;
        RECT  1.480 1.150 2.120 1.310 ;
        RECT  1.320 0.920 1.480 1.310 ;
        RECT  0.770 0.920 1.320 1.080 ;
        RECT  0.490 0.840 0.770 1.080 ;
        RECT  0.280 0.920 0.490 1.080 ;
        RECT  0.280 1.960 0.440 3.160 ;
        RECT  0.120 0.920 0.280 3.160 ;
    END
END NAND3BX4TR

MACRO NAND3BX2TR
    CLASS CORE ;
    FOREIGN NAND3BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.240 3.120 2.360 ;
        RECT  2.880 1.000 3.040 2.810 ;
        RECT  1.930 1.000 2.880 1.160 ;
        RECT  2.250 2.650 2.880 2.810 ;
        RECT  1.970 2.650 2.250 2.930 ;
        RECT  1.290 2.650 1.970 2.810 ;
        RECT  1.650 0.880 1.930 1.160 ;
        RECT  1.010 2.650 1.290 2.930 ;
        END
        ANTENNADIFFAREA 5.028 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 2.260 2.690 2.420 ;
        RECT  0.950 1.950 1.120 2.420 ;
        RECT  0.900 1.580 0.950 2.420 ;
        RECT  0.880 1.580 0.900 2.410 ;
        RECT  0.790 1.580 0.880 2.190 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.790 2.440 1.960 ;
        RECT  1.280 1.640 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.440 0.720 2.880 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.280 3.200 0.280 ;
        RECT  2.810 -0.280 3.110 0.650 ;
        RECT  0.770 -0.280 2.810 0.280 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 3.320 3.200 3.880 ;
        RECT  1.490 2.970 1.770 3.880 ;
        RECT  0.770 3.320 1.490 3.880 ;
        RECT  0.490 3.180 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.730 1.320 2.050 1.630 ;
        RECT  1.330 1.320 1.730 1.480 ;
        RECT  1.170 1.260 1.330 1.480 ;
        RECT  0.370 1.260 1.170 1.420 ;
        RECT  0.090 1.020 0.370 2.190 ;
    END
END NAND3BX2TR

MACRO NAND3BX1TR
    CLASS CORE ;
    FOREIGN NAND3BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.440 2.320 2.720 ;
        RECT  2.080 0.440 2.150 1.560 ;
        RECT  1.090 2.440 2.150 2.720 ;
        RECT  1.850 0.790 2.080 1.070 ;
        END
        ANTENNADIFFAREA 3.328 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.910 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.510 1.590 1.960 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.550 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.280 2.400 0.280 ;
        RECT  0.690 -0.280 0.970 1.080 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 3.320 2.400 3.880 ;
        RECT  1.480 3.090 1.780 3.880 ;
        RECT  0.890 3.260 1.480 3.880 ;
        RECT  0.610 2.460 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.830 1.760 1.990 2.280 ;
        RECT  0.370 2.120 1.830 2.280 ;
        RECT  0.250 1.030 0.410 1.350 ;
        RECT  0.250 2.120 0.370 2.400 ;
        RECT  0.090 1.030 0.250 2.400 ;
    END
END NAND3BX1TR

MACRO NAND3XLTR
    CLASS CORE ;
    FOREIGN NAND3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.910 1.920 2.450 ;
        RECT  1.500 0.910 1.680 1.070 ;
        RECT  1.600 2.040 1.680 2.450 ;
        RECT  0.790 2.170 1.600 2.330 ;
        RECT  0.630 2.170 0.790 2.450 ;
        END
        ANTENNADIFFAREA 1.815 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.240 0.550 1.700 ;
        RECT  0.080 1.240 0.350 2.360 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.120 1.960 ;
        RECT  0.770 1.760 0.880 1.960 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.240 1.520 1.680 ;
        RECT  1.280 1.240 1.360 1.560 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 -0.280 2.000 0.280 ;
        RECT  0.200 -0.280 0.530 1.080 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 3.320 2.000 3.880 ;
        RECT  1.070 2.800 1.360 3.880 ;
        RECT  0.390 3.320 1.070 3.880 ;
        RECT  0.090 2.720 0.390 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END NAND3XLTR

MACRO NAND3X8TR
    CLASS CORE ;
    FOREIGN NAND3X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.140 0.480 8.620 2.960 ;
        RECT  1.660 0.480 8.140 0.960 ;
        RECT  7.880 2.240 8.140 2.960 ;
        RECT  7.540 2.350 7.880 2.960 ;
        RECT  7.260 2.350 7.540 3.160 ;
        RECT  6.580 2.350 7.260 2.820 ;
        RECT  6.300 2.350 6.580 3.160 ;
        RECT  5.540 2.350 6.300 2.820 ;
        RECT  5.260 2.350 5.540 3.160 ;
        RECT  4.420 2.350 5.260 2.820 ;
        RECT  4.140 2.350 4.420 3.160 ;
        RECT  3.460 2.350 4.140 2.830 ;
        RECT  3.180 2.350 3.460 3.160 ;
        RECT  2.340 2.520 3.180 3.000 ;
        RECT  2.060 2.520 2.340 3.160 ;
        RECT  1.300 2.520 2.060 3.000 ;
        RECT  1.020 2.520 1.300 3.160 ;
        END
        ANTENNADIFFAREA 19.16 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.720 1.330 7.980 1.610 ;
        RECT  7.700 1.330 7.720 2.190 ;
        RECT  7.560 1.450 7.700 2.190 ;
        RECT  5.740 2.030 7.560 2.190 ;
        RECT  4.980 1.910 5.740 2.190 ;
        RECT  2.820 2.030 4.980 2.190 ;
        RECT  2.740 1.950 2.820 2.350 ;
        RECT  2.480 1.950 2.740 2.360 ;
        RECT  1.020 2.200 2.480 2.360 ;
        RECT  0.860 1.910 1.020 2.360 ;
        RECT  0.740 1.910 0.860 2.190 ;
        END
        ANTENNAGATEAREA 1.2 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.120 1.570 7.400 1.850 ;
        RECT  6.300 1.690 7.120 1.850 ;
        RECT  6.020 1.590 6.300 1.870 ;
        RECT  4.780 1.590 6.020 1.750 ;
        RECT  4.620 1.590 4.780 1.870 ;
        RECT  3.250 1.690 4.620 1.870 ;
        RECT  2.980 1.550 3.250 1.870 ;
        RECT  2.320 1.550 2.980 1.710 ;
        RECT  2.080 1.550 2.320 2.000 ;
        RECT  1.220 1.780 2.080 2.000 ;
        END
        ANTENNAGATEAREA 1.2 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.540 1.130 6.870 1.530 ;
        RECT  4.140 1.130 6.540 1.290 ;
        RECT  3.860 1.130 4.140 1.530 ;
        RECT  1.920 1.130 3.860 1.290 ;
        RECT  1.620 1.130 1.920 1.590 ;
        END
        ANTENNAGATEAREA 1.2 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.020 -0.280 8.800 0.280 ;
        RECT  7.740 -0.280 8.020 0.320 ;
        RECT  5.580 -0.280 7.740 0.280 ;
        RECT  5.300 -0.280 5.580 0.320 ;
        RECT  3.180 -0.280 5.300 0.280 ;
        RECT  2.900 -0.280 3.180 0.320 ;
        RECT  0.780 -0.280 2.900 0.280 ;
        RECT  0.500 -0.280 0.780 1.260 ;
        RECT  0.000 -0.280 0.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.060 3.320 8.800 3.880 ;
        RECT  7.780 3.200 8.060 3.880 ;
        RECT  7.060 3.320 7.780 3.880 ;
        RECT  6.780 2.980 7.060 3.880 ;
        RECT  6.060 3.320 6.780 3.880 ;
        RECT  5.780 3.200 6.060 3.880 ;
        RECT  5.020 3.320 5.780 3.880 ;
        RECT  4.740 3.200 5.020 3.880 ;
        RECT  3.940 3.320 4.740 3.880 ;
        RECT  3.660 2.990 3.940 3.880 ;
        RECT  2.940 3.320 3.660 3.880 ;
        RECT  2.660 3.200 2.940 3.880 ;
        RECT  1.820 3.320 2.660 3.880 ;
        RECT  1.540 3.200 1.820 3.880 ;
        RECT  0.780 3.320 1.540 3.880 ;
        RECT  0.500 2.520 0.780 3.880 ;
        RECT  0.000 3.320 0.500 3.880 ;
        END
    END VDD
END NAND3X8TR

MACRO NAND3X6TR
    CLASS CORE ;
    FOREIGN NAND3X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.380 0.500 5.720 2.960 ;
        RECT  5.360 0.500 5.380 3.090 ;
        RECT  3.970 0.500 5.360 0.860 ;
        RECT  5.080 2.190 5.360 3.090 ;
        RECT  4.340 2.480 5.080 2.840 ;
        RECT  4.060 2.480 4.340 3.150 ;
        RECT  3.380 2.480 4.060 2.840 ;
        RECT  3.640 0.500 3.970 1.180 ;
        RECT  1.260 0.500 3.640 0.860 ;
        RECT  3.100 2.480 3.380 3.150 ;
        RECT  2.100 2.480 3.100 2.840 ;
        RECT  1.820 2.480 2.100 3.150 ;
        RECT  0.900 2.480 1.820 2.840 ;
        RECT  0.620 2.480 0.900 3.150 ;
        END
        ANTENNADIFFAREA 16.672 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.120 1.560 ;
        RECT  4.790 1.320 4.880 1.560 ;
        RECT  4.630 1.320 4.790 2.310 ;
        RECT  2.590 2.150 4.630 2.310 ;
        RECT  2.310 1.680 2.590 2.310 ;
        RECT  0.570 2.150 2.310 2.310 ;
        RECT  0.410 1.570 0.570 2.310 ;
        RECT  0.340 1.570 0.410 1.870 ;
        END
        ANTENNAGATEAREA 0.8832 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.040 1.640 4.460 1.980 ;
        RECT  3.160 1.820 4.040 1.980 ;
        RECT  3.080 1.570 3.160 1.980 ;
        RECT  2.920 1.360 3.080 1.980 ;
        RECT  2.140 1.360 2.920 1.520 ;
        RECT  1.970 1.360 2.140 1.920 ;
        RECT  1.880 1.590 1.970 1.920 ;
        RECT  0.970 1.720 1.880 1.920 ;
        RECT  0.780 1.620 0.970 1.920 ;
        END
        ANTENNAGATEAREA 0.8832 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 1.430 3.800 1.660 ;
        RECT  3.320 1.040 3.480 1.660 ;
        RECT  1.670 1.040 3.320 1.200 ;
        RECT  1.220 1.040 1.670 1.560 ;
        END
        ANTENNAGATEAREA 0.8832 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.020 -0.280 6.000 0.280 ;
        RECT  4.740 -0.280 5.020 0.340 ;
        RECT  2.700 -0.280 4.740 0.280 ;
        RECT  2.420 -0.280 2.700 0.340 ;
        RECT  0.380 -0.280 2.420 0.280 ;
        RECT  0.100 -0.280 0.380 1.250 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.860 3.320 6.000 3.880 ;
        RECT  4.580 3.200 4.860 3.880 ;
        RECT  3.860 3.320 4.580 3.880 ;
        RECT  3.580 3.010 3.860 3.880 ;
        RECT  2.820 3.320 3.580 3.880 ;
        RECT  2.540 3.080 2.820 3.880 ;
        RECT  1.420 3.320 2.540 3.880 ;
        RECT  1.140 3.080 1.420 3.880 ;
        RECT  0.380 3.320 1.140 3.880 ;
        RECT  0.100 2.510 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
END NAND3X6TR

MACRO NAND3X4TR
    CLASS CORE ;
    FOREIGN NAND3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 0.840 4.320 2.250 ;
        RECT  3.900 0.840 4.080 1.080 ;
        RECT  3.600 2.010 4.080 2.250 ;
        RECT  3.620 0.480 3.900 1.080 ;
        RECT  1.220 0.480 3.620 0.720 ;
        RECT  3.280 2.010 3.600 3.160 ;
        RECT  2.640 2.010 3.280 2.250 ;
        RECT  2.400 2.010 2.640 2.720 ;
        RECT  0.860 2.430 2.400 2.720 ;
        RECT  0.580 2.430 0.860 3.160 ;
        END
        ANTENNADIFFAREA 13.81 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.650 2.520 1.820 ;
        RECT  2.080 1.650 2.240 2.270 ;
        RECT  0.580 2.110 2.080 2.270 ;
        RECT  0.320 1.640 0.580 2.270 ;
        RECT  0.080 1.190 0.320 2.410 ;
        END
        ANTENNAGATEAREA 0.6072 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.670 3.310 1.850 ;
        RECT  2.690 1.280 2.850 1.850 ;
        RECT  1.920 1.280 2.690 1.440 ;
        RECT  1.730 1.280 1.920 1.950 ;
        RECT  1.120 1.790 1.730 1.950 ;
        RECT  0.850 1.240 1.120 1.950 ;
        RECT  0.790 1.670 0.850 1.950 ;
        END
        ANTENNAGATEAREA 0.6072 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.240 3.920 1.610 ;
        RECT  3.200 1.240 3.520 1.410 ;
        RECT  3.040 0.960 3.200 1.410 ;
        RECT  1.520 0.960 3.040 1.120 ;
        RECT  1.330 0.960 1.520 1.630 ;
        END
        ANTENNAGATEAREA 0.6072 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.660 -0.280 4.400 0.280 ;
        RECT  2.380 -0.280 2.660 0.320 ;
        RECT  0.380 -0.280 2.380 0.280 ;
        RECT  0.100 -0.280 0.380 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.120 3.320 4.400 3.880 ;
        RECT  3.840 2.410 4.120 3.880 ;
        RECT  3.080 3.320 3.840 3.880 ;
        RECT  2.800 2.410 3.080 3.880 ;
        RECT  1.340 3.260 2.800 3.880 ;
        RECT  1.060 2.930 1.340 3.880 ;
        RECT  0.380 3.320 1.060 3.880 ;
        RECT  0.100 2.570 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
END NAND3X4TR

MACRO NAND3X2TR
    CLASS CORE ;
    FOREIGN NAND3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.220 1.960 2.780 ;
        RECT  0.960 2.220 1.680 2.400 ;
        RECT  0.680 0.870 1.570 1.080 ;
        RECT  0.920 2.220 0.960 2.780 ;
        RECT  0.680 2.060 0.920 2.780 ;
        RECT  0.640 0.870 0.680 2.780 ;
        RECT  0.500 0.870 0.640 2.280 ;
        END
        ANTENNADIFFAREA 5.526 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.360 2.440 3.100 ;
        RECT  0.320 2.940 2.280 3.100 ;
        RECT  0.160 1.240 0.320 3.100 ;
        RECT  0.080 1.240 0.160 2.360 ;
        END
        ANTENNAGATEAREA 0.3096 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.750 2.110 2.040 ;
        RECT  1.920 1.240 2.080 2.040 ;
        RECT  1.120 1.240 1.920 1.400 ;
        RECT  1.070 1.240 1.120 1.560 ;
        RECT  0.840 1.240 1.070 1.900 ;
        END
        ANTENNAGATEAREA 0.3096 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.560 1.620 1.840 ;
        RECT  1.280 1.560 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.3096 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 -0.280 2.800 0.280 ;
        RECT  2.390 -0.280 2.680 1.070 ;
        RECT  0.400 -0.280 2.390 0.340 ;
        RECT  0.340 -0.280 0.400 0.560 ;
        RECT  0.120 -0.280 0.340 0.800 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 3.320 2.800 3.880 ;
        RECT  1.160 3.260 1.440 3.880 ;
        RECT  0.400 3.320 1.160 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND3X2TR

MACRO NAND3X1TR
    CLASS CORE ;
    FOREIGN NAND3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.740 1.920 3.160 ;
        RECT  1.480 0.740 1.760 1.020 ;
        RECT  1.680 2.040 1.760 3.160 ;
        RECT  0.590 2.320 1.680 2.540 ;
        END
        ANTENNADIFFAREA 3.328 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.380 0.680 1.660 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.720 1.160 2.000 ;
        RECT  0.880 1.600 1.120 2.000 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.470 1.600 1.750 ;
        RECT  1.320 1.240 1.520 1.750 ;
        RECT  1.280 1.240 1.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.640 -0.280 2.000 0.280 ;
        RECT  0.360 -0.280 0.640 0.990 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 3.320 2.000 3.880 ;
        RECT  0.120 3.010 1.410 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND3X1TR

MACRO NAND2BXLTR
    CLASS CORE ;
    FOREIGN NAND2BXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.440 1.920 2.610 ;
        RECT  1.640 0.440 1.760 1.560 ;
        RECT  1.390 2.450 1.760 2.610 ;
        RECT  1.080 2.450 1.390 2.680 ;
        END
        ANTENNADIFFAREA 0.64 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.160 1.920 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.520 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 -0.280 2.000 0.280 ;
        RECT  0.740 -0.280 1.020 0.760 ;
        RECT  0.000 -0.280 0.740 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.620 2.770 1.910 3.880 ;
        RECT  0.900 3.320 1.620 3.880 ;
        RECT  0.620 2.440 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.720 1.600 1.990 ;
        RECT  1.320 0.920 1.480 2.280 ;
        RECT  0.480 0.920 1.320 1.080 ;
        RECT  0.390 2.120 1.320 2.280 ;
        RECT  0.200 0.920 0.480 1.250 ;
        RECT  0.090 2.120 0.390 2.540 ;
    END
END NAND2BXLTR

MACRO NAND2BX4TR
    CLASS CORE ;
    FOREIGN NAND2BX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.530 0.980 3.770 2.380 ;
        RECT  1.900 0.980 3.530 1.220 ;
        RECT  3.520 2.140 3.530 2.380 ;
        RECT  3.280 2.140 3.520 2.960 ;
        RECT  2.540 2.140 3.280 2.380 ;
        RECT  2.270 2.140 2.540 3.160 ;
        RECT  1.560 2.140 2.270 2.380 ;
        RECT  1.680 0.520 1.900 1.220 ;
        RECT  1.320 2.140 1.560 3.160 ;
        END
        ANTENNADIFFAREA 7.329 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.380 2.820 1.600 ;
        RECT  1.520 1.380 2.520 1.560 ;
        RECT  1.280 1.240 1.520 1.560 ;
        RECT  1.240 1.380 1.280 1.560 ;
        RECT  1.080 1.380 1.240 1.660 ;
        END
        ANTENNAGATEAREA 0.588 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.24 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.280 4.000 0.280 ;
        RECT  2.420 -0.280 2.710 0.820 ;
        RECT  1.100 -0.280 2.420 0.280 ;
        RECT  0.820 -0.280 1.100 1.140 ;
        RECT  0.000 -0.280 0.820 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.020 3.320 4.000 3.880 ;
        RECT  2.720 2.550 3.020 3.880 ;
        RECT  2.060 3.320 2.720 3.880 ;
        RECT  1.770 2.540 2.060 3.880 ;
        RECT  1.100 3.320 1.770 3.880 ;
        RECT  0.810 2.450 1.100 3.880 ;
        RECT  0.000 3.320 0.810 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.060 1.800 3.370 1.980 ;
        RECT  2.160 1.820 3.060 1.980 ;
        RECT  1.430 1.720 2.160 1.980 ;
        RECT  1.040 1.820 1.430 1.980 ;
        RECT  0.880 1.820 1.040 2.290 ;
        RECT  0.640 2.120 0.880 2.290 ;
        RECT  0.340 2.120 0.640 2.840 ;
        RECT  0.340 0.520 0.620 1.310 ;
        RECT  0.280 1.150 0.340 1.310 ;
        RECT  0.280 2.120 0.340 2.290 ;
        RECT  0.120 1.150 0.280 2.290 ;
    END
END NAND2BX4TR

MACRO NAND2BX2TR
    CLASS CORE ;
    FOREIGN NAND2BX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        RECT  2.320 1.240 2.480 1.400 ;
        RECT  1.580 2.200 2.480 2.360 ;
        RECT  2.160 0.980 2.320 1.400 ;
        RECT  1.900 0.980 2.160 1.140 ;
        RECT  1.620 0.860 1.900 1.140 ;
        RECT  1.300 2.200 1.580 3.160 ;
        END
        ANTENNADIFFAREA 3.348 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.760 2.290 2.040 ;
        RECT  1.560 1.880 2.070 2.040 ;
        RECT  1.300 1.640 1.560 2.040 ;
        RECT  1.020 1.620 1.300 2.040 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.620 0.780 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 -0.280 2.800 0.280 ;
        RECT  2.480 -0.280 2.700 0.990 ;
        RECT  1.060 -0.280 2.480 0.280 ;
        RECT  0.780 -0.280 1.060 1.030 ;
        RECT  0.000 -0.280 0.780 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.100 3.320 2.800 3.880 ;
        RECT  1.820 2.560 2.100 3.880 ;
        RECT  1.060 3.320 1.820 3.880 ;
        RECT  0.780 2.440 1.060 3.880 ;
        RECT  0.000 3.320 0.780 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 1.300 2.000 1.580 ;
        RECT  0.540 1.300 1.720 1.460 ;
        RECT  0.320 1.030 0.540 1.460 ;
        RECT  0.320 2.120 0.540 2.400 ;
        RECT  0.260 1.030 0.320 2.400 ;
        RECT  0.160 1.300 0.260 2.400 ;
    END
END NAND2BX2TR

MACRO NAND2BX1TR
    CLASS CORE ;
    FOREIGN NAND2BX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.440 1.920 2.610 ;
        RECT  1.680 0.440 1.760 1.560 ;
        RECT  1.390 2.450 1.760 2.610 ;
        RECT  1.640 0.840 1.680 1.160 ;
        RECT  1.080 2.450 1.390 2.680 ;
        END
        ANTENNADIFFAREA 2.112 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.160 1.920 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.520 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 -0.280 2.000 0.280 ;
        RECT  0.740 -0.280 1.020 0.400 ;
        RECT  0.000 -0.280 0.740 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.620 2.770 1.910 3.880 ;
        RECT  0.900 3.320 1.620 3.880 ;
        RECT  0.620 2.440 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.720 1.600 1.990 ;
        RECT  1.320 0.920 1.480 2.280 ;
        RECT  0.480 0.920 1.320 1.080 ;
        RECT  0.390 2.120 1.320 2.280 ;
        RECT  0.200 0.920 0.480 1.250 ;
        RECT  0.090 2.100 0.390 2.320 ;
    END
END NAND2BX1TR

MACRO NAND2XLTR
    CLASS CORE ;
    FOREIGN NAND2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.800 1.240 1.080 ;
        RECT  0.690 0.920 0.930 1.080 ;
        RECT  0.690 2.040 0.920 2.410 ;
        RECT  0.530 0.920 0.690 2.410 ;
        RECT  0.480 2.040 0.530 2.410 ;
        END
        ANTENNADIFFAREA 0.64 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.530 0.370 1.810 ;
        RECT  0.080 1.530 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.240 1.160 1.660 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.370 -0.280 1.600 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 3.320 1.600 3.880 ;
        RECT  1.180 2.030 1.440 3.880 ;
        RECT  0.380 3.260 1.180 3.880 ;
        RECT  0.140 2.920 0.380 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
END NAND2XLTR

MACRO NAND2X8TR
    CLASS CORE ;
    FOREIGN NAND2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.770 1.840 4.920 2.590 ;
        RECT  4.280 0.500 4.770 2.590 ;
        RECT  4.250 0.500 4.280 1.080 ;
        RECT  3.890 2.110 4.280 2.590 ;
        RECT  2.850 0.600 4.250 1.080 ;
        RECT  3.610 2.110 3.890 3.160 ;
        RECT  2.850 2.110 3.610 2.590 ;
        RECT  2.570 0.440 2.850 1.080 ;
        RECT  2.570 2.110 2.850 3.160 ;
        RECT  1.170 0.590 2.570 1.080 ;
        RECT  1.810 2.110 2.570 2.590 ;
        RECT  1.530 2.110 1.810 3.160 ;
        RECT  0.850 2.110 1.530 2.580 ;
        RECT  0.890 0.440 1.170 1.080 ;
        RECT  0.570 2.110 0.850 3.160 ;
        END
        ANTENNADIFFAREA 13.772 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.560 3.480 1.950 ;
        RECT  2.170 1.790 3.200 1.950 ;
        RECT  1.890 1.560 2.170 1.950 ;
        RECT  0.570 1.790 1.890 1.950 ;
        RECT  0.320 1.630 0.570 1.950 ;
        RECT  0.080 1.190 0.320 2.410 ;
        END
        ANTENNAGATEAREA 1.1088 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.670 4.120 1.950 ;
        RECT  3.800 1.240 3.960 1.950 ;
        RECT  3.640 1.240 3.800 1.560 ;
        RECT  3.040 1.240 3.640 1.400 ;
        RECT  2.760 1.240 3.040 1.630 ;
        RECT  1.370 1.240 2.760 1.400 ;
        RECT  1.210 1.240 1.370 1.610 ;
        RECT  0.730 1.380 1.210 1.610 ;
        END
        ANTENNAGATEAREA 1.1088 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 -0.280 5.200 0.280 ;
        RECT  3.410 -0.280 3.690 0.400 ;
        RECT  2.010 -0.280 3.410 0.280 ;
        RECT  1.730 -0.280 2.010 0.400 ;
        RECT  0.370 -0.280 1.730 0.280 ;
        RECT  0.090 -0.280 0.370 0.690 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.410 3.320 5.200 3.880 ;
        RECT  4.130 2.800 4.410 3.880 ;
        RECT  3.370 3.320 4.130 3.880 ;
        RECT  3.090 2.810 3.370 3.880 ;
        RECT  2.370 3.320 3.090 3.880 ;
        RECT  2.090 2.910 2.370 3.880 ;
        RECT  1.330 3.320 2.090 3.880 ;
        RECT  1.050 2.940 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.910 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END NAND2X8TR

MACRO NAND2X6TR
    CLASS CORE ;
    FOREIGN NAND2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.590 0.840 3.910 2.410 ;
        RECT  2.870 0.840 3.590 1.200 ;
        RECT  3.320 2.050 3.590 2.410 ;
        RECT  2.800 2.050 3.320 2.960 ;
        RECT  2.600 0.440 2.870 1.200 ;
        RECT  2.460 2.050 2.800 3.160 ;
        RECT  2.590 0.440 2.600 1.080 ;
        RECT  1.190 0.720 2.590 1.080 ;
        RECT  1.830 2.050 2.460 2.410 ;
        RECT  1.550 2.050 1.830 3.160 ;
        RECT  0.870 2.050 1.550 2.410 ;
        RECT  0.910 0.440 1.190 1.080 ;
        RECT  0.590 2.050 0.870 3.160 ;
        END
        ANTENNADIFFAREA 10.52 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.420 3.410 1.890 ;
        RECT  2.110 1.730 3.250 1.890 ;
        RECT  1.830 1.560 2.110 1.890 ;
        RECT  0.530 1.730 1.830 1.890 ;
        RECT  0.350 1.270 0.530 1.890 ;
        RECT  0.330 0.790 0.350 1.890 ;
        RECT  0.080 0.790 0.330 2.010 ;
        END
        ANTENNAGATEAREA 0.8736 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.360 3.030 1.520 ;
        RECT  2.270 1.240 2.430 1.520 ;
        RECT  1.230 1.240 2.270 1.400 ;
        RECT  0.820 1.240 1.230 1.570 ;
        END
        ANTENNAGATEAREA 0.8736 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.880 -0.280 4.000 0.280 ;
        RECT  3.600 -0.280 3.880 0.680 ;
        RECT  2.030 -0.280 3.600 0.280 ;
        RECT  1.750 -0.280 2.030 0.400 ;
        RECT  0.390 -0.280 1.750 0.280 ;
        RECT  0.100 -0.280 0.390 0.630 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 3.320 4.000 3.880 ;
        RECT  3.130 3.120 3.400 3.880 ;
        RECT  2.300 3.320 3.130 3.880 ;
        RECT  2.030 2.570 2.300 3.880 ;
        RECT  1.350 3.320 2.030 3.880 ;
        RECT  1.070 2.570 1.350 3.880 ;
        RECT  0.400 3.320 1.070 3.880 ;
        RECT  0.110 2.390 0.400 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
END NAND2X6TR

MACRO NAND2X4TR
    CLASS CORE ;
    FOREIGN NAND2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.440 3.120 2.360 ;
        RECT  2.710 0.440 2.880 1.360 ;
        RECT  2.600 2.120 2.880 2.360 ;
        RECT  2.480 0.640 2.710 1.360 ;
        RECT  2.320 2.120 2.600 3.160 ;
        RECT  1.040 0.650 2.480 0.930 ;
        RECT  1.640 2.120 2.320 2.360 ;
        RECT  1.360 2.120 1.640 3.160 ;
        END
        ANTENNADIFFAREA 7.362 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.360 2.320 1.640 ;
        RECT  1.640 1.090 1.800 1.640 ;
        RECT  0.720 1.090 1.640 1.250 ;
        RECT  0.370 1.090 0.720 1.700 ;
        END
        ANTENNAGATEAREA 0.5928 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.540 2.720 1.960 ;
        RECT  1.360 1.800 2.520 1.960 ;
        RECT  0.880 1.410 1.360 1.960 ;
        END
        ANTENNAGATEAREA 0.5928 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 -0.280 3.200 0.280 ;
        RECT  1.880 -0.280 2.160 0.400 ;
        RECT  0.540 -0.280 1.880 0.280 ;
        RECT  0.240 -0.280 0.540 0.930 ;
        RECT  0.000 -0.280 0.240 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.080 3.320 3.200 3.880 ;
        RECT  2.800 2.580 3.080 3.880 ;
        RECT  2.120 3.320 2.800 3.880 ;
        RECT  1.840 2.590 2.120 3.880 ;
        RECT  1.120 3.320 1.840 3.880 ;
        RECT  0.870 3.200 1.120 3.880 ;
        RECT  0.590 2.270 0.870 3.880 ;
        RECT  0.000 3.320 0.590 3.880 ;
        END
    END VDD
END NAND2X4TR

MACRO NAND2X2TR
    CLASS CORE ;
    FOREIGN NAND2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.000 1.920 2.240 ;
        RECT  1.520 1.000 1.760 1.160 ;
        RECT  1.390 2.080 1.760 2.240 ;
        RECT  1.280 0.840 1.520 1.160 ;
        RECT  1.110 2.080 1.390 3.160 ;
        RECT  1.130 0.840 1.280 1.000 ;
        RECT  0.830 0.720 1.130 1.000 ;
        END
        ANTENNADIFFAREA 3.348 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.620 1.600 1.920 ;
        RECT  0.460 1.760 1.380 1.920 ;
        RECT  0.320 1.320 0.460 1.920 ;
        RECT  0.080 0.830 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.240 1.120 1.600 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.630 2.400 1.910 3.880 ;
        RECT  0.870 3.320 1.630 3.880 ;
        RECT  0.590 2.080 0.870 3.880 ;
        RECT  0.000 3.320 0.590 3.880 ;
        END
    END VDD
END NAND2X2TR

MACRO NAND2X1TR
    CLASS CORE ;
    FOREIGN NAND2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 0.800 1.240 1.080 ;
        RECT  0.690 2.040 0.920 2.410 ;
        RECT  0.530 0.800 0.690 2.410 ;
        RECT  0.480 2.040 0.530 2.410 ;
        END
        ANTENNADIFFAREA 2.112 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.370 1.810 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.240 1.160 1.730 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.370 -0.280 1.600 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 3.320 1.600 3.880 ;
        RECT  1.160 2.030 1.440 3.880 ;
        RECT  0.400 3.260 1.160 3.880 ;
        RECT  0.120 2.570 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END NAND2X1TR

MACRO MXI4XLTR
    CLASS CORE ;
    FOREIGN MXI4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.940 0.450 9.120 3.160 ;
        RECT  8.730 0.450 8.940 0.610 ;
        RECT  8.830 2.040 8.940 3.160 ;
        END
        ANTENNADIFFAREA 1.188 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.240 7.920 1.750 ;
        RECT  7.560 1.470 7.680 1.750 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.150 2.720 1.560 ;
        RECT  2.320 1.150 2.480 1.430 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.240 3.520 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.580 5.240 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 1.590 2.320 1.960 ;
        RECT  2.040 1.470 2.150 1.960 ;
        RECT  1.870 1.470 2.040 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.520 -0.280 9.200 0.280 ;
        RECT  7.800 -0.280 8.520 0.610 ;
        RECT  5.450 -0.280 7.800 0.340 ;
        RECT  5.170 -0.280 5.450 0.460 ;
        RECT  3.310 -0.280 5.170 0.400 ;
        RECT  3.030 -0.280 3.310 1.080 ;
        RECT  2.270 -0.280 3.030 0.340 ;
        RECT  1.990 -0.280 2.270 0.610 ;
        RECT  0.370 -0.280 1.990 0.280 ;
        RECT  0.090 -0.280 0.370 0.860 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.620 3.320 9.200 3.880 ;
        RECT  8.340 2.700 8.620 3.880 ;
        RECT  8.080 3.320 8.340 3.880 ;
        RECT  7.800 3.260 8.080 3.880 ;
        RECT  5.450 3.320 7.800 3.880 ;
        RECT  5.170 3.260 5.450 3.880 ;
        RECT  3.170 3.320 5.170 3.880 ;
        RECT  2.890 2.990 3.170 3.880 ;
        RECT  2.270 3.320 2.890 3.880 ;
        RECT  1.990 2.990 2.270 3.880 ;
        RECT  0.370 3.320 1.990 3.880 ;
        RECT  0.090 2.620 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.620 0.770 8.780 1.800 ;
        RECT  6.620 0.770 8.620 0.930 ;
        RECT  8.240 1.970 8.480 2.130 ;
        RECT  8.240 1.090 8.460 1.310 ;
        RECT  8.160 2.370 8.290 2.530 ;
        RECT  8.080 1.090 8.240 2.130 ;
        RECT  8.000 2.370 8.160 3.040 ;
        RECT  7.840 1.960 8.080 2.130 ;
        RECT  3.610 2.880 8.000 3.040 ;
        RECT  7.680 1.960 7.840 2.650 ;
        RECT  6.940 2.370 7.680 2.650 ;
        RECT  7.400 1.090 7.520 1.310 ;
        RECT  7.400 1.910 7.520 2.190 ;
        RECT  7.240 1.090 7.400 2.190 ;
        RECT  7.100 1.490 7.240 1.770 ;
        RECT  6.940 1.090 7.060 1.310 ;
        RECT  6.780 1.090 6.940 2.650 ;
        RECT  6.340 0.520 6.620 2.440 ;
        RECT  6.000 0.900 6.010 1.180 ;
        RECT  5.840 0.900 6.000 2.440 ;
        RECT  5.730 0.900 5.840 1.180 ;
        RECT  5.400 1.830 5.680 2.720 ;
        RECT  4.390 2.560 5.400 2.720 ;
        RECT  4.730 0.900 5.010 1.180 ;
        RECT  4.720 2.120 5.010 2.400 ;
        RECT  4.720 1.020 4.730 1.180 ;
        RECT  4.560 1.020 4.720 2.400 ;
        RECT  4.230 0.900 4.390 2.720 ;
        RECT  3.910 0.960 4.070 2.320 ;
        RECT  3.890 0.960 3.910 1.160 ;
        RECT  3.730 2.160 3.910 2.320 ;
        RECT  3.670 0.900 3.890 1.160 ;
        RECT  2.830 1.720 3.750 2.000 ;
        RECT  3.450 2.160 3.730 2.440 ;
        RECT  3.450 2.670 3.610 3.040 ;
        RECT  1.370 2.670 3.450 2.830 ;
        RECT  2.550 0.710 2.830 0.990 ;
        RECT  2.550 1.720 2.830 2.510 ;
        RECT  1.390 0.770 2.550 0.930 ;
        RECT  1.390 2.350 2.550 2.510 ;
        RECT  1.710 1.090 1.830 1.310 ;
        RECT  1.710 1.910 1.830 2.190 ;
        RECT  1.550 1.090 1.710 2.190 ;
        RECT  1.230 0.770 1.390 2.510 ;
        RECT  1.090 2.670 1.370 2.950 ;
        RECT  1.070 2.670 1.090 2.830 ;
        RECT  0.910 0.520 1.070 2.830 ;
        RECT  0.790 0.520 0.910 0.800 ;
        RECT  0.530 1.030 0.750 2.250 ;
    END
END MXI4XLTR

MACRO MXI4X4TR
    CLASS CORE ;
    FOREIGN MXI4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.290 0.450 9.530 3.150 ;
        RECT  9.150 0.450 9.290 1.240 ;
        RECT  9.150 1.840 9.290 3.150 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.580 1.580 7.920 1.960 ;
        END
        ANTENNAGATEAREA 0.3528 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.140 2.810 1.620 ;
        END
        ANTENNAGATEAREA 0.576 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.240 3.540 1.710 ;
        END
        ANTENNAGATEAREA 0.1896 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.220 1.620 5.520 1.960 ;
        END
        ANTENNAGATEAREA 0.2088 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.400 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1896 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.520 0.470 1.840 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.850 -0.280 10.000 0.280 ;
        RECT  9.690 -0.280 9.850 1.310 ;
        RECT  8.910 -0.280 9.690 0.280 ;
        RECT  8.630 -0.280 8.910 0.330 ;
        RECT  7.920 -0.280 8.630 0.280 ;
        RECT  7.640 -0.280 7.920 0.490 ;
        RECT  5.520 -0.280 7.640 0.280 ;
        RECT  5.360 -0.280 5.520 1.290 ;
        RECT  3.540 -0.280 5.360 0.280 ;
        RECT  3.260 -0.280 3.540 0.980 ;
        RECT  2.550 -0.280 3.260 0.280 ;
        RECT  2.270 -0.280 2.550 0.600 ;
        RECT  0.310 -0.280 2.270 0.280 ;
        RECT  0.150 -0.280 0.310 0.930 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.850 3.320 10.000 3.880 ;
        RECT  9.690 1.930 9.850 3.880 ;
        RECT  8.950 3.320 9.690 3.880 ;
        RECT  8.670 2.990 8.950 3.880 ;
        RECT  8.040 3.320 8.670 3.880 ;
        RECT  7.760 3.260 8.040 3.880 ;
        RECT  5.700 3.320 7.760 3.880 ;
        RECT  5.420 3.260 5.700 3.880 ;
        RECT  3.420 3.320 5.420 3.880 ;
        RECT  3.140 2.950 3.420 3.880 ;
        RECT  2.390 3.320 3.140 3.880 ;
        RECT  2.110 2.950 2.390 3.880 ;
        RECT  0.380 3.320 2.110 3.880 ;
        RECT  0.090 2.650 0.380 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.970 1.400 9.130 1.680 ;
        RECT  8.940 1.400 8.970 1.560 ;
        RECT  8.780 0.650 8.940 1.560 ;
        RECT  8.720 1.860 8.880 2.830 ;
        RECT  6.640 0.650 8.780 0.810 ;
        RECT  8.610 1.860 8.720 2.020 ;
        RECT  8.500 2.670 8.720 2.830 ;
        RECT  8.450 1.600 8.610 2.020 ;
        RECT  8.290 2.200 8.560 2.360 ;
        RECT  8.340 2.670 8.500 2.920 ;
        RECT  8.290 1.030 8.380 1.330 ;
        RECT  7.600 2.760 8.340 2.920 ;
        RECT  8.220 1.030 8.290 2.360 ;
        RECT  8.110 1.170 8.220 2.360 ;
        RECT  7.930 2.170 8.110 2.600 ;
        RECT  7.280 2.440 7.930 2.600 ;
        RECT  7.420 2.120 7.680 2.280 ;
        RECT  7.440 2.760 7.600 3.160 ;
        RECT  6.020 3.000 7.440 3.160 ;
        RECT  7.260 0.980 7.420 2.280 ;
        RECT  7.120 2.440 7.280 2.840 ;
        RECT  7.120 1.380 7.260 1.640 ;
        RECT  6.960 2.440 7.120 2.600 ;
        RECT  6.800 1.040 6.960 2.600 ;
        RECT  6.480 0.650 6.640 2.840 ;
        RECT  6.250 0.890 6.480 1.050 ;
        RECT  6.000 1.270 6.160 2.660 ;
        RECT  5.860 2.940 6.020 3.160 ;
        RECT  5.840 0.460 6.000 1.440 ;
        RECT  4.020 2.940 5.860 3.100 ;
        RECT  5.680 1.620 5.840 2.720 ;
        RECT  4.720 2.560 5.680 2.720 ;
        RECT  5.040 2.120 5.180 2.280 ;
        RECT  4.880 0.590 5.040 2.280 ;
        RECT  4.560 0.600 4.720 2.720 ;
        RECT  4.260 0.600 4.560 0.760 ;
        RECT  4.420 2.560 4.560 2.720 ;
        RECT  4.240 0.980 4.400 2.400 ;
        RECT  4.000 0.980 4.240 1.140 ;
        RECT  3.940 2.240 4.240 2.400 ;
        RECT  3.920 1.560 4.080 2.080 ;
        RECT  3.860 2.630 4.020 3.100 ;
        RECT  3.840 0.860 4.000 1.140 ;
        RECT  2.850 1.920 3.920 2.080 ;
        RECT  1.270 2.630 3.860 2.790 ;
        RECT  2.850 0.760 3.010 0.980 ;
        RECT  1.590 0.760 2.850 0.920 ;
        RECT  2.690 1.920 2.850 2.470 ;
        RECT  1.430 2.310 2.690 2.470 ;
        RECT  1.910 1.080 2.030 1.240 ;
        RECT  1.750 1.080 1.910 2.150 ;
        RECT  1.590 1.990 1.750 2.150 ;
        RECT  1.430 0.760 1.590 1.650 ;
        RECT  1.270 1.490 1.430 2.470 ;
        RECT  1.110 0.760 1.270 1.040 ;
        RECT  1.110 2.630 1.270 2.910 ;
        RECT  0.950 0.880 1.110 2.790 ;
        RECT  0.630 0.630 0.790 2.950 ;
    END
END MXI4X4TR

MACRO MXI4X2TR
    CLASS CORE ;
    FOREIGN MXI4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.480 0.440 9.520 2.100 ;
        RECT  9.280 0.440 9.480 3.160 ;
        RECT  9.200 0.440 9.280 1.300 ;
        RECT  9.200 1.940 9.280 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.580 1.580 7.920 1.960 ;
        END
        ANTENNAGATEAREA 0.2832 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.610 3.120 1.960 ;
        RECT  2.880 1.300 3.090 1.960 ;
        END
        ANTENNAGATEAREA 0.4584 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.260 3.580 1.570 ;
        RECT  3.280 1.090 3.520 1.570 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.340 1.170 5.560 1.560 ;
        RECT  5.230 1.240 5.340 1.560 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.210 2.720 1.660 ;
        RECT  2.350 1.500 2.480 1.660 ;
        RECT  2.130 1.500 2.350 1.780 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.610 0.450 1.930 ;
        RECT  0.080 1.320 0.320 2.280 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.960 -0.280 9.600 0.280 ;
        RECT  8.680 -0.280 8.960 0.400 ;
        RECT  7.960 -0.280 8.680 0.280 ;
        RECT  7.680 -0.280 7.960 0.400 ;
        RECT  5.580 -0.280 7.680 0.340 ;
        RECT  5.300 -0.280 5.580 0.870 ;
        RECT  3.590 -0.280 5.300 0.340 ;
        RECT  3.310 -0.280 3.590 0.930 ;
        RECT  2.610 -0.280 3.310 0.280 ;
        RECT  2.330 -0.280 2.610 0.580 ;
        RECT  0.370 -0.280 2.330 0.340 ;
        RECT  0.090 -0.280 0.370 1.040 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.000 3.320 9.600 3.880 ;
        RECT  8.720 2.930 9.000 3.880 ;
        RECT  7.960 3.320 8.720 3.880 ;
        RECT  7.680 3.200 7.960 3.880 ;
        RECT  5.620 3.260 7.680 3.880 ;
        RECT  5.340 3.200 5.620 3.880 ;
        RECT  3.410 3.260 5.340 3.880 ;
        RECT  3.130 3.020 3.410 3.880 ;
        RECT  2.430 3.320 3.130 3.880 ;
        RECT  2.150 3.020 2.430 3.880 ;
        RECT  0.370 3.260 2.150 3.880 ;
        RECT  0.090 2.540 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.000 1.460 9.120 1.740 ;
        RECT  8.960 0.650 9.000 1.740 ;
        RECT  8.840 0.650 8.960 1.620 ;
        RECT  6.620 0.650 8.840 0.810 ;
        RECT  8.680 1.780 8.800 2.770 ;
        RECT  8.640 1.660 8.680 2.770 ;
        RECT  8.400 1.660 8.640 1.940 ;
        RECT  8.560 2.610 8.640 2.770 ;
        RECT  8.400 2.610 8.560 3.040 ;
        RECT  8.240 0.990 8.480 1.270 ;
        RECT  8.240 2.100 8.480 2.450 ;
        RECT  3.730 2.880 8.400 3.040 ;
        RECT  8.200 0.990 8.240 2.720 ;
        RECT  8.080 1.110 8.200 2.720 ;
        RECT  7.100 2.560 8.080 2.720 ;
        RECT  7.420 0.970 7.560 1.250 ;
        RECT  7.420 2.120 7.560 2.400 ;
        RECT  7.260 0.970 7.420 2.400 ;
        RECT  7.100 1.450 7.260 1.730 ;
        RECT  6.940 1.010 7.100 1.290 ;
        RECT  6.940 2.290 7.100 2.720 ;
        RECT  6.820 1.010 6.940 2.720 ;
        RECT  6.780 1.130 6.820 2.720 ;
        RECT  6.340 0.650 6.620 2.570 ;
        RECT  6.020 0.590 6.180 2.630 ;
        RECT  5.860 0.590 6.020 1.310 ;
        RECT  5.860 2.220 6.020 2.630 ;
        RECT  5.390 1.720 5.860 2.000 ;
        RECT  5.230 1.720 5.390 2.720 ;
        RECT  4.630 2.560 5.230 2.720 ;
        RECT  4.790 0.860 5.070 2.400 ;
        RECT  4.470 0.770 4.630 2.720 ;
        RECT  4.270 0.770 4.470 1.050 ;
        RECT  4.130 2.440 4.470 2.720 ;
        RECT  4.150 1.210 4.310 2.280 ;
        RECT  4.070 1.210 4.150 1.370 ;
        RECT  3.930 2.120 4.150 2.280 ;
        RECT  3.910 0.860 4.070 1.370 ;
        RECT  3.770 1.610 3.990 1.960 ;
        RECT  3.710 2.120 3.930 2.400 ;
        RECT  3.790 0.860 3.910 1.140 ;
        RECT  3.550 1.800 3.770 1.960 ;
        RECT  3.570 2.700 3.730 3.040 ;
        RECT  1.370 2.700 3.570 2.860 ;
        RECT  3.390 1.800 3.550 2.520 ;
        RECT  1.470 2.360 3.390 2.520 ;
        RECT  2.850 0.760 3.070 1.040 ;
        RECT  1.650 0.760 2.850 0.920 ;
        RECT  1.970 1.080 2.090 1.300 ;
        RECT  1.810 1.080 1.970 2.200 ;
        RECT  1.630 2.040 1.810 2.200 ;
        RECT  1.490 0.760 1.650 1.780 ;
        RECT  1.470 1.500 1.490 1.780 ;
        RECT  1.310 1.500 1.470 2.520 ;
        RECT  1.150 2.700 1.370 2.920 ;
        RECT  1.150 0.800 1.330 1.080 ;
        RECT  1.050 0.800 1.150 2.920 ;
        RECT  0.990 0.920 1.050 2.920 ;
        RECT  0.610 1.030 0.830 2.920 ;
        RECT  0.570 1.030 0.610 1.310 ;
    END
END MXI4X2TR

MACRO MXI4X1TR
    CLASS CORE ;
    FOREIGN MXI4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.880 0.510 9.120 2.360 ;
        RECT  8.870 2.040 8.880 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.150 1.170 7.520 1.690 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.420 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2208 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.150 1.690 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.180 5.190 1.560 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.650 ;
        RECT  1.960 1.420 2.080 1.650 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.560 0.400 2.760 ;
        RECT  0.080 1.640 0.240 2.760 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.630 -0.280 9.200 0.280 ;
        RECT  8.350 -0.280 8.630 0.660 ;
        RECT  7.700 -0.280 8.350 0.280 ;
        RECT  7.480 -0.280 7.700 0.340 ;
        RECT  5.380 -0.280 7.480 0.280 ;
        RECT  5.100 -0.280 5.380 0.340 ;
        RECT  3.340 -0.280 5.100 0.280 ;
        RECT  3.060 -0.280 3.340 1.080 ;
        RECT  2.320 -0.280 3.060 0.280 ;
        RECT  2.040 -0.280 2.320 0.610 ;
        RECT  0.410 -0.280 2.040 0.280 ;
        RECT  0.150 -0.280 0.410 1.310 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 3.320 9.200 3.880 ;
        RECT  7.920 2.950 8.530 3.880 ;
        RECT  5.300 3.320 7.920 3.880 ;
        RECT  5.020 3.160 5.300 3.880 ;
        RECT  3.250 3.320 5.020 3.880 ;
        RECT  2.960 2.930 3.250 3.880 ;
        RECT  2.320 3.320 2.960 3.880 ;
        RECT  2.040 2.930 2.320 3.880 ;
        RECT  0.410 3.320 2.040 3.880 ;
        RECT  0.120 3.100 0.410 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.560 0.850 8.720 1.230 ;
        RECT  7.310 0.850 8.560 1.010 ;
        RECT  8.290 1.670 8.450 2.780 ;
        RECT  8.200 1.670 8.290 1.830 ;
        RECT  7.760 2.620 8.290 2.780 ;
        RECT  8.040 1.610 8.200 1.830 ;
        RECT  7.840 1.170 8.130 1.330 ;
        RECT  7.840 2.170 8.080 2.340 ;
        RECT  7.680 1.170 7.840 2.340 ;
        RECT  7.600 2.620 7.760 3.120 ;
        RECT  7.310 2.170 7.680 2.340 ;
        RECT  5.620 2.960 7.600 3.120 ;
        RECT  7.150 0.440 7.310 1.010 ;
        RECT  7.150 2.170 7.310 2.800 ;
        RECT  6.280 0.440 7.150 0.600 ;
        RECT  6.440 2.640 7.150 2.800 ;
        RECT  6.830 0.760 6.990 2.340 ;
        RECT  6.640 0.760 6.830 0.920 ;
        RECT  6.730 1.690 6.830 2.340 ;
        RECT  6.600 1.690 6.730 1.970 ;
        RECT  6.510 1.240 6.670 1.520 ;
        RECT  6.440 1.360 6.510 1.520 ;
        RECT  6.280 1.360 6.440 2.800 ;
        RECT  6.120 0.440 6.280 0.850 ;
        RECT  5.960 0.690 6.120 2.640 ;
        RECT  5.640 0.800 5.740 2.300 ;
        RECT  5.580 0.800 5.640 2.420 ;
        RECT  5.460 2.840 5.620 3.120 ;
        RECT  5.480 2.140 5.580 2.420 ;
        RECT  3.690 2.840 5.460 3.000 ;
        RECT  5.110 1.720 5.380 1.980 ;
        RECT  4.950 1.720 5.110 2.680 ;
        RECT  4.240 2.520 4.950 2.680 ;
        RECT  4.670 0.860 4.900 1.020 ;
        RECT  4.670 2.200 4.780 2.360 ;
        RECT  4.500 0.860 4.670 2.360 ;
        RECT  4.240 0.820 4.320 1.110 ;
        RECT  4.080 0.820 4.240 2.680 ;
        RECT  3.760 0.860 3.920 2.380 ;
        RECT  3.620 0.860 3.760 1.020 ;
        RECT  3.520 2.220 3.760 2.380 ;
        RECT  3.530 2.610 3.690 3.000 ;
        RECT  3.440 1.470 3.600 2.060 ;
        RECT  1.330 2.610 3.530 2.770 ;
        RECT  3.230 1.900 3.440 2.060 ;
        RECT  3.070 1.900 3.230 2.450 ;
        RECT  1.480 2.290 3.070 2.450 ;
        RECT  2.660 0.770 2.820 1.060 ;
        RECT  1.480 0.770 2.660 0.930 ;
        RECT  1.800 1.090 1.920 1.250 ;
        RECT  1.800 1.910 1.890 2.130 ;
        RECT  1.640 1.090 1.800 2.130 ;
        RECT  1.320 0.770 1.480 2.450 ;
        RECT  1.170 2.610 1.330 2.890 ;
        RECT  1.160 2.610 1.170 2.770 ;
        RECT  1.000 0.440 1.160 2.770 ;
        RECT  0.680 1.030 0.840 2.450 ;
        RECT  0.630 2.170 0.680 2.450 ;
    END
END MXI4X1TR

MACRO MXI3XLTR
    CLASS CORE ;
    FOREIGN MXI3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 0.440 7.120 2.860 ;
        RECT  6.890 0.440 6.960 0.720 ;
        RECT  6.880 1.640 6.960 2.860 ;
        RECT  6.800 2.580 6.880 2.860 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.640 6.480 1.960 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 2.840 1.160 3.160 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.560 3.520 1.960 ;
        RECT  3.160 1.560 3.240 1.840 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.400 1.640 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.400 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.550 -0.280 7.200 0.280 ;
        RECT  6.270 -0.280 6.550 0.400 ;
        RECT  5.720 -0.280 6.270 0.280 ;
        RECT  5.560 -0.280 5.720 0.840 ;
        RECT  3.620 -0.280 5.560 0.340 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  2.440 -0.280 3.340 0.280 ;
        RECT  2.160 -0.280 2.440 1.080 ;
        RECT  0.370 -0.280 2.160 0.280 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.600 3.320 7.200 3.880 ;
        RECT  6.320 2.690 6.600 3.880 ;
        RECT  5.980 3.320 6.320 3.880 ;
        RECT  5.760 2.560 5.980 3.880 ;
        RECT  2.340 3.260 5.760 3.880 ;
        RECT  2.060 2.940 2.340 3.880 ;
        RECT  0.370 3.320 2.060 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.680 0.870 6.800 1.150 ;
        RECT  6.520 0.580 6.680 1.150 ;
        RECT  5.920 2.120 6.540 2.400 ;
        RECT  6.040 0.580 6.520 0.740 ;
        RECT  6.200 0.900 6.360 1.480 ;
        RECT  5.920 1.320 6.200 1.480 ;
        RECT  5.880 0.580 6.040 1.160 ;
        RECT  5.760 1.320 5.920 2.400 ;
        RECT  5.400 1.000 5.880 1.160 ;
        RECT  5.360 1.490 5.760 1.650 ;
        RECT  5.380 1.990 5.600 3.100 ;
        RECT  5.240 0.500 5.400 1.160 ;
        RECT  2.660 2.940 5.380 3.100 ;
        RECT  5.080 1.490 5.360 1.770 ;
        RECT  4.600 0.500 5.240 0.660 ;
        RECT  5.000 1.930 5.220 2.600 ;
        RECT  4.920 0.820 5.080 1.100 ;
        RECT  4.920 1.930 5.000 2.090 ;
        RECT  4.760 0.820 4.920 2.090 ;
        RECT  4.600 2.250 4.800 2.530 ;
        RECT  4.440 0.500 4.600 2.530 ;
        RECT  4.380 0.780 4.440 1.060 ;
        RECT  4.220 1.910 4.280 2.720 ;
        RECT  4.120 0.920 4.220 2.720 ;
        RECT  4.060 0.800 4.120 2.720 ;
        RECT  3.840 0.800 4.060 1.080 ;
        RECT  3.680 1.240 3.900 2.780 ;
        RECT  3.320 1.240 3.680 1.400 ;
        RECT  3.080 2.500 3.680 2.780 ;
        RECT  3.160 0.690 3.320 1.400 ;
        RECT  3.060 0.690 3.160 0.850 ;
        RECT  2.780 0.570 3.060 0.850 ;
        RECT  2.900 1.030 3.000 1.860 ;
        RECT  2.720 1.030 2.900 2.460 ;
        RECT  2.620 1.800 2.720 2.460 ;
        RECT  2.500 2.620 2.660 3.100 ;
        RECT  1.920 1.800 2.620 1.960 ;
        RECT  1.480 2.620 2.500 2.780 ;
        RECT  1.700 1.680 1.920 1.960 ;
        RECT  1.620 2.120 1.900 2.340 ;
        RECT  1.600 1.010 1.880 1.320 ;
        RECT  1.540 2.120 1.620 2.280 ;
        RECT  1.540 1.160 1.600 1.320 ;
        RECT  1.380 1.160 1.540 2.280 ;
        RECT  1.340 0.440 1.480 0.660 ;
        RECT  1.320 2.440 1.480 2.780 ;
        RECT  1.220 0.440 1.340 1.000 ;
        RECT  1.220 2.440 1.320 2.600 ;
        RECT  1.180 0.440 1.220 2.600 ;
        RECT  1.060 0.840 1.180 2.600 ;
        RECT  0.620 0.990 0.900 2.550 ;
    END
END MXI3XLTR

MACRO MXI3X4TR
    CLASS CORE ;
    FOREIGN MXI3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.810 0.440 7.920 1.440 ;
        RECT  7.570 0.440 7.810 3.160 ;
        RECT  7.470 1.930 7.570 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.640 6.320 1.960 ;
        RECT  5.920 1.640 6.080 1.800 ;
        END
        ANTENNAGATEAREA 0.3528 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.140 3.120 1.560 ;
        END
        ANTENNAGATEAREA 0.2976 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.600 3.640 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.410 2.720 1.960 ;
        RECT  2.280 1.410 2.440 1.690 ;
        END
        ANTENNAGATEAREA 0.1896 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.650 0.680 1.900 ;
        RECT  0.330 1.240 0.340 1.900 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.2088 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.310 -0.280 8.400 0.280 ;
        RECT  8.080 -0.280 8.310 1.310 ;
        RECT  7.310 -0.280 8.080 0.280 ;
        RECT  7.030 -0.280 7.310 0.340 ;
        RECT  6.400 -0.280 7.030 0.280 ;
        RECT  6.120 -0.280 6.400 0.340 ;
        RECT  3.940 -0.280 6.120 0.280 ;
        RECT  3.640 -0.280 3.940 0.640 ;
        RECT  2.760 -0.280 3.640 0.280 ;
        RECT  2.480 -0.280 2.760 0.610 ;
        RECT  0.600 -0.280 2.480 0.280 ;
        RECT  0.270 -0.280 0.600 0.940 ;
        RECT  0.000 -0.280 0.270 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.230 3.320 8.400 3.880 ;
        RECT  7.970 1.910 8.230 3.880 ;
        RECT  7.230 3.320 7.970 3.880 ;
        RECT  6.920 3.070 7.230 3.880 ;
        RECT  6.340 3.320 6.920 3.880 ;
        RECT  6.060 3.260 6.340 3.880 ;
        RECT  3.940 3.320 6.060 3.880 ;
        RECT  3.660 3.260 3.940 3.880 ;
        RECT  2.600 3.320 3.660 3.880 ;
        RECT  2.320 2.930 2.600 3.880 ;
        RECT  0.580 3.320 2.320 3.880 ;
        RECT  0.300 2.540 0.580 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.250 0.500 7.410 1.640 ;
        RECT  4.880 0.500 7.250 0.660 ;
        RECT  6.960 1.900 7.120 2.910 ;
        RECT  6.800 1.470 6.960 2.060 ;
        RECT  5.900 2.750 6.960 2.910 ;
        RECT  6.700 1.030 6.860 1.310 ;
        RECT  6.640 2.220 6.800 2.590 ;
        RECT  6.640 1.150 6.700 1.310 ;
        RECT  6.480 1.150 6.640 2.590 ;
        RECT  5.580 2.430 6.480 2.590 ;
        RECT  5.780 0.820 5.940 1.100 ;
        RECT  5.760 1.960 5.920 2.270 ;
        RECT  5.740 2.750 5.900 3.160 ;
        RECT  5.760 0.940 5.780 1.100 ;
        RECT  5.640 0.940 5.760 2.270 ;
        RECT  4.260 3.000 5.740 3.160 ;
        RECT  5.600 0.940 5.640 2.120 ;
        RECT  5.520 1.410 5.600 1.690 ;
        RECT  5.360 2.430 5.580 2.840 ;
        RECT  5.200 0.820 5.360 2.840 ;
        RECT  4.880 2.050 5.040 2.840 ;
        RECT  4.720 0.500 4.880 2.220 ;
        RECT  4.280 0.440 4.440 2.780 ;
        RECT  4.240 0.440 4.280 1.310 ;
        RECT  4.100 2.940 4.260 3.160 ;
        RECT  3.960 1.430 4.120 1.710 ;
        RECT  2.920 2.940 4.100 3.100 ;
        RECT  3.800 1.150 3.960 2.730 ;
        RECT  3.440 1.150 3.800 1.310 ;
        RECT  3.140 2.570 3.800 2.730 ;
        RECT  3.280 1.030 3.440 1.310 ;
        RECT  3.140 0.550 3.280 0.710 ;
        RECT  2.980 0.550 3.140 0.930 ;
        RECT  2.840 2.100 3.120 2.280 ;
        RECT  1.800 0.770 2.980 0.930 ;
        RECT  2.760 2.610 2.920 3.100 ;
        RECT  2.440 2.120 2.840 2.280 ;
        RECT  1.500 2.610 2.760 2.770 ;
        RECT  2.280 2.120 2.440 2.450 ;
        RECT  1.640 2.290 2.280 2.450 ;
        RECT  2.120 1.090 2.240 1.250 ;
        RECT  1.960 1.090 2.120 2.130 ;
        RECT  1.800 1.970 1.960 2.130 ;
        RECT  1.640 0.770 1.800 1.770 ;
        RECT  1.480 1.610 1.640 2.450 ;
        RECT  1.340 2.610 1.500 2.890 ;
        RECT  1.320 0.880 1.480 1.160 ;
        RECT  1.320 2.610 1.340 2.770 ;
        RECT  1.160 1.000 1.320 2.770 ;
        RECT  0.840 0.590 1.000 3.160 ;
    END
END MXI3X4TR

MACRO MXI3X2TR
    CLASS CORE ;
    FOREIGN MXI3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.360 0.440 7.520 3.160 ;
        RECT  7.230 0.440 7.360 1.310 ;
        RECT  7.230 1.970 7.360 3.160 ;
        END
        ANTENNADIFFAREA 3.456 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.640 6.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.840 1.240 3.160 ;
        END
        ANTENNAGATEAREA 0.2304 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.340 1.630 3.520 2.020 ;
        RECT  3.190 1.640 3.340 2.020 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.210 2.360 1.600 ;
        RECT  2.030 1.320 2.040 1.600 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.030 -0.280 7.600 0.280 ;
        RECT  6.750 -0.280 7.030 0.670 ;
        RECT  6.470 -0.280 6.750 0.280 ;
        RECT  6.190 -0.280 6.470 0.670 ;
        RECT  3.690 -0.280 6.190 0.280 ;
        RECT  3.510 -0.280 3.690 1.040 ;
        RECT  3.410 -0.280 3.510 0.400 ;
        RECT  2.470 -0.280 3.410 0.280 ;
        RECT  2.190 -0.280 2.470 0.990 ;
        RECT  0.370 -0.280 2.190 0.340 ;
        RECT  0.090 -0.280 0.370 1.030 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.030 3.320 7.600 3.880 ;
        RECT  6.750 2.580 7.030 3.880 ;
        RECT  6.150 3.320 6.750 3.880 ;
        RECT  5.930 2.610 6.150 3.880 ;
        RECT  3.890 3.260 5.930 3.880 ;
        RECT  3.610 3.200 3.890 3.880 ;
        RECT  2.510 3.260 3.610 3.880 ;
        RECT  2.230 2.860 2.510 3.880 ;
        RECT  0.370 3.320 2.230 3.880 ;
        RECT  0.090 2.550 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.070 1.470 7.200 1.750 ;
        RECT  6.910 0.830 7.070 1.750 ;
        RECT  6.030 0.830 6.910 0.990 ;
        RECT  6.090 1.150 6.670 1.370 ;
        RECT  6.090 2.120 6.670 2.400 ;
        RECT  5.930 1.150 6.090 2.400 ;
        RECT  5.870 0.450 6.030 0.990 ;
        RECT  5.710 1.150 5.930 1.370 ;
        RECT  4.610 0.450 5.870 0.610 ;
        RECT  5.550 1.640 5.770 2.780 ;
        RECT  5.550 0.770 5.710 1.370 ;
        RECT  5.010 0.770 5.550 0.930 ;
        RECT  2.830 2.620 5.550 2.780 ;
        RECT  5.170 1.090 5.390 2.370 ;
        RECT  4.850 0.770 5.010 1.700 ;
        RECT  4.850 2.090 4.970 2.370 ;
        RECT  4.770 1.420 4.850 1.700 ;
        RECT  4.690 1.860 4.850 2.370 ;
        RECT  4.610 0.770 4.690 1.050 ;
        RECT  4.610 1.860 4.690 2.020 ;
        RECT  4.450 0.450 4.610 2.020 ;
        RECT  4.290 2.180 4.410 2.460 ;
        RECT  4.130 0.880 4.290 2.460 ;
        RECT  3.930 0.880 4.130 1.160 ;
        RECT  3.840 1.420 3.970 1.700 ;
        RECT  3.680 1.310 3.840 2.340 ;
        RECT  3.350 1.310 3.680 1.470 ;
        RECT  3.450 2.180 3.680 2.340 ;
        RECT  3.170 2.180 3.450 2.460 ;
        RECT  3.190 0.570 3.350 1.470 ;
        RECT  2.890 0.570 3.190 0.850 ;
        RECT  2.990 1.030 3.030 1.310 ;
        RECT  2.750 1.030 2.990 2.380 ;
        RECT  2.670 2.540 2.830 2.780 ;
        RECT  2.710 1.760 2.750 2.380 ;
        RECT  1.870 1.760 2.710 1.920 ;
        RECT  1.510 2.540 2.670 2.700 ;
        RECT  1.710 2.080 1.990 2.380 ;
        RECT  1.760 0.840 1.880 1.120 ;
        RECT  1.650 1.510 1.870 1.920 ;
        RECT  1.600 0.840 1.760 1.350 ;
        RECT  1.490 2.080 1.710 2.240 ;
        RECT  1.490 1.190 1.600 1.350 ;
        RECT  1.350 2.400 1.510 2.700 ;
        RECT  1.330 1.190 1.490 2.240 ;
        RECT  1.170 0.810 1.400 1.030 ;
        RECT  1.170 2.400 1.350 2.680 ;
        RECT  1.010 0.810 1.170 2.680 ;
        RECT  0.570 0.920 0.850 2.680 ;
    END
END MXI3X2TR

MACRO MXI3X1TR
    CLASS CORE ;
    FOREIGN MXI3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 0.440 7.120 3.000 ;
        RECT  6.860 0.440 6.960 0.720 ;
        RECT  6.880 1.640 6.960 3.000 ;
        RECT  6.800 2.580 6.880 3.000 ;
        END
        ANTENNADIFFAREA 1.664 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.640 6.480 1.960 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 2.840 1.120 3.160 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.640 3.520 2.080 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.240 2.360 1.660 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.200 0.400 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.560 -0.280 7.200 0.280 ;
        RECT  6.280 -0.280 6.560 0.400 ;
        RECT  5.660 -0.280 6.280 0.280 ;
        RECT  5.500 -0.280 5.660 0.840 ;
        RECT  3.560 -0.280 5.500 0.340 ;
        RECT  3.280 -0.280 3.560 0.400 ;
        RECT  2.440 -0.280 3.280 0.340 ;
        RECT  2.160 -0.280 2.440 1.080 ;
        RECT  0.370 -0.280 2.160 0.280 ;
        RECT  0.090 -0.280 0.370 0.350 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.600 3.320 7.200 3.880 ;
        RECT  6.320 2.830 6.600 3.880 ;
        RECT  5.980 3.320 6.320 3.880 ;
        RECT  5.760 2.610 5.980 3.880 ;
        RECT  3.900 3.260 5.760 3.880 ;
        RECT  3.620 3.200 3.900 3.880 ;
        RECT  2.440 3.260 3.620 3.880 ;
        RECT  2.160 3.000 2.440 3.880 ;
        RECT  0.370 3.320 2.160 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.680 1.100 6.800 1.380 ;
        RECT  6.520 0.670 6.680 1.380 ;
        RECT  5.920 2.120 6.540 2.400 ;
        RECT  5.980 0.670 6.520 0.830 ;
        RECT  6.140 0.990 6.360 1.480 ;
        RECT  5.920 1.320 6.140 1.480 ;
        RECT  5.820 0.670 5.980 1.160 ;
        RECT  5.760 1.320 5.920 2.400 ;
        RECT  5.340 1.000 5.820 1.160 ;
        RECT  5.380 1.320 5.760 1.480 ;
        RECT  5.440 2.010 5.600 3.020 ;
        RECT  5.380 2.010 5.440 2.290 ;
        RECT  2.760 2.860 5.440 3.020 ;
        RECT  5.100 1.320 5.380 1.850 ;
        RECT  5.180 0.560 5.340 1.160 ;
        RECT  5.060 2.010 5.220 2.700 ;
        RECT  4.620 0.560 5.180 0.720 ;
        RECT  4.940 2.010 5.060 2.170 ;
        RECT  4.940 0.880 5.020 1.160 ;
        RECT  4.780 0.880 4.940 2.170 ;
        RECT  4.620 2.330 4.800 2.610 ;
        RECT  4.460 0.560 4.620 2.610 ;
        RECT  4.320 0.820 4.460 1.100 ;
        RECT  4.160 1.260 4.300 2.520 ;
        RECT  4.060 0.940 4.160 2.520 ;
        RECT  4.020 0.820 4.060 2.520 ;
        RECT  4.000 0.820 4.020 1.360 ;
        RECT  3.780 0.820 4.000 1.100 ;
        RECT  3.680 1.260 3.840 2.400 ;
        RECT  3.320 1.260 3.680 1.480 ;
        RECT  3.340 2.240 3.680 2.400 ;
        RECT  3.060 2.240 3.340 2.520 ;
        RECT  3.160 0.690 3.320 1.480 ;
        RECT  3.000 0.690 3.160 0.850 ;
        RECT  2.720 0.570 3.000 0.850 ;
        RECT  2.880 1.030 3.000 1.980 ;
        RECT  2.720 1.030 2.880 2.520 ;
        RECT  2.600 2.680 2.760 3.020 ;
        RECT  2.600 1.820 2.720 2.520 ;
        RECT  1.880 1.820 2.600 1.980 ;
        RECT  1.520 2.680 2.600 2.840 ;
        RECT  1.600 1.680 1.880 1.980 ;
        RECT  1.760 2.300 1.880 2.520 ;
        RECT  1.590 1.030 1.870 1.310 ;
        RECT  1.600 2.140 1.760 2.520 ;
        RECT  1.440 2.140 1.600 2.300 ;
        RECT  1.440 1.150 1.590 1.310 ;
        RECT  1.440 2.680 1.520 3.160 ;
        RECT  1.280 1.150 1.440 2.300 ;
        RECT  1.280 2.460 1.440 3.160 ;
        RECT  1.120 0.440 1.310 0.730 ;
        RECT  1.120 2.460 1.280 2.620 ;
        RECT  0.960 0.440 1.120 2.620 ;
        RECT  0.640 1.030 0.800 2.550 ;
    END
END MXI3X1TR

MACRO MXI2XLTR
    CLASS CORE ;
    FOREIGN MXI2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.520 2.110 3.160 ;
        RECT  1.650 0.520 1.950 0.780 ;
        RECT  1.500 2.840 1.950 3.160 ;
        END
        ANTENNADIFFAREA 2.048 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.840 2.720 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.850 1.060 2.130 ;
        RECT  0.480 1.850 0.760 2.360 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.120 2.360 ;
        RECT  2.840 1.240 2.880 1.730 ;
        RECT  2.650 1.450 2.840 1.730 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.280 3.200 0.280 ;
        RECT  2.820 -0.280 3.110 0.740 ;
        RECT  0.930 -0.280 2.820 0.280 ;
        RECT  0.650 -0.280 0.930 1.290 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 3.320 3.200 3.880 ;
        RECT  2.880 2.770 3.110 3.880 ;
        RECT  0.940 3.320 2.880 3.880 ;
        RECT  0.660 2.960 0.940 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 1.010 2.550 1.290 ;
        RECT  2.270 1.010 2.490 2.550 ;
        RECT  1.630 0.960 1.790 2.530 ;
        RECT  1.370 0.960 1.630 1.120 ;
        RECT  1.340 2.370 1.630 2.530 ;
        RECT  1.250 1.530 1.470 1.960 ;
        RECT  1.210 0.460 1.370 1.120 ;
        RECT  1.060 2.370 1.340 2.650 ;
        RECT  0.370 1.530 1.250 1.690 ;
        RECT  1.090 0.460 1.210 0.740 ;
        RECT  0.320 1.010 0.370 1.690 ;
        RECT  0.160 1.010 0.320 2.550 ;
        RECT  0.090 1.010 0.160 1.290 ;
        RECT  0.090 2.270 0.160 2.550 ;
    END
END MXI2XLTR

MACRO MXI2X8TR
    CLASS CORE ;
    FOREIGN MXI2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.080 0.460 15.800 2.990 ;
        RECT  2.390 0.460 15.080 0.940 ;
        RECT  2.330 2.510 15.080 2.990 ;
        END
        ANTENNADIFFAREA 21.312 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.080 1.450 14.390 1.610 ;
        RECT  8.920 1.450 9.080 2.030 ;
        RECT  7.450 1.870 8.920 2.030 ;
        RECT  7.170 1.810 7.450 2.030 ;
        RECT  5.770 1.870 7.170 2.030 ;
        RECT  5.490 1.810 5.770 2.030 ;
        RECT  4.090 1.870 5.490 2.030 ;
        RECT  3.810 1.810 4.090 2.030 ;
        RECT  2.470 1.870 3.810 2.030 ;
        RECT  2.250 1.810 2.470 2.030 ;
        RECT  0.760 1.870 2.250 2.030 ;
        RECT  0.480 1.600 0.760 2.030 ;
        END
        ANTENNAGATEAREA 1.8456 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.760 1.100 14.920 1.700 ;
        RECT  8.720 1.100 14.760 1.290 ;
        RECT  8.480 1.100 8.720 1.570 ;
        END
        ANTENNAGATEAREA 1.4208 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.130 8.310 1.290 ;
        RECT  1.770 0.840 1.920 1.290 ;
        RECT  1.510 0.840 1.770 1.370 ;
        END
        ANTENNAGATEAREA 1.4208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.430 -0.280 16.000 0.280 ;
        RECT  15.150 -0.280 15.430 0.300 ;
        RECT  13.750 -0.280 15.150 0.280 ;
        RECT  13.470 -0.280 13.750 0.300 ;
        RECT  11.950 -0.280 13.470 0.280 ;
        RECT  11.670 -0.280 11.950 0.300 ;
        RECT  10.230 -0.280 11.670 0.280 ;
        RECT  9.950 -0.280 10.230 0.300 ;
        RECT  8.550 -0.280 9.950 0.280 ;
        RECT  8.270 -0.280 8.550 0.300 ;
        RECT  6.870 -0.280 8.270 0.280 ;
        RECT  6.590 -0.280 6.870 0.300 ;
        RECT  5.190 -0.280 6.590 0.280 ;
        RECT  4.910 -0.280 5.190 0.300 ;
        RECT  3.510 -0.280 4.910 0.280 ;
        RECT  3.230 -0.280 3.510 0.300 ;
        RECT  1.810 -0.280 3.230 0.280 ;
        RECT  1.530 -0.280 1.810 0.680 ;
        RECT  0.850 -0.280 1.530 0.280 ;
        RECT  0.570 -0.280 0.850 0.720 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.310 3.320 16.000 3.880 ;
        RECT  15.030 3.200 15.310 3.880 ;
        RECT  13.630 3.320 15.030 3.880 ;
        RECT  13.350 3.200 13.630 3.880 ;
        RECT  11.950 3.320 13.350 3.880 ;
        RECT  11.670 3.200 11.950 3.880 ;
        RECT  10.270 3.320 11.670 3.880 ;
        RECT  9.990 3.200 10.270 3.880 ;
        RECT  8.550 3.320 9.990 3.880 ;
        RECT  8.270 3.200 8.550 3.880 ;
        RECT  6.810 3.320 8.270 3.880 ;
        RECT  6.530 3.200 6.810 3.880 ;
        RECT  5.130 3.320 6.530 3.880 ;
        RECT  4.850 3.200 5.130 3.880 ;
        RECT  3.450 3.320 4.850 3.880 ;
        RECT  3.170 3.200 3.450 3.880 ;
        RECT  1.810 3.320 3.170 3.880 ;
        RECT  1.530 2.510 1.810 3.880 ;
        RECT  0.850 3.320 1.530 3.880 ;
        RECT  0.570 2.510 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  14.190 1.800 14.310 2.080 ;
        RECT  14.030 1.800 14.190 2.350 ;
        RECT  12.710 2.190 14.030 2.350 ;
        RECT  12.430 1.800 12.710 2.350 ;
        RECT  11.320 2.190 12.430 2.350 ;
        RECT  11.030 1.800 11.320 2.350 ;
        RECT  9.600 2.190 11.030 2.350 ;
        RECT  9.380 1.800 9.600 2.350 ;
        RECT  1.330 2.190 9.380 2.350 ;
        RECT  2.090 1.460 7.870 1.630 ;
        RECT  1.930 1.460 2.090 1.710 ;
        RECT  1.330 1.550 1.930 1.710 ;
        RECT  1.170 0.440 1.330 1.710 ;
        RECT  1.050 2.190 1.330 2.790 ;
        RECT  1.050 0.440 1.170 1.240 ;
        RECT  0.370 1.080 1.050 1.240 ;
        RECT  0.370 2.190 1.050 2.350 ;
        RECT  0.310 0.440 0.370 1.240 ;
        RECT  0.310 2.190 0.370 2.790 ;
        RECT  0.150 0.440 0.310 2.790 ;
        RECT  0.090 0.440 0.150 1.240 ;
        RECT  0.090 1.930 0.150 2.790 ;
    END
END MXI2X8TR

MACRO MXI2X6TR
    CLASS CORE ;
    FOREIGN MXI2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.710 0.480 11.720 2.560 ;
        RECT  11.360 0.480 11.710 2.720 ;
        RECT  6.920 0.480 11.360 0.780 ;
        RECT  11.080 1.840 11.360 2.720 ;
        RECT  0.920 2.340 11.080 2.720 ;
        RECT  0.960 0.480 6.920 0.640 ;
        END
        ANTENNADIFFAREA 11.88 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.200 1.260 10.720 1.420 ;
        RECT  10.040 1.260 10.200 1.560 ;
        RECT  9.440 1.400 10.040 1.560 ;
        RECT  9.280 1.260 9.440 1.560 ;
        RECT  8.600 1.260 9.280 1.420 ;
        RECT  8.440 1.260 8.600 1.550 ;
        RECT  7.900 1.390 8.440 1.550 ;
        RECT  7.740 1.260 7.900 1.550 ;
        RECT  7.080 1.260 7.740 1.420 ;
        RECT  6.920 1.260 7.080 1.560 ;
        RECT  5.960 1.400 6.920 1.560 ;
        RECT  5.840 1.240 5.960 1.560 ;
        RECT  5.680 1.240 5.840 1.840 ;
        RECT  4.360 1.680 5.680 1.840 ;
        RECT  4.080 1.560 4.360 1.840 ;
        RECT  2.680 1.680 4.080 1.840 ;
        RECT  2.400 1.560 2.680 1.840 ;
        RECT  1.040 1.680 2.400 1.840 ;
        RECT  0.820 1.560 1.040 1.840 ;
        END
        ANTENNAGATEAREA 1.1088 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.020 0.940 11.180 1.660 ;
        RECT  9.820 0.940 11.020 1.100 ;
        RECT  9.600 0.940 9.820 1.240 ;
        RECT  8.220 0.940 9.600 1.100 ;
        RECT  8.060 0.940 8.220 1.230 ;
        RECT  6.760 0.940 8.060 1.100 ;
        RECT  6.720 0.940 6.760 1.160 ;
        RECT  6.440 0.840 6.720 1.160 ;
        END
        ANTENNAGATEAREA 0.792 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.080 0.920 5.200 1.200 ;
        RECT  4.920 0.830 5.080 1.200 ;
        RECT  3.560 0.830 4.920 0.990 ;
        RECT  3.280 0.830 3.560 1.200 ;
        RECT  1.880 0.830 3.280 0.990 ;
        RECT  1.600 0.830 1.880 1.200 ;
        RECT  0.320 0.830 1.600 0.990 ;
        RECT  0.180 0.830 0.320 1.960 ;
        RECT  0.080 0.840 0.180 1.960 ;
        END
        ANTENNAGATEAREA 0.792 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.760 -0.280 12.000 0.280 ;
        RECT  11.480 -0.280 11.760 0.320 ;
        RECT  10.080 -0.280 11.480 0.280 ;
        RECT  9.800 -0.280 10.080 0.320 ;
        RECT  8.330 -0.280 9.800 0.280 ;
        RECT  8.050 -0.280 8.330 0.320 ;
        RECT  6.520 -0.280 8.050 0.280 ;
        RECT  6.240 -0.280 6.520 0.320 ;
        RECT  5.970 -0.280 6.240 0.280 ;
        RECT  5.160 -0.280 5.970 0.320 ;
        RECT  3.760 -0.280 5.160 0.280 ;
        RECT  3.480 -0.280 3.760 0.320 ;
        RECT  2.080 -0.280 3.480 0.280 ;
        RECT  1.800 -0.280 2.080 0.320 ;
        RECT  0.400 -0.280 1.800 0.280 ;
        RECT  0.120 -0.280 0.400 0.670 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.540 3.320 12.000 3.880 ;
        RECT  11.240 2.940 11.540 3.880 ;
        RECT  9.840 3.320 11.240 3.880 ;
        RECT  9.560 3.010 9.840 3.880 ;
        RECT  8.240 3.320 9.560 3.880 ;
        RECT  7.960 3.010 8.240 3.880 ;
        RECT  6.480 3.320 7.960 3.880 ;
        RECT  6.200 2.940 6.480 3.880 ;
        RECT  5.440 3.280 6.200 3.880 ;
        RECT  5.160 2.940 5.440 3.880 ;
        RECT  3.720 3.280 5.160 3.880 ;
        RECT  3.440 2.880 3.720 3.880 ;
        RECT  2.040 3.280 3.440 3.880 ;
        RECT  1.760 2.880 2.040 3.880 ;
        RECT  0.400 3.280 1.760 3.880 ;
        RECT  0.120 2.370 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.360 1.600 10.640 1.880 ;
        RECT  9.040 1.720 10.360 1.880 ;
        RECT  8.760 1.600 9.040 1.880 ;
        RECT  7.560 1.720 8.760 1.880 ;
        RECT  7.270 1.660 7.560 1.880 ;
        RECT  6.160 1.720 7.270 1.880 ;
        RECT  6.000 1.720 6.160 2.160 ;
        RECT  5.520 0.800 6.000 1.080 ;
        RECT  0.660 2.000 6.000 2.160 ;
        RECT  5.360 0.800 5.520 1.520 ;
        RECT  4.760 1.360 5.360 1.520 ;
        RECT  4.600 1.150 4.760 1.520 ;
        RECT  4.480 1.150 4.600 1.430 ;
        RECT  3.880 1.150 4.480 1.310 ;
        RECT  3.720 1.150 3.880 1.520 ;
        RECT  3.120 1.360 3.720 1.520 ;
        RECT  2.960 1.150 3.120 1.520 ;
        RECT  2.840 1.150 2.960 1.430 ;
        RECT  2.200 1.150 2.840 1.310 ;
        RECT  2.040 1.150 2.200 1.520 ;
        RECT  1.440 1.360 2.040 1.520 ;
        RECT  1.280 1.150 1.440 1.520 ;
        RECT  1.160 1.150 1.280 1.430 ;
        RECT  0.660 1.150 1.160 1.310 ;
        RECT  0.500 1.150 0.660 2.160 ;
    END
END MXI2X6TR

MACRO MXI2X4TR
    CLASS CORE ;
    FOREIGN MXI2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.870 0.940 4.950 1.920 ;
        RECT  4.710 0.940 4.870 2.270 ;
        RECT  3.920 0.940 4.710 1.180 ;
        RECT  4.590 1.840 4.710 2.270 ;
        RECT  3.950 1.840 4.590 2.080 ;
        RECT  3.680 1.840 3.950 2.720 ;
        RECT  3.670 0.480 3.920 1.180 ;
        RECT  2.670 2.440 3.680 2.720 ;
        RECT  2.810 0.480 3.670 0.720 ;
        END
        ANTENNADIFFAREA 8.962 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.840 2.840 5.120 3.160 ;
        RECT  4.800 2.880 4.840 3.160 ;
        RECT  0.760 2.880 4.800 3.040 ;
        RECT  0.510 2.690 0.760 3.040 ;
        END
        ANTENNAGATEAREA 0.7224 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.360 2.230 1.640 ;
        RECT  1.240 1.240 1.560 1.640 ;
        RECT  1.210 1.360 1.240 1.640 ;
        END
        ANTENNAGATEAREA 0.528 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.560 1.600 5.970 1.880 ;
        RECT  5.240 1.600 5.560 1.960 ;
        END
        ANTENNAGATEAREA 0.528 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 -0.280 6.400 0.280 ;
        RECT  5.530 -0.280 5.810 1.070 ;
        RECT  2.090 -0.280 5.530 0.280 ;
        RECT  0.090 -0.280 2.090 0.340 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 3.320 6.400 3.880 ;
        RECT  5.530 2.440 5.810 3.880 ;
        RECT  2.210 3.320 5.530 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  1.170 3.320 1.930 3.880 ;
        RECT  0.890 3.200 1.170 3.880 ;
        RECT  0.370 3.260 0.890 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.130 0.440 6.290 3.160 ;
        RECT  6.010 0.440 6.130 1.390 ;
        RECT  6.010 2.120 6.130 3.160 ;
        RECT  5.330 1.230 6.010 1.390 ;
        RECT  5.330 2.120 6.010 2.280 ;
        RECT  5.110 0.440 5.330 1.390 ;
        RECT  5.050 2.120 5.330 2.680 ;
        RECT  4.370 0.440 5.110 0.600 ;
        RECT  4.390 2.460 5.050 2.680 ;
        RECT  3.380 1.410 4.510 1.570 ;
        RECT  4.110 2.390 4.390 2.680 ;
        RECT  4.100 0.440 4.370 0.720 ;
        RECT  3.290 0.880 3.510 1.160 ;
        RECT  1.690 2.120 3.430 2.280 ;
        RECT  3.210 1.410 3.380 1.960 ;
        RECT  2.610 1.000 3.290 1.160 ;
        RECT  0.770 1.800 3.210 1.960 ;
        RECT  2.330 0.550 2.610 1.160 ;
        RECT  1.690 0.920 2.330 1.080 ;
        RECT  1.570 0.800 1.690 1.080 ;
        RECT  1.410 2.120 1.690 2.530 ;
        RECT  1.410 0.710 1.570 1.080 ;
        RECT  0.330 0.710 1.410 0.870 ;
        RECT  0.330 2.370 1.410 2.530 ;
        RECT  0.610 1.030 0.770 2.210 ;
        RECT  0.490 1.030 0.610 1.310 ;
        RECT  0.490 1.930 0.610 2.210 ;
        RECT  0.170 0.710 0.330 2.530 ;
    END
END MXI2X4TR

MACRO MXI2X2TR
    CLASS CORE ;
    FOREIGN MXI2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.610 2.960 2.760 ;
        RECT  2.380 0.610 2.800 0.770 ;
        RECT  2.480 2.440 2.800 2.760 ;
        RECT  1.900 2.560 2.480 2.720 ;
        RECT  2.100 0.490 2.380 0.770 ;
        RECT  1.740 2.270 1.900 2.720 ;
        RECT  1.620 2.270 1.740 2.490 ;
        END
        ANTENNADIFFAREA 4.752 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 2.880 2.170 3.100 ;
        RECT  0.750 2.880 1.950 3.040 ;
        RECT  0.470 2.440 0.750 3.040 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.570 1.370 1.790 ;
        RECT  0.880 1.570 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.2256 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.320 3.920 2.280 ;
        RECT  3.670 1.640 3.680 2.280 ;
        RECT  3.440 1.640 3.670 1.960 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.280 4.000 0.280 ;
        RECT  3.540 -0.280 3.820 1.060 ;
        RECT  1.230 -0.280 3.540 0.280 ;
        RECT  0.900 -0.280 1.230 1.060 ;
        RECT  0.000 -0.280 0.900 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 3.320 4.000 3.880 ;
        RECT  3.540 2.590 3.820 3.880 ;
        RECT  0.920 3.320 3.540 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.120 0.440 3.280 3.160 ;
        RECT  2.480 0.930 2.640 2.110 ;
        RECT  1.780 0.930 2.480 1.090 ;
        RECT  2.320 1.950 2.480 2.110 ;
        RECT  2.100 1.250 2.320 1.790 ;
        RECT  2.100 1.950 2.320 2.390 ;
        RECT  0.640 1.250 2.100 1.410 ;
        RECT  1.440 1.950 2.100 2.110 ;
        RECT  1.500 0.810 1.780 1.090 ;
        RECT  1.280 1.950 1.440 2.550 ;
        RECT  1.160 2.230 1.280 2.550 ;
        RECT  0.440 0.730 0.640 1.410 ;
        RECT  0.360 0.730 0.440 2.270 ;
        RECT  0.280 1.210 0.360 2.270 ;
        RECT  0.160 2.050 0.280 2.270 ;
    END
END MXI2X2TR

MACRO MXI2X1TR
    CLASS CORE ;
    FOREIGN MXI2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.780 2.150 2.760 ;
        RECT  1.760 0.780 1.990 1.060 ;
        RECT  1.680 2.440 1.990 2.760 ;
        END
        ANTENNADIFFAREA 2.046 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.940 2.290 3.100 ;
        RECT  1.280 2.770 1.520 3.160 ;
        RECT  0.570 2.770 1.280 2.930 ;
        RECT  0.260 2.650 0.570 2.930 ;
        END
        ANTENNAGATEAREA 0.1896 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.860 1.100 2.140 ;
        RECT  0.480 1.860 0.760 2.360 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.190 3.120 2.360 ;
        RECT  2.630 1.190 2.860 1.630 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.010 -0.280 3.200 0.280 ;
        RECT  2.730 -0.280 3.010 1.030 ;
        RECT  1.020 -0.280 2.730 0.340 ;
        RECT  0.720 -0.280 1.020 1.030 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 3.320 3.200 3.880 ;
        RECT  2.720 2.550 3.000 3.880 ;
        RECT  0.970 3.320 2.720 3.880 ;
        RECT  0.660 3.200 0.970 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.310 0.930 2.470 2.780 ;
        RECT  1.670 1.220 1.830 2.200 ;
        RECT  1.560 1.220 1.670 1.380 ;
        RECT  1.490 2.040 1.670 2.200 ;
        RECT  1.280 0.930 1.560 1.380 ;
        RECT  1.270 1.540 1.510 1.880 ;
        RECT  1.300 2.040 1.490 2.490 ;
        RECT  0.370 1.540 1.270 1.700 ;
        RECT  0.320 0.930 0.370 1.700 ;
        RECT  0.160 0.930 0.320 2.490 ;
        RECT  0.090 0.930 0.160 1.210 ;
        RECT  0.090 2.210 0.160 2.490 ;
    END
END MXI2X1TR

MACRO MX4XLTR
    CLASS CORE ;
    FOREIGN MX4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.260 2.010 8.300 2.360 ;
        RECT  8.090 0.440 8.260 2.360 ;
        RECT  7.680 2.010 8.090 2.360 ;
        END
        ANTENNADIFFAREA 1.202 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.600 0.440 5.920 0.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.510 2.800 1.670 ;
        RECT  2.520 0.840 2.720 1.670 ;
        RECT  2.480 0.840 2.520 1.160 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.230 2.320 1.580 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.200 0.490 1.580 ;
        RECT  0.080 1.200 0.340 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.840 3.520 1.270 ;
        END
        ANTENNAGATEAREA 0.0552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.220 5.220 1.580 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.750 -0.280 8.400 0.280 ;
        RECT  7.470 -0.280 7.750 0.340 ;
        RECT  5.440 -0.280 7.470 0.280 ;
        RECT  5.220 -0.280 5.440 0.980 ;
        RECT  3.100 -0.280 5.220 0.280 ;
        RECT  2.880 -0.280 3.100 0.890 ;
        RECT  2.490 -0.280 2.880 0.280 ;
        RECT  2.220 -0.280 2.490 0.680 ;
        RECT  0.310 -0.280 2.220 0.280 ;
        RECT  0.150 -0.280 0.310 0.740 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.780 3.320 8.400 3.880 ;
        RECT  7.560 2.520 7.780 3.880 ;
        RECT  5.260 3.320 7.560 3.880 ;
        RECT  4.980 3.000 5.260 3.880 ;
        RECT  3.100 3.320 4.980 3.880 ;
        RECT  2.820 2.720 3.100 3.880 ;
        RECT  2.490 3.320 2.820 3.880 ;
        RECT  2.210 2.720 2.490 3.880 ;
        RECT  0.370 3.320 2.210 3.880 ;
        RECT  0.090 2.800 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.750 0.500 7.910 1.100 ;
        RECT  6.930 0.500 7.750 0.660 ;
        RECT  7.400 0.890 7.570 1.050 ;
        RECT  7.240 0.890 7.400 2.840 ;
        RECT  3.580 2.680 7.240 2.840 ;
        RECT  6.850 0.500 6.930 1.060 ;
        RECT  6.670 0.500 6.850 2.390 ;
        RECT  6.360 0.640 6.480 2.520 ;
        RECT  6.320 0.470 6.360 2.520 ;
        RECT  6.200 0.470 6.320 0.800 ;
        RECT  4.320 2.360 6.320 2.520 ;
        RECT  6.060 1.300 6.140 1.680 ;
        RECT  5.980 0.990 6.060 1.680 ;
        RECT  5.790 0.990 5.980 2.200 ;
        RECT  5.420 2.040 5.790 2.200 ;
        RECT  4.680 0.760 4.940 0.920 ;
        RECT  4.680 2.040 4.840 2.200 ;
        RECT  4.520 0.760 4.680 2.200 ;
        RECT  4.160 0.690 4.320 2.520 ;
        RECT  3.940 2.360 4.160 2.520 ;
        RECT  3.840 0.510 4.000 2.200 ;
        RECT  3.300 0.510 3.840 0.670 ;
        RECT  3.380 2.040 3.840 2.200 ;
        RECT  3.520 1.520 3.680 1.790 ;
        RECT  3.420 2.400 3.580 2.840 ;
        RECT  3.120 1.580 3.520 1.790 ;
        RECT  1.480 2.400 3.420 2.560 ;
        RECT  3.040 1.190 3.120 2.190 ;
        RECT  2.960 1.070 3.040 2.190 ;
        RECT  2.880 1.070 2.960 1.350 ;
        RECT  2.370 2.030 2.960 2.190 ;
        RECT  2.210 1.760 2.370 2.190 ;
        RECT  1.770 1.760 2.210 1.920 ;
        RECT  1.450 2.080 2.050 2.240 ;
        RECT  1.760 0.910 2.040 1.070 ;
        RECT  1.610 1.640 1.770 1.920 ;
        RECT  1.600 0.910 1.760 1.440 ;
        RECT  1.450 1.280 1.600 1.440 ;
        RECT  1.230 2.400 1.480 2.840 ;
        RECT  1.290 1.280 1.450 2.240 ;
        RECT  1.130 0.830 1.440 1.120 ;
        RECT  1.130 2.400 1.230 2.560 ;
        RECT  0.970 0.830 1.130 2.560 ;
        RECT  0.650 0.970 0.810 2.490 ;
    END
END MX4XLTR

MACRO MX4X4TR
    CLASS CORE ;
    FOREIGN MX4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.430 0.640 9.520 1.360 ;
        RECT  9.150 0.440 9.430 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.360 1.380 8.470 3.000 ;
        RECT  8.310 1.380 8.360 3.160 ;
        RECT  8.190 1.380 8.310 1.660 ;
        RECT  8.040 2.840 8.310 3.160 ;
        RECT  6.700 2.840 8.040 3.120 ;
        END
        ANTENNAGATEAREA 0.3624 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 2.880 5.130 3.160 ;
        RECT  4.210 0.440 4.490 0.720 ;
        RECT  3.590 0.560 4.210 0.720 ;
        RECT  4.040 2.840 4.200 3.160 ;
        RECT  1.560 2.840 4.040 3.000 ;
        RECT  3.310 0.560 3.590 0.870 ;
        RECT  2.180 0.560 3.310 0.720 ;
        RECT  1.900 0.440 2.180 0.720 ;
        RECT  1.110 0.560 1.900 0.720 ;
        RECT  1.280 2.840 1.560 3.160 ;
        RECT  1.110 3.000 1.280 3.160 ;
        RECT  0.950 0.560 1.110 3.160 ;
        END
        ANTENNAGATEAREA 0.72 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.760 2.760 2.360 ;
        RECT  2.440 1.640 2.630 2.360 ;
        RECT  2.350 1.640 2.440 1.920 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.360 0.410 1.640 ;
        RECT  0.320 0.920 0.360 1.640 ;
        RECT  0.080 0.920 0.320 1.880 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.320 4.080 1.600 ;
        RECT  3.640 1.240 3.960 1.600 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.640 6.360 1.960 ;
        RECT  5.760 1.520 6.040 1.800 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.910 -0.280 10.000 0.280 ;
        RECT  9.680 -0.280 9.910 1.310 ;
        RECT  8.950 -0.280 9.680 0.280 ;
        RECT  8.730 -0.280 8.950 0.800 ;
        RECT  6.000 -0.280 8.730 0.340 ;
        RECT  3.690 -0.280 6.000 0.280 ;
        RECT  3.410 -0.280 3.690 0.400 ;
        RECT  0.370 -0.280 3.410 0.280 ;
        RECT  0.090 -0.280 0.370 0.680 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.910 3.320 10.000 3.880 ;
        RECT  9.630 1.910 9.910 3.880 ;
        RECT  8.910 3.320 9.630 3.880 ;
        RECT  8.630 1.910 8.910 3.880 ;
        RECT  6.340 3.320 8.630 3.880 ;
        RECT  6.060 3.200 6.340 3.880 ;
        RECT  3.880 3.320 6.060 3.880 ;
        RECT  3.600 3.200 3.880 3.880 ;
        RECT  2.830 3.260 3.600 3.880 ;
        RECT  2.550 3.180 2.830 3.880 ;
        RECT  0.370 3.320 2.550 3.880 ;
        RECT  0.090 2.110 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.710 0.960 8.990 1.640 ;
        RECT  8.570 0.960 8.710 1.120 ;
        RECT  8.410 0.620 8.570 1.120 ;
        RECT  7.710 0.620 8.410 0.780 ;
        RECT  8.030 0.940 8.250 1.220 ;
        RECT  8.030 1.970 8.150 2.680 ;
        RECT  7.870 1.060 8.030 2.680 ;
        RECT  1.550 2.520 7.870 2.680 ;
        RECT  7.430 0.500 7.710 2.250 ;
        RECT  7.390 1.970 7.430 2.250 ;
        RECT  7.190 0.500 7.230 1.310 ;
        RECT  7.030 0.500 7.190 2.250 ;
        RECT  7.010 0.500 7.030 1.310 ;
        RECT  6.910 1.970 7.030 2.250 ;
        RECT  5.280 0.500 7.010 0.660 ;
        RECT  6.700 1.380 6.850 1.660 ;
        RECT  6.540 0.980 6.700 2.360 ;
        RECT  6.420 0.980 6.540 1.260 ;
        RECT  6.420 2.140 6.540 2.360 ;
        RECT  5.600 1.960 5.820 2.240 ;
        RECT  5.600 0.990 5.760 1.270 ;
        RECT  5.540 0.990 5.600 2.240 ;
        RECT  5.440 0.990 5.540 2.120 ;
        RECT  5.160 0.440 5.280 1.270 ;
        RECT  5.160 1.930 5.280 2.210 ;
        RECT  5.000 0.440 5.160 2.210 ;
        RECT  4.680 1.000 4.840 2.360 ;
        RECT  4.600 1.000 4.680 1.160 ;
        RECT  4.120 2.080 4.680 2.360 ;
        RECT  4.230 0.880 4.600 1.160 ;
        RECT  4.240 1.600 4.520 1.920 ;
        RECT  3.350 1.760 4.240 1.920 ;
        RECT  3.190 1.030 3.350 2.250 ;
        RECT  3.070 1.030 3.190 1.480 ;
        RECT  3.070 1.970 3.190 2.250 ;
        RECT  2.190 1.320 3.070 1.480 ;
        RECT  1.810 0.880 2.430 1.160 ;
        RECT  2.000 2.080 2.280 2.360 ;
        RECT  1.970 1.320 2.190 1.900 ;
        RECT  1.810 2.080 2.000 2.240 ;
        RECT  1.650 0.880 1.810 2.240 ;
        RECT  1.490 2.400 1.550 2.680 ;
        RECT  1.270 1.030 1.490 2.680 ;
        RECT  0.570 0.440 0.790 3.160 ;
    END
END MX4X4TR

MACRO MX4X2TR
    CLASS CORE ;
    FOREIGN MX4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.340 1.210 9.520 2.430 ;
        RECT  9.300 1.210 9.340 3.160 ;
        RECT  9.140 0.440 9.300 3.160 ;
        END
        ANTENNADIFFAREA 3.584 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.360 1.470 8.490 3.000 ;
        RECT  8.330 1.470 8.360 3.160 ;
        RECT  8.270 1.470 8.330 1.720 ;
        RECT  8.040 2.840 8.330 3.160 ;
        RECT  7.020 2.840 8.040 3.020 ;
        RECT  6.750 2.840 7.020 3.120 ;
        END
        ANTENNAGATEAREA 0.3624 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.870 2.880 5.180 3.160 ;
        RECT  3.210 2.880 4.870 3.060 ;
        RECT  4.260 0.440 4.540 0.720 ;
        RECT  3.640 0.560 4.260 0.720 ;
        RECT  3.360 0.560 3.640 0.870 ;
        RECT  2.240 0.560 3.360 0.720 ;
        RECT  3.050 2.840 3.210 3.060 ;
        RECT  1.560 2.840 3.050 3.000 ;
        RECT  1.960 0.440 2.240 0.720 ;
        RECT  1.170 0.560 1.960 0.720 ;
        RECT  1.240 2.840 1.560 3.160 ;
        RECT  1.170 2.840 1.240 3.000 ;
        RECT  1.010 0.560 1.170 3.000 ;
        END
        ANTENNAGATEAREA 0.7272 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.640 2.760 2.010 ;
        RECT  2.410 1.640 2.440 1.920 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.920 0.380 1.880 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.320 4.130 1.600 ;
        RECT  3.640 1.240 3.960 1.600 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.090 1.640 6.360 1.960 ;
        RECT  6.040 1.520 6.090 1.960 ;
        RECT  5.810 1.520 6.040 1.800 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.880 -0.280 9.600 0.280 ;
        RECT  8.600 -0.280 8.880 0.610 ;
        RECT  6.050 -0.280 8.600 0.340 ;
        RECT  3.810 -0.280 6.050 0.280 ;
        RECT  3.170 -0.280 3.810 0.390 ;
        RECT  0.370 -0.280 3.170 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.820 3.320 9.600 3.880 ;
        RECT  8.660 2.140 8.820 3.880 ;
        RECT  6.390 3.320 8.660 3.880 ;
        RECT  6.110 3.200 6.390 3.880 ;
        RECT  2.890 3.320 6.110 3.880 ;
        RECT  2.610 3.200 2.890 3.880 ;
        RECT  0.370 3.320 2.610 3.880 ;
        RECT  0.090 2.400 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.820 0.770 8.980 1.740 ;
        RECT  7.790 0.770 8.820 0.930 ;
        RECT  8.110 1.090 8.360 1.310 ;
        RECT  8.110 2.000 8.170 2.680 ;
        RECT  7.950 1.090 8.110 2.680 ;
        RECT  1.610 2.520 7.950 2.680 ;
        RECT  7.730 0.500 7.790 0.930 ;
        RECT  7.510 0.500 7.730 2.250 ;
        RECT  7.440 1.970 7.510 2.250 ;
        RECT  7.240 0.500 7.310 1.310 ;
        RECT  7.080 0.500 7.240 2.250 ;
        RECT  7.030 0.500 7.080 1.310 ;
        RECT  6.960 1.970 7.080 2.250 ;
        RECT  5.330 0.500 7.030 0.660 ;
        RECT  6.760 1.380 6.870 1.660 ;
        RECT  6.750 1.380 6.760 2.360 ;
        RECT  6.590 0.980 6.750 2.360 ;
        RECT  6.470 0.980 6.590 1.260 ;
        RECT  6.480 2.080 6.590 2.360 ;
        RECT  5.650 1.960 5.870 2.240 ;
        RECT  5.650 0.990 5.810 1.270 ;
        RECT  5.490 0.990 5.650 2.240 ;
        RECT  5.170 0.440 5.330 2.210 ;
        RECT  5.050 0.440 5.170 1.270 ;
        RECT  5.050 1.930 5.170 2.210 ;
        RECT  4.730 0.880 4.890 2.360 ;
        RECT  4.120 0.880 4.730 1.160 ;
        RECT  4.050 2.080 4.730 2.360 ;
        RECT  4.290 1.580 4.570 1.920 ;
        RECT  3.410 1.760 4.290 1.920 ;
        RECT  3.250 1.030 3.410 2.250 ;
        RECT  3.130 1.030 3.250 1.480 ;
        RECT  3.130 1.970 3.250 2.250 ;
        RECT  2.250 1.320 3.130 1.480 ;
        RECT  1.870 0.880 2.490 1.160 ;
        RECT  2.000 2.080 2.280 2.360 ;
        RECT  2.030 1.320 2.250 1.900 ;
        RECT  1.870 2.080 2.000 2.240 ;
        RECT  1.710 0.880 1.870 2.240 ;
        RECT  1.550 2.400 1.610 2.680 ;
        RECT  1.330 1.030 1.550 2.680 ;
        RECT  0.570 0.440 0.850 3.160 ;
    END
END MX4X2TR

MACRO MX4X1TR
    CLASS CORE ;
    FOREIGN MX4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.920 8.320 2.420 ;
        RECT  8.000 0.920 8.080 1.200 ;
        RECT  8.000 1.910 8.080 2.420 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 0.440 5.960 0.780 ;
        RECT  5.580 0.500 5.640 0.780 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.4272 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.200 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.500 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.240 3.580 1.620 ;
        END
        ANTENNAGATEAREA 0.1512 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.360 1.640 5.560 1.960 ;
        RECT  5.240 1.520 5.360 1.960 ;
        RECT  5.140 1.520 5.240 1.800 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.880 -0.280 8.400 0.280 ;
        RECT  7.600 -0.280 7.880 0.400 ;
        RECT  5.420 -0.280 7.600 0.280 ;
        RECT  5.140 -0.280 5.420 0.930 ;
        RECT  3.420 -0.280 5.140 0.340 ;
        RECT  3.200 -0.280 3.420 1.040 ;
        RECT  2.480 -0.280 3.200 0.280 ;
        RECT  2.200 -0.280 2.480 1.040 ;
        RECT  0.460 -0.280 2.200 0.340 ;
        RECT  0.180 -0.280 0.460 0.940 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.880 3.320 8.400 3.880 ;
        RECT  7.600 3.200 7.880 3.880 ;
        RECT  3.380 3.260 7.600 3.880 ;
        RECT  3.100 2.930 3.380 3.880 ;
        RECT  2.540 3.320 3.100 3.880 ;
        RECT  2.260 2.930 2.540 3.880 ;
        RECT  0.460 3.260 2.260 3.880 ;
        RECT  0.180 2.590 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.840 1.360 7.920 1.640 ;
        RECT  7.680 0.620 7.840 1.640 ;
        RECT  6.940 0.620 7.680 0.780 ;
        RECT  7.300 0.940 7.420 1.220 ;
        RECT  7.300 2.200 7.420 2.950 ;
        RECT  7.140 0.940 7.300 3.090 ;
        RECT  3.700 2.930 7.140 3.090 ;
        RECT  6.660 0.620 6.940 2.480 ;
        RECT  6.460 1.060 6.500 2.490 ;
        RECT  6.350 0.940 6.460 2.490 ;
        RECT  6.340 0.940 6.350 2.770 ;
        RECT  6.180 0.940 6.340 1.220 ;
        RECT  6.180 2.170 6.340 2.770 ;
        RECT  6.000 1.530 6.180 1.810 ;
        RECT  4.600 2.610 6.180 2.770 ;
        RECT  5.840 0.970 6.000 2.420 ;
        RECT  5.720 0.970 5.840 1.250 ;
        RECT  5.680 2.200 5.840 2.420 ;
        RECT  4.760 0.650 4.980 2.390 ;
        RECT  4.660 0.650 4.760 0.930 ;
        RECT  4.440 1.090 4.600 2.770 ;
        RECT  4.380 1.090 4.440 1.250 ;
        RECT  4.100 2.610 4.440 2.770 ;
        RECT  4.100 0.910 4.380 1.250 ;
        RECT  4.120 1.410 4.280 2.450 ;
        RECT  3.900 1.410 4.120 1.570 ;
        RECT  3.620 2.170 4.120 2.450 ;
        RECT  3.740 1.730 3.960 2.010 ;
        RECT  3.740 0.760 3.900 1.570 ;
        RECT  3.620 0.760 3.740 1.040 ;
        RECT  3.040 1.850 3.740 2.010 ;
        RECT  3.540 2.610 3.700 3.090 ;
        RECT  1.440 2.610 3.540 2.770 ;
        RECT  2.880 0.800 3.040 2.410 ;
        RECT  2.680 0.800 2.880 1.080 ;
        RECT  2.320 2.250 2.880 2.410 ;
        RECT  2.160 1.850 2.320 2.410 ;
        RECT  1.840 1.850 2.160 2.010 ;
        RECT  1.870 0.780 2.000 1.030 ;
        RECT  1.520 2.240 1.930 2.400 ;
        RECT  1.710 0.780 1.870 1.480 ;
        RECT  1.680 1.730 1.840 2.010 ;
        RECT  1.520 1.320 1.710 1.480 ;
        RECT  1.240 0.880 1.520 1.160 ;
        RECT  1.360 1.320 1.520 2.400 ;
        RECT  1.200 2.610 1.440 2.890 ;
        RECT  1.200 1.000 1.240 1.160 ;
        RECT  1.040 1.000 1.200 2.890 ;
        RECT  0.660 0.880 0.880 2.890 ;
    END
END MX4X1TR

MACRO MX3XLTR
    CLASS CORE ;
    FOREIGN MX3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 0.600 6.320 3.160 ;
        RECT  6.090 0.600 6.110 0.890 ;
        RECT  6.080 1.910 6.110 3.160 ;
        END
        ANTENNADIFFAREA 1.174 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.820 0.440 4.360 0.760 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.840 1.140 3.160 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.720 1.640 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.520 3.560 1.960 ;
        RECT  3.220 1.520 3.280 1.800 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.850 -0.280 6.400 0.280 ;
        RECT  5.510 -0.280 5.850 0.340 ;
        RECT  3.560 -0.280 5.510 0.280 ;
        RECT  3.280 -0.280 3.560 0.390 ;
        RECT  1.560 -0.280 3.280 0.340 ;
        RECT  1.280 -0.280 1.560 1.030 ;
        RECT  0.380 -0.280 1.280 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.900 3.320 6.400 3.880 ;
        RECT  5.620 3.000 5.900 3.880 ;
        RECT  3.640 3.320 5.620 3.880 ;
        RECT  3.360 3.260 3.640 3.880 ;
        RECT  1.520 3.320 3.360 3.880 ;
        RECT  1.300 2.780 1.520 3.880 ;
        RECT  0.380 3.320 1.300 3.880 ;
        RECT  0.100 3.200 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.870 1.370 5.950 1.650 ;
        RECT  5.710 0.670 5.870 1.650 ;
        RECT  5.080 0.670 5.710 0.830 ;
        RECT  5.520 1.030 5.550 1.420 ;
        RECT  5.400 1.030 5.520 2.530 ;
        RECT  5.360 1.030 5.400 3.100 ;
        RECT  5.220 2.250 5.360 3.100 ;
        RECT  1.840 2.940 5.220 3.100 ;
        RECT  4.960 0.670 5.080 1.390 ;
        RECT  4.910 0.670 4.960 2.660 ;
        RECT  4.800 1.040 4.910 2.660 ;
        RECT  4.680 2.160 4.800 2.660 ;
        RECT  4.480 1.140 4.640 2.000 ;
        RECT  4.320 1.140 4.480 1.300 ;
        RECT  4.320 1.840 4.480 2.780 ;
        RECT  4.140 1.460 4.320 1.680 ;
        RECT  2.740 2.560 4.320 2.780 ;
        RECT  3.860 0.920 4.140 2.360 ;
        RECT  3.060 2.080 3.120 2.360 ;
        RECT  2.900 0.760 3.060 2.360 ;
        RECT  2.590 1.060 2.740 2.780 ;
        RECT  2.580 0.820 2.590 2.780 ;
        RECT  2.340 0.820 2.580 1.220 ;
        RECT  2.240 2.500 2.580 2.780 ;
        RECT  2.260 1.380 2.420 2.300 ;
        RECT  2.060 1.380 2.260 1.540 ;
        RECT  1.760 2.140 2.260 2.300 ;
        RECT  1.880 1.700 2.100 1.980 ;
        RECT  1.880 0.800 2.060 1.540 ;
        RECT  1.120 1.820 1.880 1.980 ;
        RECT  1.680 2.460 1.840 3.100 ;
        RECT  0.800 2.460 1.680 2.620 ;
        RECT  0.960 0.490 1.120 2.220 ;
        RECT  0.720 0.490 0.960 0.770 ;
        RECT  0.840 1.940 0.960 2.220 ;
        RECT  0.680 1.030 0.800 1.310 ;
        RECT  0.680 2.460 0.800 2.680 ;
        RECT  0.520 1.030 0.680 2.680 ;
    END
END MX3XLTR

MACRO MX3X4TR
    CLASS CORE ;
    FOREIGN MX3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 0.600 7.520 3.160 ;
        RECT  7.080 0.600 7.240 0.880 ;
        RECT  7.080 2.120 7.240 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.070 1.800 6.440 2.360 ;
        RECT  6.040 1.800 6.070 2.720 ;
        RECT  5.910 2.200 6.040 2.720 ;
        RECT  4.280 2.440 5.910 2.720 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.560 3.180 2.840 ;
        RECT  2.740 2.440 2.760 2.840 ;
        RECT  2.480 2.440 2.740 2.780 ;
        RECT  2.260 0.440 2.540 0.700 ;
        RECT  1.040 2.500 2.480 2.780 ;
        RECT  1.290 0.540 2.260 0.700 ;
        RECT  1.130 0.540 1.290 0.720 ;
        RECT  1.040 1.330 1.160 1.610 ;
        RECT  1.010 0.560 1.130 0.720 ;
        RECT  1.010 1.330 1.040 2.780 ;
        RECT  0.880 0.560 1.010 2.780 ;
        RECT  0.850 0.560 0.880 1.490 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 2.040 0.720 2.360 ;
        RECT  0.480 1.600 0.690 2.360 ;
        RECT  0.470 1.600 0.480 2.070 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 2.050 1.580 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.070 1.240 4.360 1.560 ;
        RECT  4.040 1.240 4.070 1.580 ;
        RECT  3.790 1.300 4.040 1.580 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.910 -0.280 8.000 0.280 ;
        RECT  7.680 -0.280 7.910 1.310 ;
        RECT  6.880 -0.280 7.680 0.280 ;
        RECT  6.600 -0.280 6.880 0.670 ;
        RECT  4.030 -0.280 6.600 0.340 ;
        RECT  1.770 -0.280 4.030 0.280 ;
        RECT  1.490 -0.280 1.770 0.380 ;
        RECT  0.970 -0.280 1.490 0.340 ;
        RECT  0.690 -0.280 0.970 0.400 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.910 3.320 8.000 3.880 ;
        RECT  7.680 1.910 7.910 3.880 ;
        RECT  6.880 3.320 7.680 3.880 ;
        RECT  6.600 2.910 6.880 3.880 ;
        RECT  4.110 3.260 6.600 3.880 ;
        RECT  1.780 3.320 4.110 3.880 ;
        RECT  0.650 3.260 1.780 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.920 1.040 7.080 1.960 ;
        RECT  6.390 1.040 6.920 1.200 ;
        RECT  6.760 1.800 6.920 1.960 ;
        RECT  6.480 1.360 6.760 1.640 ;
        RECT  6.600 1.800 6.760 2.680 ;
        RECT  6.390 2.520 6.600 2.680 ;
        RECT  5.750 1.480 6.480 1.640 ;
        RECT  6.110 0.500 6.390 1.200 ;
        RECT  6.230 2.520 6.390 3.100 ;
        RECT  3.500 2.880 6.230 3.100 ;
        RECT  5.670 0.500 5.790 1.270 ;
        RECT  5.670 1.480 5.750 2.210 ;
        RECT  5.510 0.500 5.670 2.210 ;
        RECT  5.470 1.480 5.510 2.210 ;
        RECT  5.030 0.500 5.310 2.210 ;
        RECT  3.250 0.500 5.030 0.660 ;
        RECT  4.990 1.930 5.030 2.210 ;
        RECT  4.750 1.260 4.870 1.540 ;
        RECT  4.590 0.860 4.750 2.210 ;
        RECT  4.470 0.860 4.590 1.080 ;
        RECT  4.470 1.930 4.590 2.210 ;
        RECT  3.630 1.930 3.870 2.720 ;
        RECT  3.630 0.860 3.750 1.140 ;
        RECT  3.470 0.860 3.630 2.720 ;
        RECT  3.340 2.880 3.500 3.160 ;
        RECT  2.100 3.000 3.340 3.160 ;
        RECT  3.130 0.500 3.250 1.250 ;
        RECT  3.130 1.930 3.250 2.210 ;
        RECT  2.970 0.500 3.130 2.210 ;
        RECT  2.650 0.860 2.810 2.220 ;
        RECT  2.050 0.860 2.650 1.080 ;
        RECT  2.300 2.060 2.650 2.220 ;
        RECT  2.210 1.580 2.490 1.900 ;
        RECT  2.020 2.060 2.300 2.340 ;
        RECT  1.480 1.740 2.210 1.900 ;
        RECT  1.940 2.940 2.100 3.160 ;
        RECT  0.310 2.940 1.940 3.100 ;
        RECT  1.420 0.890 1.480 1.930 ;
        RECT  1.320 0.890 1.420 2.210 ;
        RECT  1.170 0.890 1.320 1.170 ;
        RECT  1.200 1.770 1.320 2.210 ;
        RECT  0.310 0.440 0.410 1.310 ;
        RECT  0.090 0.440 0.310 3.100 ;
    END
END MX3X4TR

MACRO MX3X2TR
    CLASS CORE ;
    FOREIGN MX3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.360 0.540 7.520 3.160 ;
        RECT  6.980 0.540 7.360 0.820 ;
        RECT  6.980 2.040 7.360 3.160 ;
        END
        ANTENNADIFFAREA 3.424 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.360 1.740 6.370 2.020 ;
        RECT  6.040 1.740 6.360 2.360 ;
        RECT  6.000 2.200 6.040 2.360 ;
        RECT  5.840 2.200 6.000 2.660 ;
        RECT  4.230 2.470 5.840 2.660 ;
        END
        ANTENNAGATEAREA 0.3336 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 2.440 3.160 2.840 ;
        RECT  2.840 2.440 2.850 2.780 ;
        RECT  1.040 2.500 2.840 2.780 ;
        RECT  2.210 0.440 2.490 0.700 ;
        RECT  1.280 0.540 2.210 0.700 ;
        RECT  1.120 0.540 1.280 0.720 ;
        RECT  1.040 1.330 1.160 1.610 ;
        RECT  0.920 0.560 1.120 0.720 ;
        RECT  0.920 1.330 1.040 2.780 ;
        RECT  0.880 0.560 0.920 2.780 ;
        RECT  0.760 0.560 0.880 1.490 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.790 0.720 2.360 ;
        RECT  0.440 1.790 0.480 2.070 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 2.080 1.580 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.040 1.240 4.360 1.560 ;
        RECT  3.760 1.300 4.040 1.580 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.780 -0.280 7.600 0.280 ;
        RECT  6.500 -0.280 6.780 0.670 ;
        RECT  4.000 -0.280 6.500 0.340 ;
        RECT  1.760 -0.280 4.000 0.280 ;
        RECT  1.480 -0.280 1.760 0.380 ;
        RECT  0.960 -0.280 1.480 0.340 ;
        RECT  0.680 -0.280 0.960 0.400 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.780 3.320 7.600 3.880 ;
        RECT  6.500 2.910 6.780 3.880 ;
        RECT  4.340 3.260 6.500 3.880 ;
        RECT  4.060 3.200 4.340 3.880 ;
        RECT  1.840 3.320 4.060 3.880 ;
        RECT  0.690 3.260 1.840 3.880 ;
        RECT  0.000 3.320 0.690 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.040 0.980 7.200 1.880 ;
        RECT  6.320 0.980 7.040 1.140 ;
        RECT  6.690 1.720 7.040 1.880 ;
        RECT  6.600 1.300 6.880 1.560 ;
        RECT  6.530 1.720 6.690 2.680 ;
        RECT  5.840 1.400 6.600 1.560 ;
        RECT  6.320 2.520 6.530 2.680 ;
        RECT  6.040 0.520 6.320 1.240 ;
        RECT  6.160 2.520 6.320 3.040 ;
        RECT  3.480 2.820 6.160 3.040 ;
        RECT  5.680 0.520 5.840 1.560 ;
        RECT  5.560 0.520 5.680 2.280 ;
        RECT  5.520 1.420 5.560 2.280 ;
        RECT  5.400 1.990 5.520 2.280 ;
        RECT  5.240 0.500 5.360 1.220 ;
        RECT  5.080 0.500 5.240 2.200 ;
        RECT  3.280 0.500 5.080 0.660 ;
        RECT  4.920 1.920 5.080 2.200 ;
        RECT  4.740 1.250 4.920 1.530 ;
        RECT  4.580 0.820 4.740 2.200 ;
        RECT  4.460 0.820 4.580 1.100 ;
        RECT  4.430 1.920 4.580 2.200 ;
        RECT  3.600 1.920 3.820 2.660 ;
        RECT  3.600 0.860 3.760 1.140 ;
        RECT  3.440 0.860 3.600 2.660 ;
        RECT  3.320 2.820 3.480 3.160 ;
        RECT  2.140 3.000 3.320 3.160 ;
        RECT  3.160 0.500 3.280 1.250 ;
        RECT  3.160 1.920 3.280 2.200 ;
        RECT  3.000 0.500 3.160 2.200 ;
        RECT  2.680 0.860 2.840 2.220 ;
        RECT  2.000 0.860 2.680 1.080 ;
        RECT  2.360 2.060 2.680 2.220 ;
        RECT  2.240 1.570 2.520 1.900 ;
        RECT  2.080 2.060 2.360 2.340 ;
        RECT  1.480 1.740 2.240 1.900 ;
        RECT  2.000 2.940 2.140 3.160 ;
        RECT  0.320 2.940 2.000 3.100 ;
        RECT  1.360 1.010 1.480 2.200 ;
        RECT  1.320 0.890 1.360 2.200 ;
        RECT  1.080 0.890 1.320 1.170 ;
        RECT  1.200 1.770 1.320 2.200 ;
        RECT  0.280 0.570 0.440 1.310 ;
        RECT  0.280 2.190 0.320 3.100 ;
        RECT  0.120 0.570 0.280 3.100 ;
        RECT  0.100 2.190 0.120 3.100 ;
    END
END MX3X2TR

MACRO MX3X1TR
    CLASS CORE ;
    FOREIGN MX3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 0.530 6.320 3.160 ;
        RECT  6.090 0.530 6.110 0.840 ;
        RECT  6.080 1.910 6.110 3.160 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.440 4.360 0.760 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.840 1.140 3.160 ;
        END
        ANTENNAGATEAREA 0.2232 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.720 1.640 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.520 3.560 1.960 ;
        RECT  3.220 1.520 3.280 1.800 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.790 -0.280 6.400 0.280 ;
        RECT  5.510 -0.280 5.790 0.510 ;
        RECT  3.600 -0.280 5.510 0.280 ;
        RECT  3.280 -0.280 3.600 0.870 ;
        RECT  1.560 -0.280 3.280 0.340 ;
        RECT  1.280 -0.280 1.560 1.030 ;
        RECT  0.380 -0.280 1.280 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.900 3.320 6.400 3.880 ;
        RECT  5.620 3.000 5.900 3.880 ;
        RECT  3.640 3.320 5.620 3.880 ;
        RECT  3.360 3.260 3.640 3.880 ;
        RECT  1.520 3.320 3.360 3.880 ;
        RECT  1.300 2.780 1.520 3.880 ;
        RECT  0.380 3.320 1.300 3.880 ;
        RECT  0.100 3.200 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.870 1.370 5.950 1.650 ;
        RECT  5.710 0.670 5.870 1.650 ;
        RECT  5.080 0.670 5.710 0.830 ;
        RECT  5.520 1.030 5.550 1.420 ;
        RECT  5.400 1.030 5.520 2.530 ;
        RECT  5.360 1.030 5.400 3.100 ;
        RECT  5.220 2.250 5.360 3.100 ;
        RECT  1.840 2.940 5.220 3.100 ;
        RECT  4.960 0.670 5.080 1.220 ;
        RECT  4.800 0.670 4.960 2.440 ;
        RECT  4.680 2.160 4.800 2.440 ;
        RECT  4.480 0.960 4.640 2.000 ;
        RECT  4.320 0.960 4.480 1.240 ;
        RECT  4.320 1.840 4.480 2.780 ;
        RECT  4.140 1.400 4.320 1.680 ;
        RECT  2.740 2.560 4.320 2.780 ;
        RECT  3.860 0.920 4.140 2.360 ;
        RECT  3.060 2.080 3.120 2.360 ;
        RECT  2.900 0.620 3.060 2.360 ;
        RECT  2.780 0.620 2.900 0.900 ;
        RECT  2.580 1.060 2.740 2.780 ;
        RECT  2.520 1.060 2.580 1.220 ;
        RECT  2.240 2.500 2.580 2.780 ;
        RECT  2.240 0.820 2.520 1.220 ;
        RECT  2.260 1.380 2.420 2.300 ;
        RECT  2.040 1.380 2.260 1.540 ;
        RECT  1.760 2.140 2.260 2.300 ;
        RECT  1.880 1.700 2.100 1.980 ;
        RECT  1.880 0.800 2.040 1.540 ;
        RECT  1.760 0.800 1.880 1.080 ;
        RECT  1.120 1.820 1.880 1.980 ;
        RECT  1.680 2.460 1.840 3.100 ;
        RECT  0.800 2.460 1.680 2.620 ;
        RECT  0.960 0.490 1.120 2.220 ;
        RECT  0.720 0.490 0.960 0.770 ;
        RECT  0.840 1.940 0.960 2.220 ;
        RECT  0.680 1.030 0.800 1.310 ;
        RECT  0.680 2.460 0.800 2.680 ;
        RECT  0.520 1.030 0.680 2.680 ;
    END
END MX3X1TR

MACRO MX2XLTR
    CLASS CORE ;
    FOREIGN MX2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.480 3.520 3.080 ;
        RECT  3.140 0.480 3.360 0.760 ;
        RECT  3.280 2.120 3.360 3.080 ;
        RECT  3.240 2.440 3.280 3.080 ;
        END
        ANTENNADIFFAREA 1.612 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 2.440 0.720 2.840 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.640 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.160 1.750 ;
        RECT  2.610 1.470 2.840 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.960 -0.280 3.600 0.280 ;
        RECT  2.680 -0.280 2.960 0.800 ;
        RECT  0.930 -0.280 2.680 0.340 ;
        RECT  0.650 -0.280 0.930 0.800 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.080 3.320 3.600 3.880 ;
        RECT  2.800 3.200 3.080 3.880 ;
        RECT  1.040 3.320 2.800 3.880 ;
        RECT  0.880 2.880 1.040 3.880 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.770 1.960 3.110 2.240 ;
        RECT  2.610 1.960 2.770 2.890 ;
        RECT  2.080 2.730 2.610 2.890 ;
        RECT  2.450 1.030 2.510 1.310 ;
        RECT  2.240 1.030 2.450 2.570 ;
        RECT  1.920 0.520 2.080 2.890 ;
        RECT  1.670 0.520 1.920 0.800 ;
        RECT  1.810 2.730 1.920 2.890 ;
        RECT  1.530 2.730 1.810 3.160 ;
        RECT  1.600 1.000 1.760 2.450 ;
        RECT  1.390 1.000 1.600 1.160 ;
        RECT  1.370 2.290 1.600 2.450 ;
        RECT  1.280 1.320 1.440 1.980 ;
        RECT  1.110 0.880 1.390 1.160 ;
        RECT  1.090 2.290 1.370 2.570 ;
        RECT  0.370 1.320 1.280 1.480 ;
        RECT  0.320 1.030 0.370 1.480 ;
        RECT  0.160 1.030 0.320 2.280 ;
        RECT  0.090 1.030 0.160 1.310 ;
        RECT  0.090 2.000 0.160 2.280 ;
    END
END MX2XLTR

MACRO MX2X8TR
    CLASS CORE ;
    FOREIGN MX2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.440 6.120 2.170 ;
        RECT  5.800 0.520 5.850 2.170 ;
        RECT  5.540 0.520 5.800 3.090 ;
        RECT  5.500 0.520 5.540 2.570 ;
        RECT  5.370 0.870 5.500 2.570 ;
        RECT  4.790 0.870 5.370 1.280 ;
        RECT  4.780 2.090 5.370 2.570 ;
        RECT  4.500 0.480 4.790 1.280 ;
        RECT  4.500 2.090 4.780 3.090 ;
        END
        ANTENNADIFFAREA 8.018 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 2.710 0.720 3.160 ;
        END
        ANTENNAGATEAREA 0.3432 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.600 1.280 1.790 ;
        RECT  0.820 1.600 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.860 1.240 4.320 1.600 ;
        END
        ANTENNAGATEAREA 0.2448 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.280 -0.280 6.400 0.280 ;
        RECT  6.010 -0.280 6.280 1.100 ;
        RECT  5.300 -0.280 6.010 0.280 ;
        RECT  5.020 -0.280 5.300 0.660 ;
        RECT  4.260 -0.280 5.020 0.280 ;
        RECT  3.980 -0.280 4.260 0.940 ;
        RECT  2.060 -0.280 3.980 0.280 ;
        RECT  1.780 -0.280 2.060 0.800 ;
        RECT  0.980 -0.280 1.780 0.280 ;
        RECT  0.700 -0.280 0.980 1.090 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.260 3.320 6.400 3.880 ;
        RECT  6.000 2.510 6.260 3.880 ;
        RECT  5.300 3.320 6.000 3.880 ;
        RECT  5.020 2.890 5.300 3.880 ;
        RECT  4.260 3.320 5.020 3.880 ;
        RECT  3.980 2.760 4.260 3.880 ;
        RECT  1.770 3.320 3.980 3.880 ;
        RECT  1.800 2.010 1.960 2.430 ;
        RECT  1.770 2.270 1.800 2.430 ;
        RECT  1.610 2.270 1.770 3.880 ;
        RECT  1.090 3.320 1.610 3.880 ;
        RECT  0.910 2.250 1.090 3.880 ;
        RECT  0.700 2.250 0.910 2.520 ;
        RECT  0.000 3.320 0.910 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.800 1.520 5.190 1.800 ;
        RECT  4.550 1.520 4.800 1.920 ;
        RECT  4.090 1.760 4.550 1.920 ;
        RECT  3.930 1.760 4.090 2.530 ;
        RECT  3.360 2.370 3.930 2.530 ;
        RECT  3.520 0.460 3.680 2.210 ;
        RECT  3.230 0.690 3.360 2.530 ;
        RECT  3.200 0.690 3.230 2.890 ;
        RECT  3.160 0.690 3.200 0.850 ;
        RECT  2.980 2.260 3.200 2.890 ;
        RECT  2.880 0.570 3.160 0.850 ;
        RECT  2.880 1.010 3.040 2.100 ;
        RECT  2.170 2.590 2.980 2.750 ;
        RECT  2.580 1.010 2.880 1.170 ;
        RECT  2.640 1.940 2.880 2.100 ;
        RECT  2.600 1.610 2.720 1.770 ;
        RECT  2.360 1.940 2.640 2.220 ;
        RECT  2.440 1.330 2.600 1.770 ;
        RECT  2.300 0.490 2.580 1.170 ;
        RECT  1.640 1.330 2.440 1.490 ;
        RECT  2.280 1.940 2.360 2.100 ;
        RECT  1.500 0.960 2.300 1.120 ;
        RECT  2.120 1.650 2.280 2.100 ;
        RECT  1.950 2.590 2.170 2.880 ;
        RECT  1.640 1.650 2.120 1.810 ;
        RECT  1.480 1.280 1.640 1.490 ;
        RECT  1.480 1.650 1.640 2.110 ;
        RECT  1.220 0.810 1.500 1.120 ;
        RECT  0.370 1.280 1.480 1.440 ;
        RECT  1.440 1.950 1.480 2.110 ;
        RECT  1.280 1.950 1.440 2.790 ;
        RECT  0.140 0.800 0.370 2.440 ;
        RECT  0.100 0.800 0.140 1.130 ;
        RECT  0.100 2.160 0.140 2.440 ;
    END
END MX2X8TR

MACRO MX2X6TR
    CLASS CORE ;
    FOREIGN MX2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.580 0.540 5.860 3.090 ;
        RECT  5.050 1.000 5.580 2.440 ;
        RECT  4.830 1.000 5.050 1.360 ;
        RECT  4.830 2.080 5.050 2.440 ;
        RECT  4.540 0.530 4.830 1.360 ;
        RECT  4.530 2.080 4.830 3.040 ;
        END
        ANTENNADIFFAREA 8.14 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 2.840 0.720 3.160 ;
        RECT  0.410 2.710 0.570 3.160 ;
        END
        ANTENNAGATEAREA 0.3528 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.600 1.320 1.790 ;
        RECT  0.880 1.600 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.900 1.240 4.320 1.600 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.350 -0.280 6.000 0.280 ;
        RECT  5.060 -0.280 5.350 0.720 ;
        RECT  4.300 -0.280 5.060 0.290 ;
        RECT  4.020 -0.280 4.300 0.970 ;
        RECT  2.060 -0.280 4.020 0.290 ;
        RECT  1.780 -0.280 2.060 0.800 ;
        RECT  0.980 -0.280 1.780 0.290 ;
        RECT  0.700 -0.280 0.980 1.060 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.340 3.320 6.000 3.880 ;
        RECT  5.060 2.750 5.340 3.880 ;
        RECT  4.300 3.320 5.060 3.880 ;
        RECT  4.020 2.690 4.300 3.880 ;
        RECT  1.760 3.320 4.020 3.880 ;
        RECT  1.800 2.070 1.960 2.430 ;
        RECT  1.760 2.270 1.800 2.430 ;
        RECT  1.600 2.270 1.760 3.880 ;
        RECT  1.050 3.320 1.600 3.880 ;
        RECT  0.880 2.250 1.050 3.880 ;
        RECT  0.640 2.250 0.880 2.410 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.480 1.520 4.640 1.920 ;
        RECT  4.130 1.760 4.480 1.920 ;
        RECT  3.970 1.760 4.130 2.530 ;
        RECT  3.400 2.370 3.970 2.530 ;
        RECT  3.560 0.530 3.720 2.210 ;
        RECT  3.240 0.590 3.400 2.530 ;
        RECT  2.920 0.590 3.240 0.750 ;
        RECT  3.200 2.370 3.240 2.530 ;
        RECT  2.920 2.370 3.200 2.910 ;
        RECT  2.920 0.960 3.080 2.210 ;
        RECT  2.560 0.960 2.920 1.120 ;
        RECT  2.680 2.050 2.920 2.210 ;
        RECT  2.080 2.750 2.920 2.910 ;
        RECT  2.620 1.660 2.740 1.820 ;
        RECT  2.400 2.050 2.680 2.560 ;
        RECT  2.460 1.280 2.620 1.820 ;
        RECT  2.280 0.560 2.560 1.120 ;
        RECT  0.380 1.280 2.460 1.440 ;
        RECT  2.300 2.050 2.400 2.210 ;
        RECT  2.140 1.720 2.300 2.210 ;
        RECT  1.500 0.960 2.280 1.120 ;
        RECT  1.640 1.720 2.140 1.880 ;
        RECT  1.920 2.590 2.080 2.910 ;
        RECT  1.480 1.720 1.640 2.110 ;
        RECT  1.220 0.840 1.500 1.120 ;
        RECT  1.440 1.950 1.480 2.110 ;
        RECT  1.280 1.950 1.440 2.820 ;
        RECT  1.220 2.480 1.280 2.820 ;
        RECT  0.220 0.800 0.380 2.390 ;
        RECT  0.100 0.800 0.220 1.130 ;
        RECT  0.100 2.080 0.220 2.390 ;
    END
END MX2X6TR

MACRO MX2X4TR
    CLASS CORE ;
    FOREIGN MX2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.470 0.840 4.670 2.290 ;
        RECT  4.200 0.840 4.470 1.060 ;
        RECT  4.320 2.090 4.470 2.290 ;
        RECT  4.200 2.090 4.320 2.980 ;
        RECT  3.920 0.550 4.200 1.060 ;
        RECT  3.920 2.090 4.200 3.090 ;
        END
        ANTENNADIFFAREA 4.2 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 2.980 2.400 3.160 ;
        RECT  2.130 0.440 2.280 2.360 ;
        RECT  2.120 0.440 2.130 3.160 ;
        RECT  1.450 0.440 2.120 0.620 ;
        RECT  1.970 2.200 2.120 3.160 ;
        RECT  1.680 2.730 1.970 3.160 ;
        RECT  0.530 2.730 1.680 2.910 ;
        RECT  0.230 2.730 0.530 2.980 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.600 1.110 1.780 ;
        RECT  0.480 1.600 0.800 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.240 3.750 1.560 ;
        RECT  3.260 1.240 3.500 1.600 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.280 4.800 0.280 ;
        RECT  4.420 -0.280 4.700 0.660 ;
        RECT  3.700 -0.280 4.420 0.280 ;
        RECT  3.420 -0.280 3.700 0.940 ;
        RECT  0.970 -0.280 3.420 0.280 ;
        RECT  0.700 -0.280 0.970 0.400 ;
        RECT  0.000 -0.280 0.700 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.480 2.450 4.700 3.880 ;
        RECT  3.700 3.320 4.480 3.880 ;
        RECT  3.420 2.970 3.700 3.880 ;
        RECT  1.020 3.320 3.420 3.880 ;
        RECT  0.660 3.200 1.020 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.940 1.520 4.120 1.920 ;
        RECT  3.600 1.760 3.940 1.920 ;
        RECT  3.440 1.760 3.600 2.750 ;
        RECT  2.600 2.590 3.440 2.750 ;
        RECT  3.100 1.990 3.200 2.290 ;
        RECT  2.940 0.530 3.100 2.290 ;
        RECT  2.890 1.980 2.940 2.290 ;
        RECT  2.440 0.530 2.600 2.750 ;
        RECT  2.310 2.520 2.440 2.750 ;
        RECT  1.800 0.960 1.960 2.040 ;
        RECT  1.700 0.960 1.800 1.120 ;
        RECT  1.480 1.880 1.800 2.040 ;
        RECT  1.420 0.830 1.700 1.120 ;
        RECT  1.560 1.400 1.640 1.700 ;
        RECT  1.400 1.280 1.560 1.700 ;
        RECT  1.320 1.880 1.480 2.390 ;
        RECT  0.420 1.280 1.400 1.440 ;
        RECT  0.320 0.900 0.420 1.440 ;
        RECT  0.160 0.900 0.320 2.440 ;
        RECT  0.140 0.900 0.160 1.280 ;
    END
END MX2X4TR

MACRO MX2X2TR
    CLASS CORE ;
    FOREIGN MX2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.240 3.920 2.360 ;
        RECT  3.820 1.240 3.880 3.160 ;
        RECT  3.660 0.500 3.820 3.160 ;
        END
        ANTENNADIFFAREA 4.364 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.230 1.700 1.590 ;
        RECT  1.090 1.230 1.540 1.450 ;
        RECT  0.930 0.570 1.090 1.450 ;
        RECT  0.260 0.570 0.930 0.740 ;
        RECT  0.470 2.780 0.770 3.160 ;
        RECT  0.260 2.780 0.470 2.960 ;
        RECT  0.100 0.570 0.260 2.960 ;
        END
        ANTENNAGATEAREA 0.2928 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.640 1.350 1.810 ;
        RECT  0.880 1.640 1.160 2.150 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.120 1.670 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.280 4.000 0.280 ;
        RECT  2.970 -0.280 3.270 0.410 ;
        RECT  0.000 -0.280 2.970 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.300 3.320 4.000 3.880 ;
        RECT  3.020 3.200 3.300 3.880 ;
        RECT  1.290 3.260 3.020 3.880 ;
        RECT  1.010 2.670 1.290 3.880 ;
        RECT  0.000 3.320 1.010 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.280 0.570 3.440 3.040 ;
        RECT  2.120 0.570 3.280 0.730 ;
        RECT  2.280 2.880 3.280 3.040 ;
        RECT  2.660 1.910 2.780 2.720 ;
        RECT  2.500 0.890 2.660 2.720 ;
        RECT  2.180 1.200 2.340 2.510 ;
        RECT  2.000 2.670 2.280 3.040 ;
        RECT  0.690 2.350 2.180 2.510 ;
        RECT  1.840 0.450 2.120 0.730 ;
        RECT  1.860 0.890 2.020 2.150 ;
        RECT  1.640 0.890 1.860 1.050 ;
        RECT  1.470 1.990 1.860 2.150 ;
        RECT  1.360 0.770 1.640 1.050 ;
        RECT  0.530 0.900 0.690 2.510 ;
        RECT  0.420 0.900 0.530 1.210 ;
    END
END MX2X2TR

MACRO MX2X1TR
    CLASS CORE ;
    FOREIGN MX2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.440 3.520 2.900 ;
        RECT  3.280 0.440 3.360 1.560 ;
        RECT  3.220 2.480 3.360 2.900 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 2.840 0.720 3.160 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.950 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.680 1.240 3.120 1.650 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.280 3.600 0.280 ;
        RECT  2.690 -0.280 2.970 0.400 ;
        RECT  0.960 -0.280 2.690 0.280 ;
        RECT  0.680 -0.280 0.960 1.150 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 3.320 3.600 3.880 ;
        RECT  2.690 3.200 2.970 3.880 ;
        RECT  1.080 3.320 2.690 3.880 ;
        RECT  0.880 2.520 1.080 3.880 ;
        RECT  0.790 2.520 0.880 2.680 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.060 1.890 3.200 2.210 ;
        RECT  2.900 1.890 3.060 2.900 ;
        RECT  2.140 2.740 2.900 2.900 ;
        RECT  2.300 0.950 2.520 2.580 ;
        RECT  1.980 0.870 2.140 2.900 ;
        RECT  1.640 0.870 1.980 1.150 ;
        RECT  1.760 2.390 1.980 2.670 ;
        RECT  1.660 1.310 1.820 2.230 ;
        RECT  1.440 1.310 1.660 1.470 ;
        RECT  1.560 2.070 1.660 2.230 ;
        RECT  1.400 2.070 1.560 2.590 ;
        RECT  1.280 1.630 1.500 1.910 ;
        RECT  1.160 0.950 1.440 1.470 ;
        RECT  1.280 2.310 1.400 2.590 ;
        RECT  0.340 1.630 1.280 1.790 ;
        RECT  0.340 2.400 0.390 2.680 ;
        RECT  0.180 1.030 0.340 2.680 ;
        RECT  0.120 2.400 0.180 2.680 ;
    END
END MX2X1TR

MACRO MDFFHQX8TR
    CLASS CORE ;
    FOREIGN MDFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.350 2.370 1.630 ;
        RECT  1.680 1.240 1.960 1.630 ;
        END
        ANTENNAGATEAREA 0.5616 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.540 0.440 15.820 3.160 ;
        RECT  14.960 1.250 15.540 1.730 ;
        RECT  14.860 1.250 14.960 2.560 ;
        RECT  14.580 0.440 14.860 3.160 ;
        RECT  14.240 1.720 14.580 2.560 ;
        END
        ANTENNADIFFAREA 7.956 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.440 0.560 1.670 ;
        RECT  0.080 0.840 0.330 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.150 1.230 5.660 1.560 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.300 -0.280 16.400 0.280 ;
        RECT  16.020 -0.280 16.300 1.210 ;
        RECT  15.340 -0.280 16.020 0.280 ;
        RECT  15.060 -0.280 15.340 1.090 ;
        RECT  14.380 -0.280 15.060 0.280 ;
        RECT  14.100 -0.280 14.380 1.250 ;
        RECT  9.890 -0.280 14.100 0.340 ;
        RECT  9.610 -0.280 9.890 0.400 ;
        RECT  8.570 -0.280 9.610 0.340 ;
        RECT  7.130 -0.280 8.570 0.280 ;
        RECT  6.850 -0.280 7.130 0.610 ;
        RECT  5.630 -0.280 6.850 0.280 ;
        RECT  5.350 -0.280 5.630 0.670 ;
        RECT  4.170 -0.280 5.350 0.280 ;
        RECT  3.890 -0.280 4.170 0.360 ;
        RECT  2.750 -0.280 3.890 0.280 ;
        RECT  2.470 -0.280 2.750 0.360 ;
        RECT  1.710 -0.280 2.470 0.340 ;
        RECT  1.430 -0.280 1.710 0.400 ;
        RECT  0.370 -0.280 1.430 0.280 ;
        RECT  0.090 -0.280 0.370 0.680 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.300 3.320 16.400 3.880 ;
        RECT  16.000 2.070 16.300 3.880 ;
        RECT  15.350 3.320 16.000 3.880 ;
        RECT  15.120 2.090 15.350 3.880 ;
        RECT  14.380 3.320 15.120 3.880 ;
        RECT  14.090 2.790 14.380 3.880 ;
        RECT  13.650 3.320 14.090 3.880 ;
        RECT  13.370 3.200 13.650 3.880 ;
        RECT  10.930 3.260 13.370 3.880 ;
        RECT  10.650 3.200 10.930 3.880 ;
        RECT  9.890 3.320 10.650 3.880 ;
        RECT  9.610 3.200 9.890 3.880 ;
        RECT  8.780 3.260 9.610 3.880 ;
        RECT  8.500 3.200 8.780 3.880 ;
        RECT  7.090 3.320 8.500 3.880 ;
        RECT  6.810 3.200 7.090 3.880 ;
        RECT  6.050 3.320 6.810 3.880 ;
        RECT  5.770 3.200 6.050 3.880 ;
        RECT  4.210 3.320 5.770 3.880 ;
        RECT  3.930 3.200 4.210 3.880 ;
        RECT  2.750 3.320 3.930 3.880 ;
        RECT  2.470 3.200 2.750 3.880 ;
        RECT  1.710 3.260 2.470 3.880 ;
        RECT  1.430 3.200 1.710 3.880 ;
        RECT  0.370 3.320 1.430 3.880 ;
        RECT  0.090 2.430 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.710 0.860 13.920 1.160 ;
        RECT  13.710 2.350 13.920 2.630 ;
        RECT  13.550 0.860 13.710 2.630 ;
        RECT  13.410 1.680 13.550 1.960 ;
        RECT  13.250 1.240 13.390 1.520 ;
        RECT  13.090 0.660 13.250 2.620 ;
        RECT  12.230 0.660 13.090 0.820 ;
        RECT  12.150 2.400 13.090 2.620 ;
        RECT  12.770 0.980 12.930 2.240 ;
        RECT  11.750 0.980 12.770 1.140 ;
        RECT  11.950 2.080 12.770 2.240 ;
        RECT  12.360 2.820 12.640 3.100 ;
        RECT  12.390 1.360 12.610 1.920 ;
        RECT  10.530 1.360 12.390 1.520 ;
        RECT  8.460 2.820 12.360 2.980 ;
        RECT  11.950 0.540 12.230 0.820 ;
        RECT  11.470 2.400 12.150 2.560 ;
        RECT  11.270 0.540 11.950 0.700 ;
        RECT  11.670 1.850 11.950 2.240 ;
        RECT  11.470 0.860 11.750 1.140 ;
        RECT  10.410 1.850 11.670 2.010 ;
        RECT  10.850 0.980 11.470 1.140 ;
        RECT  11.190 2.220 11.470 2.560 ;
        RECT  11.050 0.540 11.270 0.820 ;
        RECT  10.690 0.680 10.850 1.140 ;
        RECT  10.410 0.680 10.690 0.840 ;
        RECT  10.370 1.000 10.530 1.520 ;
        RECT  10.130 0.590 10.410 0.840 ;
        RECT  10.130 1.850 10.410 2.660 ;
        RECT  9.570 1.000 10.370 1.160 ;
        RECT  9.930 1.320 10.210 1.600 ;
        RECT  9.720 2.350 10.130 2.510 ;
        RECT  9.250 1.440 9.930 1.600 ;
        RECT  9.440 2.350 9.720 2.630 ;
        RECT  9.410 0.710 9.570 1.160 ;
        RECT  9.130 0.590 9.410 0.870 ;
        RECT  9.090 1.030 9.250 2.190 ;
        RECT  7.530 0.710 9.130 0.870 ;
        RECT  7.690 1.030 9.090 1.250 ;
        RECT  7.660 1.910 9.090 2.190 ;
        RECT  8.650 1.470 8.930 1.750 ;
        RECT  7.500 1.590 8.650 1.750 ;
        RECT  8.300 2.500 8.460 2.980 ;
        RECT  7.500 2.500 8.300 2.700 ;
        RECT  3.210 2.860 8.140 3.040 ;
        RECT  7.350 0.710 7.530 0.930 ;
        RECT  7.340 1.180 7.500 2.700 ;
        RECT  6.690 0.770 7.350 0.930 ;
        RECT  7.050 1.180 7.340 1.340 ;
        RECT  4.560 2.540 7.340 2.700 ;
        RECT  6.690 1.520 7.180 1.800 ;
        RECT  6.570 0.770 6.690 2.220 ;
        RECT  6.530 0.530 6.570 2.280 ;
        RECT  6.290 0.530 6.530 1.250 ;
        RECT  6.290 2.060 6.530 2.280 ;
        RECT  6.130 1.620 6.370 1.900 ;
        RECT  5.320 2.060 6.290 2.220 ;
        RECT  6.090 0.650 6.130 1.900 ;
        RECT  5.970 0.650 6.090 1.880 ;
        RECT  5.830 0.650 5.970 0.930 ;
        RECT  4.880 1.720 5.970 1.880 ;
        RECT  5.040 2.060 5.320 2.300 ;
        RECT  5.030 0.590 5.150 0.870 ;
        RECT  4.870 0.590 5.030 1.070 ;
        RECT  4.720 1.720 4.880 2.000 ;
        RECT  4.560 0.910 4.870 1.070 ;
        RECT  4.410 0.470 4.690 0.750 ;
        RECT  4.400 0.910 4.560 2.700 ;
        RECT  4.240 0.590 4.410 0.750 ;
        RECT  4.080 0.590 4.240 2.090 ;
        RECT  3.650 0.590 4.080 0.750 ;
        RECT  3.690 1.930 4.080 2.090 ;
        RECT  3.410 1.930 3.690 2.660 ;
        RECT  3.430 0.470 3.650 0.750 ;
        RECT  3.210 0.820 3.240 2.040 ;
        RECT  3.080 0.820 3.210 3.040 ;
        RECT  2.850 0.820 3.080 1.100 ;
        RECT  2.930 1.930 3.080 3.040 ;
        RECT  1.370 2.440 2.930 2.600 ;
        RECT  2.690 1.260 2.920 1.540 ;
        RECT  2.530 0.920 2.690 1.950 ;
        RECT  2.280 0.920 2.530 1.080 ;
        RECT  2.230 1.790 2.530 1.950 ;
        RECT  1.950 0.800 2.280 1.080 ;
        RECT  1.950 1.790 2.230 2.280 ;
        RECT  1.520 1.790 1.950 1.950 ;
        RECT  1.360 1.670 1.520 1.950 ;
        RECT  1.200 1.000 1.370 1.280 ;
        RECT  1.200 2.320 1.370 2.600 ;
        RECT  1.040 1.000 1.200 2.600 ;
        RECT  0.720 0.440 0.880 3.160 ;
        RECT  0.610 0.440 0.720 1.280 ;
        RECT  0.610 1.940 0.720 3.160 ;
    END
END MDFFHQX8TR

MACRO MDFFHQX4TR
    CLASS CORE ;
    FOREIGN MDFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.350 2.370 1.630 ;
        RECT  1.680 1.240 1.960 1.630 ;
        END
        ANTENNAGATEAREA 0.5616 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.630 1.810 14.720 2.570 ;
        RECT  14.350 0.440 14.630 3.160 ;
        END
        ANTENNADIFFAREA 3.978 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.440 0.560 1.670 ;
        RECT  0.080 0.840 0.330 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.240 3.920 1.650 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.150 1.230 5.660 1.560 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.110 -0.280 15.200 0.280 ;
        RECT  14.830 -0.280 15.110 1.250 ;
        RECT  14.150 -0.280 14.830 0.280 ;
        RECT  13.870 -0.280 14.150 1.250 ;
        RECT  9.890 -0.280 13.870 0.340 ;
        RECT  9.610 -0.280 9.890 0.400 ;
        RECT  8.570 -0.280 9.610 0.340 ;
        RECT  7.130 -0.280 8.570 0.280 ;
        RECT  6.850 -0.280 7.130 0.610 ;
        RECT  5.630 -0.280 6.850 0.280 ;
        RECT  5.350 -0.280 5.630 0.670 ;
        RECT  4.170 -0.280 5.350 0.280 ;
        RECT  3.890 -0.280 4.170 0.360 ;
        RECT  2.750 -0.280 3.890 0.280 ;
        RECT  2.470 -0.280 2.750 0.360 ;
        RECT  1.710 -0.280 2.470 0.340 ;
        RECT  1.430 -0.280 1.710 0.400 ;
        RECT  0.370 -0.280 1.430 0.280 ;
        RECT  0.090 -0.280 0.370 0.680 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.110 3.320 15.200 3.880 ;
        RECT  14.880 2.080 15.110 3.880 ;
        RECT  14.110 3.320 14.880 3.880 ;
        RECT  13.370 3.200 14.110 3.880 ;
        RECT  10.930 3.260 13.370 3.880 ;
        RECT  10.650 3.200 10.930 3.880 ;
        RECT  9.890 3.320 10.650 3.880 ;
        RECT  9.610 3.200 9.890 3.880 ;
        RECT  8.780 3.260 9.610 3.880 ;
        RECT  8.500 3.200 8.780 3.880 ;
        RECT  7.090 3.320 8.500 3.880 ;
        RECT  6.810 3.200 7.090 3.880 ;
        RECT  6.050 3.320 6.810 3.880 ;
        RECT  5.770 3.200 6.050 3.880 ;
        RECT  4.210 3.320 5.770 3.880 ;
        RECT  3.930 3.200 4.210 3.880 ;
        RECT  2.750 3.320 3.930 3.880 ;
        RECT  2.470 3.200 2.750 3.880 ;
        RECT  1.710 3.260 2.470 3.880 ;
        RECT  1.430 3.200 1.710 3.880 ;
        RECT  0.370 3.320 1.430 3.880 ;
        RECT  0.090 2.430 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.710 2.350 13.810 2.630 ;
        RECT  13.550 0.800 13.710 2.630 ;
        RECT  13.410 0.800 13.550 1.080 ;
        RECT  13.410 1.680 13.550 1.960 ;
        RECT  13.530 2.350 13.550 2.630 ;
        RECT  13.250 1.240 13.390 1.520 ;
        RECT  13.090 0.660 13.250 2.620 ;
        RECT  12.230 0.660 13.090 0.820 ;
        RECT  12.150 2.400 13.090 2.620 ;
        RECT  12.770 0.980 12.930 2.240 ;
        RECT  11.750 0.980 12.770 1.140 ;
        RECT  11.950 2.080 12.770 2.240 ;
        RECT  12.360 2.820 12.640 3.100 ;
        RECT  12.390 1.360 12.610 1.920 ;
        RECT  10.530 1.360 12.390 1.520 ;
        RECT  8.460 2.820 12.360 2.980 ;
        RECT  11.950 0.540 12.230 0.820 ;
        RECT  11.470 2.400 12.150 2.560 ;
        RECT  11.270 0.540 11.950 0.700 ;
        RECT  11.670 1.850 11.950 2.240 ;
        RECT  11.470 0.860 11.750 1.140 ;
        RECT  10.410 1.850 11.670 2.010 ;
        RECT  10.850 0.980 11.470 1.140 ;
        RECT  11.190 2.220 11.470 2.560 ;
        RECT  11.050 0.540 11.270 0.820 ;
        RECT  10.690 0.680 10.850 1.140 ;
        RECT  10.410 0.680 10.690 0.840 ;
        RECT  10.370 1.000 10.530 1.520 ;
        RECT  10.130 0.590 10.410 0.840 ;
        RECT  10.130 1.850 10.410 2.660 ;
        RECT  9.570 1.000 10.370 1.160 ;
        RECT  9.930 1.320 10.210 1.600 ;
        RECT  9.720 2.350 10.130 2.510 ;
        RECT  9.250 1.440 9.930 1.600 ;
        RECT  9.440 2.350 9.720 2.630 ;
        RECT  9.410 0.710 9.570 1.160 ;
        RECT  9.130 0.590 9.410 0.870 ;
        RECT  9.090 1.030 9.250 2.190 ;
        RECT  7.530 0.710 9.130 0.870 ;
        RECT  7.690 1.030 9.090 1.250 ;
        RECT  7.660 1.910 9.090 2.190 ;
        RECT  8.650 1.470 8.930 1.750 ;
        RECT  7.500 1.590 8.650 1.750 ;
        RECT  8.300 2.500 8.460 2.980 ;
        RECT  7.500 2.500 8.300 2.700 ;
        RECT  3.210 2.860 8.140 3.040 ;
        RECT  7.350 0.710 7.530 0.930 ;
        RECT  7.340 1.180 7.500 2.700 ;
        RECT  6.690 0.770 7.350 0.930 ;
        RECT  7.050 1.180 7.340 1.340 ;
        RECT  4.560 2.540 7.340 2.700 ;
        RECT  6.690 1.520 7.180 1.800 ;
        RECT  6.570 0.770 6.690 2.220 ;
        RECT  6.530 0.530 6.570 2.280 ;
        RECT  6.290 0.530 6.530 1.250 ;
        RECT  6.290 2.060 6.530 2.280 ;
        RECT  6.130 1.620 6.370 1.900 ;
        RECT  5.320 2.060 6.290 2.220 ;
        RECT  6.090 0.650 6.130 1.900 ;
        RECT  5.970 0.650 6.090 1.880 ;
        RECT  5.830 0.650 5.970 0.930 ;
        RECT  4.880 1.720 5.970 1.880 ;
        RECT  5.040 2.060 5.320 2.300 ;
        RECT  5.030 0.590 5.150 0.870 ;
        RECT  4.870 0.590 5.030 1.070 ;
        RECT  4.720 1.720 4.880 2.000 ;
        RECT  4.560 0.910 4.870 1.070 ;
        RECT  4.410 0.470 4.690 0.750 ;
        RECT  4.400 0.910 4.560 2.700 ;
        RECT  4.240 0.590 4.410 0.750 ;
        RECT  4.080 0.590 4.240 2.090 ;
        RECT  3.650 0.590 4.080 0.750 ;
        RECT  3.690 1.930 4.080 2.090 ;
        RECT  3.410 1.930 3.690 2.660 ;
        RECT  3.430 0.470 3.650 0.750 ;
        RECT  3.210 0.820 3.240 2.040 ;
        RECT  3.080 0.820 3.210 3.040 ;
        RECT  2.850 0.820 3.080 1.100 ;
        RECT  2.930 1.930 3.080 3.040 ;
        RECT  1.370 2.440 2.930 2.600 ;
        RECT  2.690 1.260 2.920 1.540 ;
        RECT  2.530 0.920 2.690 1.950 ;
        RECT  2.280 0.920 2.530 1.080 ;
        RECT  2.230 1.790 2.530 1.950 ;
        RECT  1.950 0.800 2.280 1.080 ;
        RECT  1.950 1.790 2.230 2.280 ;
        RECT  1.520 1.790 1.950 1.950 ;
        RECT  1.360 1.670 1.520 1.950 ;
        RECT  1.200 1.000 1.370 1.280 ;
        RECT  1.200 2.320 1.370 2.600 ;
        RECT  1.040 1.000 1.200 2.600 ;
        RECT  0.720 0.440 0.880 3.160 ;
        RECT  0.610 0.440 0.720 1.280 ;
        RECT  0.610 1.940 0.720 3.160 ;
    END
END MDFFHQX4TR

MACRO MDFFHQX2TR
    CLASS CORE ;
    FOREIGN MDFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.490 1.550 2.360 ;
        RECT  0.650 0.500 1.390 0.660 ;
        RECT  1.280 2.040 1.390 2.360 ;
        RECT  0.490 0.440 0.650 0.660 ;
        RECT  0.370 0.440 0.490 0.600 ;
        END
        ANTENNAGATEAREA 0.3144 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.680 0.770 9.920 2.610 ;
        RECT  9.360 0.770 9.680 0.930 ;
        RECT  9.370 2.450 9.680 2.610 ;
        RECT  9.210 2.450 9.370 3.000 ;
        RECT  9.200 0.440 9.360 0.930 ;
        END
        ANTENNADIFFAREA 2.636 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.220 0.910 1.560 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.180 3.150 1.660 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.070 1.240 4.350 1.570 ;
        RECT  3.710 1.410 4.070 1.570 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.900 -0.280 10.000 0.280 ;
        RECT  9.620 -0.280 9.900 0.610 ;
        RECT  8.900 -0.280 9.620 0.280 ;
        RECT  8.620 -0.280 8.900 0.300 ;
        RECT  6.900 -0.280 8.620 0.280 ;
        RECT  6.620 -0.280 6.900 0.300 ;
        RECT  5.250 -0.280 6.620 0.280 ;
        RECT  4.970 -0.280 5.250 0.300 ;
        RECT  3.490 -0.280 4.970 0.280 ;
        RECT  3.180 -0.280 3.490 0.640 ;
        RECT  1.330 -0.280 3.180 0.280 ;
        RECT  1.090 -0.280 1.330 0.340 ;
        RECT  0.000 -0.280 1.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.890 3.320 10.000 3.880 ;
        RECT  9.630 2.840 9.890 3.880 ;
        RECT  8.770 3.320 9.630 3.880 ;
        RECT  8.490 2.470 8.770 3.880 ;
        RECT  6.900 3.320 8.490 3.880 ;
        RECT  6.620 3.240 6.900 3.880 ;
        RECT  5.330 3.320 6.620 3.880 ;
        RECT  5.050 3.260 5.330 3.880 ;
        RECT  3.330 3.320 5.050 3.880 ;
        RECT  3.050 3.260 3.330 3.880 ;
        RECT  1.410 3.320 3.050 3.880 ;
        RECT  1.130 3.260 1.410 3.880 ;
        RECT  0.000 3.320 1.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.320 1.090 9.480 2.130 ;
        RECT  9.180 1.090 9.320 1.250 ;
        RECT  8.640 1.970 9.320 2.130 ;
        RECT  9.020 1.480 9.160 1.780 ;
        RECT  8.860 0.500 9.020 1.780 ;
        RECT  8.000 0.500 8.860 0.660 ;
        RECT  8.480 1.400 8.640 2.130 ;
        RECT  8.160 1.070 8.320 3.160 ;
        RECT  7.220 3.000 8.160 3.160 ;
        RECT  7.840 0.500 8.000 2.000 ;
        RECT  7.680 1.840 7.840 2.820 ;
        RECT  7.520 0.520 7.680 1.540 ;
        RECT  5.110 0.520 7.520 0.680 ;
        RECT  7.200 0.840 7.360 2.430 ;
        RECT  7.060 2.590 7.220 3.160 ;
        RECT  6.450 2.270 7.200 2.430 ;
        RECT  6.210 2.590 7.060 2.750 ;
        RECT  6.650 1.170 7.040 1.450 ;
        RECT  6.490 0.960 6.650 2.090 ;
        RECT  6.070 0.960 6.490 1.120 ;
        RECT  6.030 1.930 6.490 2.090 ;
        RECT  5.710 1.610 6.330 1.770 ;
        RECT  6.050 2.560 6.210 2.750 ;
        RECT  5.910 0.840 6.070 1.120 ;
        RECT  5.710 2.560 6.050 2.720 ;
        RECT  5.870 1.930 6.030 2.210 ;
        RECT  5.610 2.910 5.890 3.150 ;
        RECT  5.550 1.230 5.710 2.720 ;
        RECT  2.400 2.910 5.610 3.070 ;
        RECT  5.430 1.230 5.550 1.390 ;
        RECT  3.550 2.560 5.550 2.720 ;
        RECT  5.270 1.110 5.430 1.390 ;
        RECT  5.110 1.550 5.390 1.830 ;
        RECT  4.950 0.520 5.110 2.320 ;
        RECT  4.450 0.520 4.950 0.760 ;
        RECT  4.030 2.160 4.950 2.320 ;
        RECT  4.670 1.170 4.790 1.330 ;
        RECT  4.510 0.920 4.670 1.980 ;
        RECT  4.290 0.920 4.510 1.080 ;
        RECT  3.870 1.820 4.510 1.980 ;
        RECT  4.130 0.450 4.290 1.080 ;
        RECT  3.670 0.450 4.130 0.610 ;
        RECT  3.730 0.850 3.930 1.130 ;
        RECT  3.710 1.770 3.870 2.100 ;
        RECT  3.550 0.970 3.730 1.130 ;
        RECT  3.390 0.970 3.550 2.720 ;
        RECT  2.720 0.810 2.960 0.980 ;
        RECT  2.720 1.970 2.930 2.590 ;
        RECT  2.640 0.810 2.720 2.590 ;
        RECT  2.560 0.810 2.640 2.130 ;
        RECT  2.330 0.880 2.400 3.070 ;
        RECT  2.230 0.760 2.330 3.070 ;
        RECT  2.170 0.760 2.230 1.040 ;
        RECT  0.310 2.910 2.230 3.070 ;
        RECT  1.870 1.200 2.070 1.480 ;
        RECT  1.710 0.560 1.870 2.750 ;
        RECT  0.630 2.590 1.710 2.750 ;
        RECT  1.100 0.900 1.230 1.880 ;
        RECT  1.070 0.900 1.100 2.420 ;
        RECT  0.570 0.900 1.070 1.060 ;
        RECT  0.940 1.720 1.070 2.420 ;
        RECT  0.790 2.090 0.940 2.420 ;
        RECT  0.630 1.720 0.760 1.880 ;
        RECT  0.470 1.720 0.630 2.750 ;
        RECT  0.150 0.930 0.310 3.070 ;
    END
END MDFFHQX2TR

MACRO MDFFHQX1TR
    CLASS CORE ;
    FOREIGN MDFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.500 1.920 1.960 ;
        RECT  1.580 0.810 1.740 1.960 ;
        RECT  1.490 0.810 1.580 0.980 ;
        RECT  1.330 0.520 1.490 0.980 ;
        RECT  0.410 0.520 1.330 0.680 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.680 0.630 9.920 2.530 ;
        RECT  9.520 0.630 9.680 0.790 ;
        RECT  9.440 2.370 9.680 2.530 ;
        RECT  9.360 0.510 9.520 0.790 ;
        RECT  9.280 2.370 9.440 3.160 ;
        END
        ANTENNADIFFAREA 2.104 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.720 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.240 3.520 1.700 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.240 4.470 1.620 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.970 -0.280 10.000 0.280 ;
        RECT  8.690 -0.280 8.970 0.340 ;
        RECT  7.050 -0.280 8.690 0.280 ;
        RECT  6.770 -0.280 7.050 0.340 ;
        RECT  5.410 -0.280 6.770 0.280 ;
        RECT  5.130 -0.280 5.410 0.340 ;
        RECT  3.470 -0.280 5.130 0.280 ;
        RECT  3.190 -0.280 3.470 0.340 ;
        RECT  1.410 -0.280 3.190 0.280 ;
        RECT  1.130 -0.280 1.410 0.340 ;
        RECT  0.000 -0.280 1.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.020 3.320 10.000 3.880 ;
        RECT  8.740 2.480 9.020 3.880 ;
        RECT  7.100 3.320 8.740 3.880 ;
        RECT  6.820 3.260 7.100 3.880 ;
        RECT  5.510 3.320 6.820 3.880 ;
        RECT  5.230 3.260 5.510 3.880 ;
        RECT  3.610 3.320 5.230 3.880 ;
        RECT  3.330 3.260 3.610 3.880 ;
        RECT  1.450 3.320 3.330 3.880 ;
        RECT  1.170 3.260 1.450 3.880 ;
        RECT  0.000 3.320 1.170 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.320 1.030 9.480 2.200 ;
        RECT  8.710 1.970 9.320 2.130 ;
        RECT  8.950 0.620 9.110 1.710 ;
        RECT  8.040 0.620 8.950 0.780 ;
        RECT  8.550 1.580 8.710 2.130 ;
        RECT  8.230 0.940 8.390 3.070 ;
        RECT  6.370 2.910 8.230 3.070 ;
        RECT  7.880 0.620 8.040 2.610 ;
        RECT  7.830 0.900 7.880 1.180 ;
        RECT  7.500 0.440 7.660 0.740 ;
        RECT  7.500 1.050 7.660 2.600 ;
        RECT  5.270 0.580 7.500 0.740 ;
        RECT  7.290 1.050 7.500 1.210 ;
        RECT  7.400 2.320 7.500 2.600 ;
        RECT  6.610 2.440 7.400 2.600 ;
        RECT  6.810 1.470 7.340 1.630 ;
        RECT  6.650 1.020 6.810 2.280 ;
        RECT  6.230 1.020 6.650 1.180 ;
        RECT  5.970 2.120 6.650 2.280 ;
        RECT  5.910 1.660 6.490 1.820 ;
        RECT  6.210 2.620 6.370 3.070 ;
        RECT  6.070 0.900 6.230 1.180 ;
        RECT  5.810 2.620 6.210 2.780 ;
        RECT  2.610 2.940 6.050 3.100 ;
        RECT  5.810 1.140 5.910 1.960 ;
        RECT  5.750 1.140 5.810 2.780 ;
        RECT  5.590 1.140 5.750 1.300 ;
        RECT  5.650 1.800 5.750 2.780 ;
        RECT  3.890 2.620 5.650 2.780 ;
        RECT  5.430 1.020 5.590 1.300 ;
        RECT  5.270 1.480 5.590 1.640 ;
        RECT  5.110 0.580 5.270 2.380 ;
        RECT  4.610 0.580 5.110 0.760 ;
        RECT  4.050 2.220 5.110 2.380 ;
        RECT  4.730 0.920 4.890 1.980 ;
        RECT  4.380 0.920 4.730 1.080 ;
        RECT  4.050 1.820 4.730 1.980 ;
        RECT  4.220 0.450 4.380 1.080 ;
        RECT  3.750 0.450 4.220 0.610 ;
        RECT  3.890 0.920 4.030 1.080 ;
        RECT  3.730 0.920 3.890 2.780 ;
        RECT  2.970 2.080 3.130 2.360 ;
        RECT  2.810 0.700 2.970 2.360 ;
        RECT  2.450 0.640 2.610 3.100 ;
        RECT  2.420 0.640 2.450 0.800 ;
        RECT  0.290 2.940 2.450 3.100 ;
        RECT  2.260 0.520 2.420 0.800 ;
        RECT  2.130 0.960 2.290 2.300 ;
        RECT  2.100 0.960 2.130 1.120 ;
        RECT  1.950 2.120 2.130 2.300 ;
        RECT  1.940 0.490 2.100 1.120 ;
        RECT  1.710 2.120 1.950 2.510 ;
        RECT  1.650 0.490 1.940 0.650 ;
        RECT  0.730 2.350 1.710 2.510 ;
        RECT  0.720 1.970 0.930 2.130 ;
        RECT  0.720 0.900 0.890 1.060 ;
        RECT  0.450 2.350 0.730 2.590 ;
        RECT  0.560 0.900 0.720 2.130 ;
        RECT  0.350 1.910 0.390 2.190 ;
        RECT  0.290 0.840 0.350 2.190 ;
        RECT  0.130 0.840 0.290 3.100 ;
    END
END MDFFHQX1TR

MACRO INVXLTR
    CLASS CORE ;
    FOREIGN INVXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.440 1.120 2.250 ;
        RECT  0.780 0.440 0.880 1.230 ;
        RECT  0.680 1.930 0.880 2.250 ;
        END
        ANTENNADIFFAREA 1.086 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.390 0.680 1.670 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 -0.280 1.200 0.280 ;
        RECT  0.160 -0.280 0.440 1.080 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 3.320 1.200 3.880 ;
        RECT  0.160 2.520 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
END INVXLTR

MACRO INVX8TR
    CLASS CORE ;
    FOREIGN INVX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.040 2.120 1.810 ;
        RECT  1.850 0.600 1.890 1.810 ;
        RECT  1.530 0.600 1.850 2.890 ;
        RECT  1.480 0.600 1.530 2.280 ;
        RECT  0.570 0.600 1.480 1.080 ;
        RECT  0.850 1.800 1.480 2.280 ;
        RECT  0.570 1.800 0.850 3.160 ;
        END
        ANTENNADIFFAREA 7.676 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 1.160 1.640 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 1.0056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 -0.280 2.800 0.280 ;
        RECT  2.090 -0.280 2.370 0.870 ;
        RECT  1.370 -0.280 2.090 0.340 ;
        RECT  1.090 -0.280 1.370 0.400 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 3.320 2.800 3.880 ;
        RECT  2.010 1.970 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.590 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.240 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END INVX8TR

MACRO INVX6TR
    CLASS CORE ;
    FOREIGN INVX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.040 2.120 1.760 ;
        RECT  1.910 0.590 2.000 1.760 ;
        RECT  1.700 0.590 1.910 3.020 ;
        RECT  1.620 1.040 1.700 3.020 ;
        RECT  1.480 1.040 1.620 2.480 ;
        RECT  0.940 1.040 1.480 1.400 ;
        RECT  0.940 2.120 1.480 2.480 ;
        RECT  0.660 0.540 0.940 1.400 ;
        RECT  0.660 2.120 0.940 3.060 ;
        END
        ANTENNADIFFAREA 7.62 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.640 1.280 1.800 ;
        RECT  0.460 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.7584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.280 2.400 0.280 ;
        RECT  1.140 -0.280 1.460 0.780 ;
        RECT  0.460 -0.280 1.140 0.280 ;
        RECT  0.180 -0.280 0.460 1.200 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 3.320 2.400 3.880 ;
        RECT  1.970 3.240 2.250 3.880 ;
        RECT  1.420 3.320 1.970 3.880 ;
        RECT  1.140 2.770 1.420 3.880 ;
        RECT  0.460 3.320 1.140 3.880 ;
        RECT  0.180 2.340 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
END INVX6TR

MACRO INVX4TR
    CLASS CORE ;
    FOREIGN INVX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.070 1.120 2.170 ;
        RECT  0.850 1.070 0.880 1.310 ;
        RECT  0.850 1.910 0.880 2.170 ;
        RECT  0.570 0.520 0.850 1.310 ;
        RECT  0.570 1.910 0.850 3.080 ;
        END
        ANTENNADIFFAREA 3.762 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.470 0.650 1.750 ;
        RECT  0.320 1.470 0.360 2.360 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.4848 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.280 1.600 0.280 ;
        RECT  1.050 -0.280 1.330 0.860 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.420 3.320 1.600 3.880 ;
        RECT  1.140 2.420 1.420 3.880 ;
        RECT  0.370 3.320 1.140 3.880 ;
        RECT  0.090 2.530 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END INVX4TR

MACRO INVX3TR
    CLASS CORE ;
    FOREIGN INVX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.630 1.120 1.990 ;
        RECT  0.930 0.800 1.050 1.990 ;
        RECT  0.880 0.800 0.930 2.750 ;
        RECT  0.650 0.800 0.880 1.080 ;
        RECT  0.650 1.830 0.880 2.750 ;
        END
        ANTENNADIFFAREA 2.898 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.240 0.720 1.580 ;
        END
        ANTENNAGATEAREA 0.3864 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.280 1.600 0.280 ;
        RECT  1.210 -0.280 1.460 1.080 ;
        RECT  0.470 -0.280 1.210 0.280 ;
        RECT  0.190 -0.280 0.470 1.080 ;
        RECT  0.000 -0.280 0.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 1.600 3.880 ;
        RECT  1.110 2.220 1.400 3.880 ;
        RECT  0.460 3.260 1.110 3.880 ;
        RECT  0.190 2.200 0.460 3.880 ;
        RECT  0.000 3.320 0.190 3.880 ;
        END
    END VDD
END INVX3TR

MACRO INVX2TR
    CLASS CORE ;
    FOREIGN INVX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.240 1.120 2.360 ;
        RECT  0.960 0.440 1.000 2.360 ;
        RECT  0.840 0.440 0.960 3.160 ;
        RECT  0.680 0.440 0.840 1.310 ;
        RECT  0.680 1.910 0.840 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.470 0.680 1.750 ;
        RECT  0.360 1.240 0.400 1.750 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 -0.280 1.200 0.280 ;
        RECT  0.160 -0.280 0.440 0.990 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 3.320 1.200 3.880 ;
        RECT  0.160 2.750 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
END INVX2TR

MACRO INVX20TR
    CLASS CORE ;
    FOREIGN INVX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 0.650 4.700 2.830 ;
        RECT  3.740 0.840 4.420 2.130 ;
        RECT  3.460 0.440 3.740 3.160 ;
        RECT  3.280 0.840 3.460 2.130 ;
        RECT  2.780 0.920 3.280 2.130 ;
        RECT  2.500 0.440 2.780 3.160 ;
        RECT  1.820 0.920 2.500 2.130 ;
        RECT  1.540 0.440 1.820 3.160 ;
        RECT  0.860 0.920 1.540 2.130 ;
        RECT  0.580 0.920 0.860 2.890 ;
        END
        ANTENNADIFFAREA 19.255 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.420 2.360 ;
        END
        ANTENNAGATEAREA 2.5416 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.180 -0.280 5.600 0.280 ;
        RECT  4.900 -0.280 5.180 1.310 ;
        RECT  4.220 -0.280 4.900 0.280 ;
        RECT  3.940 -0.280 4.220 0.670 ;
        RECT  3.260 -0.280 3.940 0.280 ;
        RECT  2.980 -0.280 3.260 0.670 ;
        RECT  2.300 -0.280 2.980 0.280 ;
        RECT  2.020 -0.280 2.300 0.670 ;
        RECT  1.340 -0.280 2.020 0.280 ;
        RECT  1.060 -0.280 1.340 0.670 ;
        RECT  0.380 -0.280 1.060 0.340 ;
        RECT  0.100 -0.280 0.380 1.020 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.200 3.320 5.600 3.880 ;
        RECT  4.900 2.020 5.200 3.880 ;
        RECT  4.220 3.320 4.900 3.880 ;
        RECT  3.940 2.490 4.220 3.880 ;
        RECT  3.260 3.320 3.940 3.880 ;
        RECT  2.980 2.480 3.260 3.880 ;
        RECT  2.300 3.320 2.980 3.880 ;
        RECT  2.020 2.490 2.300 3.880 ;
        RECT  1.340 3.320 2.020 3.880 ;
        RECT  1.060 2.480 1.340 3.880 ;
        RECT  0.380 3.260 1.060 3.880 ;
        RECT  0.100 2.520 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
END INVX20TR

MACRO INVX1TR
    CLASS CORE ;
    FOREIGN INVX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.440 1.120 2.430 ;
        RECT  0.870 0.440 0.880 1.230 ;
        RECT  0.680 2.120 0.880 2.430 ;
        RECT  0.680 0.840 0.870 1.230 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.640 0.720 1.960 ;
        RECT  0.400 1.390 0.680 1.960 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 -0.280 1.200 0.280 ;
        RECT  0.200 -0.280 0.480 1.220 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 3.320 1.200 3.880 ;
        RECT  0.200 2.190 0.480 3.880 ;
        RECT  0.000 3.320 0.200 3.880 ;
        END
    END VDD
END INVX1TR

MACRO INVX16TR
    CLASS CORE ;
    FOREIGN INVX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.040 0.840 4.320 1.960 ;
        RECT  3.760 0.440 4.040 3.160 ;
        RECT  3.280 0.840 3.760 1.970 ;
        RECT  3.080 0.990 3.280 1.970 ;
        RECT  2.800 0.440 3.080 3.160 ;
        RECT  2.120 1.000 2.800 1.960 ;
        RECT  1.840 0.440 2.120 3.160 ;
        RECT  1.160 1.000 1.840 1.960 ;
        RECT  0.880 0.650 1.160 3.080 ;
        END
        ANTENNADIFFAREA 15.608 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.240 0.720 1.640 ;
        RECT  0.160 1.390 0.430 1.640 ;
        END
        ANTENNAGATEAREA 2.076 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.280 4.800 0.280 ;
        RECT  4.240 -0.280 4.520 0.680 ;
        RECT  3.560 -0.280 4.240 0.280 ;
        RECT  3.280 -0.280 3.560 0.670 ;
        RECT  2.600 -0.280 3.280 0.280 ;
        RECT  2.320 -0.280 2.600 0.670 ;
        RECT  1.640 -0.280 2.320 0.280 ;
        RECT  1.360 -0.280 1.640 0.670 ;
        RECT  0.680 -0.280 1.360 0.340 ;
        RECT  0.400 -0.280 0.680 1.080 ;
        RECT  0.000 -0.280 0.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 3.320 4.800 3.880 ;
        RECT  4.240 2.310 4.520 3.880 ;
        RECT  3.560 3.320 4.240 3.880 ;
        RECT  3.280 2.490 3.560 3.880 ;
        RECT  2.600 3.320 3.280 3.880 ;
        RECT  2.320 2.440 2.600 3.880 ;
        RECT  1.640 3.320 2.320 3.880 ;
        RECT  1.360 2.480 1.640 3.880 ;
        RECT  0.680 3.320 1.360 3.880 ;
        RECT  0.400 1.910 0.680 3.880 ;
        RECT  0.000 3.320 0.400 3.880 ;
        END
    END VDD
END INVX16TR

MACRO INVX12TR
    CLASS CORE ;
    FOREIGN INVX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 0.440 2.790 3.160 ;
        RECT  1.830 1.040 2.510 1.760 ;
        RECT  1.550 0.440 1.830 3.160 ;
        RECT  0.870 1.040 1.550 1.760 ;
        RECT  0.590 0.650 0.870 2.890 ;
        END
        ANTENNADIFFAREA 11.572 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.430 1.680 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 1.536 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.280 3.600 0.280 ;
        RECT  2.990 -0.280 3.270 1.310 ;
        RECT  2.310 -0.280 2.990 0.280 ;
        RECT  2.030 -0.280 2.310 0.670 ;
        RECT  1.350 -0.280 2.030 0.280 ;
        RECT  1.070 -0.280 1.350 0.670 ;
        RECT  0.390 -0.280 1.070 0.340 ;
        RECT  0.110 -0.280 0.390 1.030 ;
        RECT  0.000 -0.280 0.110 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 3.320 3.600 3.880 ;
        RECT  2.990 1.910 3.270 3.880 ;
        RECT  2.310 3.320 2.990 3.880 ;
        RECT  2.030 2.130 2.310 3.880 ;
        RECT  1.350 3.320 2.030 3.880 ;
        RECT  1.070 2.120 1.350 3.880 ;
        RECT  0.390 3.260 1.070 3.880 ;
        RECT  0.110 2.610 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
END INVX12TR

MACRO HOLDX1TR
    CLASS CORE ;
    FOREIGN HOLDX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION INOUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.440 1.520 1.960 ;
        RECT  1.240 0.440 1.490 2.190 ;
        RECT  1.210 1.800 1.240 2.190 ;
        RECT  0.690 1.800 1.210 1.960 ;
        RECT  0.530 1.470 0.690 1.960 ;
        RECT  0.400 1.470 0.530 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.840 -0.280 1.600 0.280 ;
        RECT  0.560 -0.280 0.840 0.800 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 3.320 1.600 3.880 ;
        RECT  0.650 2.120 0.930 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 1.150 1.020 1.640 ;
        RECT  0.370 1.150 0.860 1.310 ;
        RECT  0.240 0.520 0.370 1.310 ;
        RECT  0.240 1.910 0.370 2.190 ;
        RECT  0.080 0.520 0.240 2.190 ;
    END
END HOLDX1TR

MACRO FILL8TR
    CLASS CORE SPACER ;
    FOREIGN FILL8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 3.200 3.880 ;
        END
    END VDD
END FILL8TR

MACRO FILL64TR
    CLASS CORE SPACER ;
    FOREIGN FILL64TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 25.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 25.600 3.880 ;
        END
    END VDD
END FILL64TR

MACRO FILL4TR
    CLASS CORE SPACER ;
    FOREIGN FILL4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 1.600 3.880 ;
        END
    END VDD
END FILL4TR

MACRO FILL32TR
    CLASS CORE SPACER ;
    FOREIGN FILL32TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 12.800 3.880 ;
        END
    END VDD
END FILL32TR

MACRO FILL2TR
    CLASS CORE SPACER ;
    FOREIGN FILL2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
END FILL2TR

MACRO FILL16TR
    CLASS CORE SPACER ;
    FOREIGN FILL16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 6.400 3.880 ;
        END
    END VDD
END FILL16TR

MACRO FILL1TR
    CLASS CORE SPACER ;
    FOREIGN FILL1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 0.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 0.400 3.880 ;
        END
    END VDD
END FILL1TR

MACRO EDFFTRXLTR
    CLASS CORE ;
    FOREIGN EDFFTRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.440 1.530 0.870 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.320 1.240 9.520 1.560 ;
        RECT  9.280 1.240 9.320 2.380 ;
        RECT  9.160 0.770 9.280 2.380 ;
        RECT  9.120 0.770 9.160 1.410 ;
        RECT  9.020 2.220 9.160 2.380 ;
        END
        ANTENNADIFFAREA 1.0745 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.250 1.640 10.320 2.760 ;
        RECT  10.080 0.480 10.250 2.760 ;
        END
        ANTENNADIFFAREA 1.7195 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.080 3.300 1.240 ;
        RECT  2.650 1.080 2.810 1.960 ;
        RECT  1.920 1.800 2.650 1.960 ;
        RECT  1.680 1.640 1.920 1.960 ;
        RECT  1.120 1.640 1.680 1.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.640 3.560 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.340 -0.280 10.400 0.280 ;
        RECT  8.180 -0.280 8.340 0.400 ;
        RECT  6.750 -0.280 8.180 0.280 ;
        RECT  6.450 -0.280 6.750 0.950 ;
        RECT  5.320 -0.280 6.450 0.280 ;
        RECT  5.160 -0.280 5.320 0.470 ;
        RECT  2.710 -0.280 5.160 0.280 ;
        RECT  2.430 -0.280 2.710 0.300 ;
        RECT  0.900 -0.280 2.430 0.280 ;
        RECT  0.620 -0.280 0.900 0.740 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.780 3.320 10.400 3.880 ;
        RECT  9.480 2.860 9.780 3.880 ;
        RECT  8.380 3.320 9.480 3.880 ;
        RECT  8.220 3.200 8.380 3.880 ;
        RECT  6.690 3.320 8.220 3.880 ;
        RECT  6.410 3.260 6.690 3.880 ;
        RECT  5.260 3.320 6.410 3.880 ;
        RECT  4.980 3.260 5.260 3.880 ;
        RECT  2.760 3.320 4.980 3.880 ;
        RECT  2.480 3.260 2.760 3.880 ;
        RECT  1.540 3.320 2.480 3.880 ;
        RECT  0.840 2.680 1.540 3.880 ;
        RECT  0.000 3.320 0.840 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.840 1.360 9.920 1.640 ;
        RECT  9.680 0.450 9.840 2.700 ;
        RECT  8.560 0.450 9.680 0.610 ;
        RECT  9.240 2.540 9.680 2.700 ;
        RECT  9.080 2.540 9.240 3.160 ;
        RECT  8.930 1.820 9.000 1.980 ;
        RECT  8.780 1.200 8.930 1.980 ;
        RECT  8.770 1.200 8.780 2.400 ;
        RECT  8.620 1.820 8.770 2.400 ;
        RECT  8.200 2.240 8.620 2.400 ;
        RECT  8.370 1.230 8.530 1.550 ;
        RECT  7.650 1.230 8.370 1.390 ;
        RECT  8.080 1.850 8.200 2.400 ;
        RECT  7.920 1.850 8.080 2.990 ;
        RECT  2.330 2.830 7.920 2.990 ;
        RECT  7.200 0.450 7.870 0.610 ;
        RECT  7.490 0.860 7.650 2.330 ;
        RECT  7.360 0.860 7.490 1.110 ;
        RECT  7.470 2.170 7.490 2.330 ;
        RECT  7.310 2.170 7.470 2.450 ;
        RECT  7.200 1.850 7.330 2.010 ;
        RECT  7.040 0.450 7.200 2.010 ;
        RECT  6.620 1.850 7.040 2.010 ;
        RECT  6.500 1.190 6.620 2.010 ;
        RECT  6.340 1.190 6.500 2.670 ;
        RECT  4.040 2.510 6.340 2.670 ;
        RECT  6.000 0.610 6.180 2.350 ;
        RECT  5.800 0.610 6.000 0.870 ;
        RECT  5.820 1.530 5.840 1.810 ;
        RECT  5.660 1.030 5.820 2.240 ;
        RECT  5.510 0.440 5.800 0.870 ;
        RECT  5.600 1.030 5.660 1.590 ;
        RECT  5.500 2.080 5.660 2.240 ;
        RECT  5.000 1.430 5.600 1.590 ;
        RECT  4.820 0.710 5.510 0.870 ;
        RECT  5.320 1.750 5.500 1.910 ;
        RECT  5.160 1.750 5.320 2.030 ;
        RECT  4.360 1.870 5.160 2.030 ;
        RECT  4.840 1.430 5.000 1.710 ;
        RECT  4.660 0.710 4.820 1.270 ;
        RECT  4.520 0.990 4.660 1.270 ;
        RECT  4.360 0.670 4.500 0.830 ;
        RECT  4.200 0.670 4.360 2.350 ;
        RECT  3.880 1.080 4.040 2.670 ;
        RECT  3.720 0.640 3.880 0.920 ;
        RECT  1.620 2.120 3.880 2.280 ;
        RECT  1.850 0.760 3.720 0.920 ;
        RECT  1.940 2.440 3.720 2.600 ;
        RECT  2.330 1.320 2.490 1.620 ;
        RECT  1.280 1.320 2.330 1.480 ;
        RECT  2.170 2.830 2.330 3.110 ;
        RECT  1.780 2.440 1.940 2.930 ;
        RECT  1.690 0.760 1.850 1.160 ;
        RECT  1.460 2.120 1.620 2.520 ;
        RECT  0.640 2.360 1.460 2.520 ;
        RECT  0.960 2.040 1.300 2.200 ;
        RECT  1.120 1.030 1.280 1.480 ;
        RECT  0.960 1.320 1.120 1.480 ;
        RECT  0.800 1.320 0.960 2.200 ;
        RECT  0.480 0.900 0.640 2.860 ;
        RECT  0.380 0.900 0.480 1.060 ;
        RECT  0.160 2.640 0.480 2.860 ;
        RECT  0.220 0.460 0.380 1.060 ;
    END
END EDFFTRXLTR

MACRO EDFFTRX4TR
    CLASS CORE ;
    FOREIGN EDFFTRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.440 1.560 0.800 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.080 1.090 10.380 2.250 ;
        END
        ANTENNADIFFAREA 4.07 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.200 0.580 11.440 3.160 ;
        RECT  11.060 0.580 11.200 1.240 ;
        RECT  11.060 1.840 11.200 3.160 ;
        RECT  10.880 1.840 11.060 2.560 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.100 3.340 1.270 ;
        RECT  2.690 1.100 2.850 1.980 ;
        RECT  1.920 1.820 2.690 1.980 ;
        RECT  1.670 1.640 1.920 1.980 ;
        RECT  1.150 1.640 1.670 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.640 3.600 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.820 -0.280 12.000 0.280 ;
        RECT  11.600 -0.280 11.820 1.320 ;
        RECT  10.880 -0.280 11.600 0.280 ;
        RECT  10.570 -0.280 10.880 0.610 ;
        RECT  9.890 -0.280 10.570 0.280 ;
        RECT  9.610 -0.280 9.890 0.610 ;
        RECT  8.400 -0.280 9.610 0.280 ;
        RECT  8.120 -0.280 8.400 0.400 ;
        RECT  6.830 -0.280 8.120 0.280 ;
        RECT  6.550 -0.280 6.830 0.990 ;
        RECT  5.420 -0.280 6.550 0.280 ;
        RECT  5.140 -0.280 5.420 0.340 ;
        RECT  2.750 -0.280 5.140 0.280 ;
        RECT  2.470 -0.280 2.750 0.340 ;
        RECT  0.900 -0.280 2.470 0.280 ;
        RECT  0.620 -0.280 0.900 0.740 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.870 3.320 12.000 3.880 ;
        RECT  11.600 2.080 11.870 3.880 ;
        RECT  10.870 3.320 11.600 3.880 ;
        RECT  10.560 2.790 10.870 3.880 ;
        RECT  9.890 3.320 10.560 3.880 ;
        RECT  9.610 2.900 9.890 3.880 ;
        RECT  8.420 3.320 9.610 3.880 ;
        RECT  8.190 2.120 8.420 3.880 ;
        RECT  1.580 3.320 8.190 3.880 ;
        RECT  0.840 2.860 1.580 3.880 ;
        RECT  0.000 3.320 0.840 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.700 1.420 11.010 1.640 ;
        RECT  10.540 0.770 10.700 2.630 ;
        RECT  9.400 0.770 10.540 0.930 ;
        RECT  9.360 2.470 10.540 2.630 ;
        RECT  9.410 1.090 9.600 1.900 ;
        RECT  8.860 1.090 9.410 1.250 ;
        RECT  8.900 1.740 9.410 1.900 ;
        RECT  9.100 0.450 9.400 0.930 ;
        RECT  9.090 2.220 9.360 2.630 ;
        RECT  8.620 1.740 8.900 3.150 ;
        RECT  8.700 0.600 8.860 1.250 ;
        RECT  8.500 1.420 8.710 1.580 ;
        RECT  8.180 1.740 8.620 1.900 ;
        RECT  8.340 0.930 8.500 1.580 ;
        RECT  7.660 0.930 8.340 1.090 ;
        RECT  8.030 1.570 8.180 1.900 ;
        RECT  7.870 1.570 8.030 3.160 ;
        RECT  7.200 0.440 7.880 0.600 ;
        RECT  2.430 3.000 7.870 3.160 ;
        RECT  7.540 0.810 7.660 2.350 ;
        RECT  7.500 0.810 7.540 2.810 ;
        RECT  7.360 0.810 7.500 1.370 ;
        RECT  7.260 2.190 7.500 2.810 ;
        RECT  7.200 1.870 7.340 2.030 ;
        RECT  7.040 0.440 7.200 2.030 ;
        RECT  6.600 1.870 7.040 2.030 ;
        RECT  6.540 1.210 6.600 2.030 ;
        RECT  6.360 1.210 6.540 2.810 ;
        RECT  4.020 2.650 6.360 2.810 ;
        RECT  6.200 0.630 6.280 0.820 ;
        RECT  6.040 0.630 6.200 2.440 ;
        RECT  5.880 0.630 6.040 0.830 ;
        RECT  5.610 0.440 5.880 0.830 ;
        RECT  5.840 1.550 5.880 1.880 ;
        RECT  5.680 1.030 5.840 2.310 ;
        RECT  5.660 1.030 5.680 1.560 ;
        RECT  5.520 2.150 5.680 2.310 ;
        RECT  4.980 1.400 5.660 1.560 ;
        RECT  4.860 0.670 5.610 0.830 ;
        RECT  5.330 1.720 5.520 1.890 ;
        RECT  5.140 1.720 5.330 2.000 ;
        RECT  4.400 1.840 5.140 2.000 ;
        RECT  4.820 1.400 4.980 1.680 ;
        RECT  4.700 0.670 4.860 1.240 ;
        RECT  4.560 0.960 4.700 1.240 ;
        RECT  4.400 0.640 4.540 0.800 ;
        RECT  4.240 0.640 4.400 2.370 ;
        RECT  4.180 2.090 4.240 2.370 ;
        RECT  4.020 1.100 4.080 1.380 ;
        RECT  3.860 1.100 4.020 2.810 ;
        RECT  3.760 0.660 3.920 0.940 ;
        RECT  1.650 2.140 3.860 2.300 ;
        RECT  1.890 0.780 3.760 0.940 ;
        RECT  1.970 2.460 3.700 2.620 ;
        RECT  2.370 1.310 2.530 1.640 ;
        RECT  2.180 2.910 2.430 3.160 ;
        RECT  1.280 1.310 2.370 1.470 ;
        RECT  1.810 2.460 1.970 3.080 ;
        RECT  1.730 0.780 1.890 1.150 ;
        RECT  1.490 2.140 1.650 2.700 ;
        RECT  0.640 2.540 1.490 2.700 ;
        RECT  1.030 2.120 1.310 2.350 ;
        RECT  1.120 1.030 1.280 1.470 ;
        RECT  0.990 1.310 1.120 1.470 ;
        RECT  0.990 2.120 1.030 2.280 ;
        RECT  0.830 1.310 0.990 2.280 ;
        RECT  0.480 0.920 0.640 2.700 ;
        RECT  0.350 0.920 0.480 1.080 ;
        RECT  0.350 2.540 0.480 2.700 ;
        RECT  0.090 0.840 0.350 1.080 ;
        RECT  0.090 2.540 0.350 3.090 ;
    END
END EDFFTRX4TR

MACRO EDFFTRX2TR
    CLASS CORE ;
    FOREIGN EDFFTRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.440 1.560 0.800 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.990 1.090 10.090 1.300 ;
        RECT  9.680 1.090 9.990 2.250 ;
        END
        ANTENNADIFFAREA 2.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.050 2.030 11.120 3.160 ;
        RECT  10.780 0.580 11.050 3.160 ;
        END
        ANTENNADIFFAREA 3.904 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.100 3.340 1.270 ;
        RECT  2.690 1.100 2.850 1.980 ;
        RECT  1.920 1.820 2.690 1.980 ;
        RECT  1.670 1.640 1.920 1.980 ;
        RECT  1.150 1.640 1.670 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.640 3.600 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.590 -0.280 11.200 0.280 ;
        RECT  10.310 -0.280 10.590 0.480 ;
        RECT  9.190 -0.280 10.310 0.280 ;
        RECT  8.900 -0.280 9.190 0.640 ;
        RECT  8.520 -0.280 8.900 0.280 ;
        RECT  8.240 -0.280 8.520 0.400 ;
        RECT  6.830 -0.280 8.240 0.280 ;
        RECT  6.550 -0.280 6.830 0.990 ;
        RECT  5.420 -0.280 6.550 0.280 ;
        RECT  5.140 -0.280 5.420 0.340 ;
        RECT  2.750 -0.280 5.140 0.280 ;
        RECT  2.470 -0.280 2.750 0.340 ;
        RECT  0.870 -0.280 2.470 0.280 ;
        RECT  0.590 -0.280 0.870 0.740 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.480 3.320 11.200 3.880 ;
        RECT  10.170 2.790 10.480 3.880 ;
        RECT  9.180 3.320 10.170 3.880 ;
        RECT  8.920 2.860 9.180 3.880 ;
        RECT  8.360 3.320 8.920 3.880 ;
        RECT  7.960 3.260 8.360 3.880 ;
        RECT  6.700 3.320 7.960 3.880 ;
        RECT  6.420 3.260 6.700 3.880 ;
        RECT  5.280 3.320 6.420 3.880 ;
        RECT  5.000 3.260 5.280 3.880 ;
        RECT  2.820 3.320 5.000 3.880 ;
        RECT  2.540 3.260 2.820 3.880 ;
        RECT  1.580 3.320 2.540 3.880 ;
        RECT  0.840 2.860 1.580 3.880 ;
        RECT  0.000 3.320 0.840 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.460 0.750 10.620 2.630 ;
        RECT  9.760 0.750 10.460 0.910 ;
        RECT  9.640 2.470 10.460 2.630 ;
        RECT  9.590 0.450 9.760 0.910 ;
        RECT  9.440 2.470 9.640 3.150 ;
        RECT  9.470 0.450 9.590 0.720 ;
        RECT  9.110 1.600 9.440 1.900 ;
        RECT  9.370 2.850 9.440 3.150 ;
        RECT  8.950 1.090 9.110 1.900 ;
        RECT  8.620 1.090 8.950 1.250 ;
        RECT  8.820 1.740 8.950 1.900 ;
        RECT  8.540 1.740 8.820 2.500 ;
        RECT  7.660 1.420 8.710 1.580 ;
        RECT  8.030 1.740 8.540 1.900 ;
        RECT  7.870 1.740 8.030 3.090 ;
        RECT  7.200 0.440 7.880 0.600 ;
        RECT  2.370 2.880 7.870 3.090 ;
        RECT  7.500 0.810 7.660 2.350 ;
        RECT  7.360 0.810 7.500 0.970 ;
        RECT  7.480 2.190 7.500 2.350 ;
        RECT  7.320 2.190 7.480 2.470 ;
        RECT  7.200 1.870 7.340 2.030 ;
        RECT  7.040 0.440 7.200 2.030 ;
        RECT  6.600 1.870 7.040 2.030 ;
        RECT  6.540 1.210 6.600 2.030 ;
        RECT  6.360 1.210 6.540 2.690 ;
        RECT  4.020 2.530 6.360 2.690 ;
        RECT  6.200 0.640 6.280 0.830 ;
        RECT  6.040 0.640 6.200 2.370 ;
        RECT  5.880 0.640 6.040 0.830 ;
        RECT  5.610 0.440 5.880 0.830 ;
        RECT  5.840 1.550 5.880 1.880 ;
        RECT  5.680 1.030 5.840 2.210 ;
        RECT  5.660 1.030 5.680 1.560 ;
        RECT  5.520 2.050 5.680 2.210 ;
        RECT  4.980 1.400 5.660 1.560 ;
        RECT  4.860 0.670 5.610 0.830 ;
        RECT  5.330 1.720 5.520 1.890 ;
        RECT  5.140 1.720 5.330 2.000 ;
        RECT  4.400 1.840 5.140 2.000 ;
        RECT  4.820 1.400 4.980 1.680 ;
        RECT  4.700 0.670 4.860 1.240 ;
        RECT  4.560 0.960 4.700 1.240 ;
        RECT  4.400 0.640 4.540 0.800 ;
        RECT  4.240 0.640 4.400 2.370 ;
        RECT  4.180 2.090 4.240 2.370 ;
        RECT  4.020 1.100 4.080 1.380 ;
        RECT  3.860 1.100 4.020 2.690 ;
        RECT  3.760 0.660 3.920 0.940 ;
        RECT  1.650 2.140 3.860 2.300 ;
        RECT  1.890 0.780 3.760 0.940 ;
        RECT  1.970 2.460 3.700 2.620 ;
        RECT  2.370 1.310 2.530 1.640 ;
        RECT  1.250 1.310 2.370 1.470 ;
        RECT  2.180 2.880 2.370 3.160 ;
        RECT  1.810 2.460 1.970 3.080 ;
        RECT  1.730 0.780 1.890 1.150 ;
        RECT  1.490 2.140 1.650 2.700 ;
        RECT  0.640 2.540 1.490 2.700 ;
        RECT  1.030 2.120 1.310 2.350 ;
        RECT  1.090 1.030 1.250 1.470 ;
        RECT  0.990 1.310 1.090 1.470 ;
        RECT  0.990 2.120 1.030 2.280 ;
        RECT  0.830 1.310 0.990 2.280 ;
        RECT  0.480 0.920 0.640 2.700 ;
        RECT  0.350 0.920 0.480 1.080 ;
        RECT  0.350 2.540 0.480 2.700 ;
        RECT  0.190 0.440 0.350 1.080 ;
        RECT  0.190 2.540 0.350 3.130 ;
    END
END EDFFTRX2TR

MACRO EDFFTRX1TR
    CLASS CORE ;
    FOREIGN EDFFTRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.440 1.560 0.800 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.340 1.090 9.520 1.560 ;
        RECT  9.320 0.970 9.340 1.560 ;
        RECT  9.160 0.970 9.320 2.250 ;
        RECT  8.950 2.080 9.160 2.250 ;
        END
        ANTENNADIFFAREA 1.728 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.270 2.030 10.320 3.160 ;
        RECT  10.080 0.820 10.270 3.160 ;
        END
        ANTENNADIFFAREA 1.824 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.100 3.340 1.270 ;
        RECT  2.690 1.100 2.850 1.980 ;
        RECT  1.920 1.820 2.690 1.980 ;
        RECT  1.670 1.640 1.920 1.980 ;
        RECT  1.150 1.640 1.670 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.640 3.600 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.340 -0.280 10.400 0.280 ;
        RECT  8.180 -0.280 8.340 0.400 ;
        RECT  6.830 -0.280 8.180 0.280 ;
        RECT  6.550 -0.280 6.830 0.990 ;
        RECT  5.420 -0.280 6.550 0.280 ;
        RECT  5.140 -0.280 5.420 0.340 ;
        RECT  2.750 -0.280 5.140 0.280 ;
        RECT  2.470 -0.280 2.750 0.340 ;
        RECT  0.870 -0.280 2.470 0.280 ;
        RECT  0.590 -0.280 0.870 0.740 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.750 3.320 10.400 3.880 ;
        RECT  9.470 2.790 9.750 3.880 ;
        RECT  8.360 3.320 9.470 3.880 ;
        RECT  8.200 3.190 8.360 3.880 ;
        RECT  6.700 3.320 8.200 3.880 ;
        RECT  6.420 3.260 6.700 3.880 ;
        RECT  5.280 3.320 6.420 3.880 ;
        RECT  5.000 3.260 5.280 3.880 ;
        RECT  2.820 3.320 5.000 3.880 ;
        RECT  2.540 3.260 2.820 3.880 ;
        RECT  1.580 3.320 2.540 3.880 ;
        RECT  0.840 2.860 1.580 3.880 ;
        RECT  0.000 3.320 0.840 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.840 1.360 9.920 1.640 ;
        RECT  9.680 0.450 9.840 2.630 ;
        RECT  8.990 0.450 9.680 0.610 ;
        RECT  9.270 2.470 9.680 2.630 ;
        RECT  9.020 2.470 9.270 3.150 ;
        RECT  8.800 0.930 8.960 1.920 ;
        RECT  8.640 0.930 8.800 1.090 ;
        RECT  8.760 1.760 8.800 1.920 ;
        RECT  8.600 1.760 8.760 2.500 ;
        RECT  8.440 1.250 8.600 1.530 ;
        RECT  8.190 1.760 8.600 1.930 ;
        RECT  7.660 1.250 8.440 1.410 ;
        RECT  8.030 1.730 8.190 1.930 ;
        RECT  7.870 1.730 8.030 3.090 ;
        RECT  7.200 0.440 7.880 0.600 ;
        RECT  2.370 2.880 7.870 3.090 ;
        RECT  7.500 0.810 7.660 2.350 ;
        RECT  7.360 0.810 7.500 0.970 ;
        RECT  7.480 2.190 7.500 2.350 ;
        RECT  7.320 2.190 7.480 2.470 ;
        RECT  7.200 1.870 7.340 2.030 ;
        RECT  7.040 0.440 7.200 2.030 ;
        RECT  6.600 1.870 7.040 2.030 ;
        RECT  6.540 1.210 6.600 2.030 ;
        RECT  6.360 1.210 6.540 2.690 ;
        RECT  4.020 2.530 6.360 2.690 ;
        RECT  6.200 0.640 6.280 0.830 ;
        RECT  6.040 0.640 6.200 2.370 ;
        RECT  5.880 0.640 6.040 0.830 ;
        RECT  5.610 0.440 5.880 0.830 ;
        RECT  5.840 1.550 5.880 1.880 ;
        RECT  5.680 1.030 5.840 2.210 ;
        RECT  5.660 1.030 5.680 1.560 ;
        RECT  5.520 2.050 5.680 2.210 ;
        RECT  4.980 1.400 5.660 1.560 ;
        RECT  4.860 0.670 5.610 0.830 ;
        RECT  5.330 1.720 5.520 1.890 ;
        RECT  5.140 1.720 5.330 2.000 ;
        RECT  4.400 1.840 5.140 2.000 ;
        RECT  4.820 1.400 4.980 1.680 ;
        RECT  4.700 0.670 4.860 1.240 ;
        RECT  4.560 0.960 4.700 1.240 ;
        RECT  4.400 0.640 4.540 0.800 ;
        RECT  4.240 0.640 4.400 2.370 ;
        RECT  4.180 2.090 4.240 2.370 ;
        RECT  4.020 1.100 4.080 1.380 ;
        RECT  3.860 1.100 4.020 2.690 ;
        RECT  3.760 0.660 3.920 0.940 ;
        RECT  1.650 2.140 3.860 2.300 ;
        RECT  1.890 0.780 3.760 0.940 ;
        RECT  1.970 2.460 3.700 2.620 ;
        RECT  2.370 1.310 2.530 1.640 ;
        RECT  1.250 1.310 2.370 1.470 ;
        RECT  2.180 2.880 2.370 3.160 ;
        RECT  1.810 2.460 1.970 3.080 ;
        RECT  1.730 0.780 1.890 1.150 ;
        RECT  1.490 2.140 1.650 2.700 ;
        RECT  0.640 2.540 1.490 2.700 ;
        RECT  1.030 2.120 1.310 2.350 ;
        RECT  1.090 1.030 1.250 1.470 ;
        RECT  0.990 1.310 1.090 1.470 ;
        RECT  0.990 2.120 1.030 2.280 ;
        RECT  0.830 1.310 0.990 2.280 ;
        RECT  0.480 0.920 0.640 2.700 ;
        RECT  0.350 0.920 0.480 1.080 ;
        RECT  0.350 2.540 0.480 2.700 ;
        RECT  0.190 0.460 0.350 1.080 ;
        RECT  0.190 2.540 0.350 2.930 ;
    END
END EDFFTRX1TR

MACRO EDFFHQX8TR
    CLASS CORE ;
    FOREIGN EDFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.910 0.450 15.190 3.150 ;
        RECT  14.230 1.440 14.910 2.160 ;
        RECT  13.950 0.440 14.230 3.160 ;
        RECT  13.880 1.440 13.950 2.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.2424 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.310 0.680 1.620 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.280 5.260 1.560 ;
        RECT  4.760 1.240 5.120 1.560 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.670 -0.280 16.000 0.280 ;
        RECT  15.390 -0.280 15.670 1.220 ;
        RECT  14.710 -0.280 15.390 0.280 ;
        RECT  14.430 -0.280 14.710 1.220 ;
        RECT  13.690 -0.280 14.430 0.280 ;
        RECT  13.530 -0.280 13.690 1.220 ;
        RECT  12.820 -0.280 13.530 0.340 ;
        RECT  12.540 -0.280 12.820 0.380 ;
        RECT  5.780 -0.280 12.540 0.280 ;
        RECT  5.500 -0.280 5.780 0.360 ;
        RECT  5.020 -0.280 5.500 0.280 ;
        RECT  4.740 -0.280 5.020 0.360 ;
        RECT  3.800 -0.280 4.740 0.280 ;
        RECT  3.520 -0.280 3.800 0.400 ;
        RECT  1.940 -0.280 3.520 0.280 ;
        RECT  1.630 -0.280 1.940 0.910 ;
        RECT  0.480 -0.280 1.630 0.280 ;
        RECT  0.200 -0.280 0.480 0.670 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.670 3.320 16.000 3.880 ;
        RECT  15.390 2.040 15.670 3.880 ;
        RECT  14.710 3.320 15.390 3.880 ;
        RECT  14.430 2.510 14.710 3.880 ;
        RECT  13.750 3.320 14.430 3.880 ;
        RECT  13.470 2.990 13.750 3.880 ;
        RECT  12.890 3.320 13.470 3.880 ;
        RECT  12.610 2.850 12.890 3.880 ;
        RECT  10.480 3.260 12.610 3.880 ;
        RECT  10.200 3.200 10.480 3.880 ;
        RECT  9.440 3.320 10.200 3.880 ;
        RECT  9.160 3.200 9.440 3.880 ;
        RECT  8.310 3.260 9.160 3.880 ;
        RECT  8.030 3.200 8.310 3.880 ;
        RECT  6.620 3.320 8.030 3.880 ;
        RECT  6.340 3.200 6.620 3.880 ;
        RECT  5.580 3.320 6.340 3.880 ;
        RECT  5.300 3.200 5.580 3.880 ;
        RECT  3.740 3.320 5.300 3.880 ;
        RECT  3.460 3.200 3.740 3.880 ;
        RECT  1.960 3.260 3.460 3.880 ;
        RECT  1.630 2.860 1.960 3.880 ;
        RECT  0.480 3.320 1.630 3.880 ;
        RECT  0.200 2.190 0.480 3.880 ;
        RECT  0.000 3.320 0.200 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.370 2.320 13.410 2.640 ;
        RECT  13.210 0.540 13.370 2.640 ;
        RECT  13.070 0.540 13.210 1.050 ;
        RECT  13.190 1.930 13.210 2.640 ;
        RECT  12.380 0.540 13.070 0.700 ;
        RECT  12.910 1.210 12.990 1.490 ;
        RECT  12.750 0.860 12.910 2.600 ;
        RECT  11.860 0.860 12.750 1.020 ;
        RECT  10.990 2.440 12.750 2.600 ;
        RECT  12.430 1.240 12.590 2.260 ;
        RECT  11.340 1.240 12.430 1.400 ;
        RECT  11.470 2.100 12.430 2.260 ;
        RECT  12.220 0.440 12.380 0.700 ;
        RECT  12.080 1.560 12.240 1.940 ;
        RECT  6.100 0.440 12.220 0.600 ;
        RECT  10.640 2.820 12.160 3.100 ;
        RECT  10.080 1.560 12.080 1.720 ;
        RECT  11.580 0.760 11.860 1.020 ;
        RECT  10.760 0.760 11.580 0.920 ;
        RECT  11.190 1.940 11.470 2.260 ;
        RECT  11.060 1.080 11.340 1.400 ;
        RECT  9.960 1.940 11.190 2.100 ;
        RECT  10.400 1.240 11.060 1.400 ;
        RECT  10.710 2.260 10.990 2.600 ;
        RECT  10.600 0.760 10.760 1.040 ;
        RECT  7.990 2.820 10.640 2.980 ;
        RECT  10.240 0.760 10.400 1.400 ;
        RECT  9.680 0.760 10.240 0.920 ;
        RECT  9.920 1.080 10.080 1.720 ;
        RECT  9.680 1.940 9.960 2.660 ;
        RECT  9.230 1.080 9.920 1.240 ;
        RECT  9.480 1.440 9.760 1.660 ;
        RECT  8.990 2.350 9.680 2.510 ;
        RECT  8.720 1.500 9.480 1.660 ;
        RECT  9.070 0.760 9.230 1.240 ;
        RECT  6.420 0.760 9.070 0.920 ;
        RECT  8.560 1.080 8.720 2.240 ;
        RECT  8.400 1.080 8.560 1.300 ;
        RECT  7.190 1.960 8.560 2.240 ;
        RECT  7.220 1.080 8.400 1.240 ;
        RECT  7.030 1.570 8.400 1.730 ;
        RECT  7.830 2.500 7.990 2.980 ;
        RECT  7.030 2.500 7.830 2.660 ;
        RECT  6.940 2.940 7.670 3.100 ;
        RECT  6.870 1.110 7.030 2.660 ;
        RECT  6.780 2.880 6.940 3.100 ;
        RECT  6.580 1.110 6.870 1.390 ;
        RECT  3.280 2.500 6.870 2.660 ;
        RECT  2.960 2.880 6.780 3.040 ;
        RECT  6.420 1.550 6.710 1.830 ;
        RECT  6.260 0.760 6.420 2.220 ;
        RECT  5.820 1.000 6.260 1.280 ;
        RECT  6.100 2.060 6.260 2.220 ;
        RECT  5.940 0.440 6.100 0.680 ;
        RECT  5.820 2.060 6.100 2.280 ;
        RECT  4.820 0.520 5.940 0.680 ;
        RECT  5.620 1.620 5.900 1.900 ;
        RECT  4.700 2.060 5.820 2.220 ;
        RECT  5.580 1.620 5.620 1.880 ;
        RECT  5.420 0.840 5.580 1.880 ;
        RECT  5.320 0.840 5.420 1.120 ;
        RECT  4.260 1.720 5.420 1.880 ;
        RECT  4.660 0.520 4.820 1.080 ;
        RECT  4.420 2.060 4.700 2.280 ;
        RECT  3.660 0.920 4.660 1.080 ;
        RECT  4.220 0.480 4.500 0.760 ;
        RECT  3.980 1.600 4.260 1.880 ;
        RECT  3.280 0.600 4.220 0.760 ;
        RECT  3.440 0.920 3.660 1.250 ;
        RECT  3.120 0.600 3.280 2.660 ;
        RECT  2.800 0.500 2.960 3.040 ;
        RECT  2.680 0.500 2.800 0.720 ;
        RECT  1.440 2.490 2.800 2.650 ;
        RECT  2.500 0.920 2.640 2.330 ;
        RECT  2.480 0.630 2.500 2.330 ;
        RECT  2.220 0.630 2.480 1.080 ;
        RECT  1.880 2.050 2.480 2.330 ;
        RECT  1.600 1.720 1.880 2.330 ;
        RECT  1.320 0.580 1.440 1.290 ;
        RECT  1.320 2.040 1.440 3.160 ;
        RECT  1.160 0.580 1.320 3.160 ;
        RECT  0.840 0.440 1.000 3.160 ;
        RECT  0.680 0.440 0.840 1.080 ;
        RECT  0.680 1.950 0.840 3.160 ;
    END
END EDFFHQX8TR

MACRO EDFFHQX4TR
    CLASS CORE ;
    FOREIGN EDFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.950 0.440 14.230 3.160 ;
        RECT  13.680 1.840 13.950 2.560 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.240 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.2424 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.310 0.680 1.620 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.280 5.260 1.560 ;
        RECT  4.760 1.240 5.120 1.560 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.710 -0.280 14.800 0.280 ;
        RECT  14.430 -0.280 14.710 1.220 ;
        RECT  13.770 -0.280 14.430 0.280 ;
        RECT  13.530 -0.280 13.770 1.220 ;
        RECT  12.820 -0.280 13.530 0.340 ;
        RECT  12.540 -0.280 12.820 0.380 ;
        RECT  5.020 -0.280 12.540 0.280 ;
        RECT  4.740 -0.280 5.020 0.360 ;
        RECT  3.800 -0.280 4.740 0.280 ;
        RECT  3.520 -0.280 3.800 0.400 ;
        RECT  1.940 -0.280 3.520 0.280 ;
        RECT  1.660 -0.280 1.940 0.860 ;
        RECT  0.480 -0.280 1.660 0.280 ;
        RECT  0.200 -0.280 0.480 0.670 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.710 3.320 14.800 3.880 ;
        RECT  14.430 1.820 14.710 3.880 ;
        RECT  13.750 3.320 14.430 3.880 ;
        RECT  13.470 2.870 13.750 3.880 ;
        RECT  12.940 3.320 13.470 3.880 ;
        RECT  12.610 2.760 12.940 3.880 ;
        RECT  10.480 3.260 12.610 3.880 ;
        RECT  10.200 3.200 10.480 3.880 ;
        RECT  9.440 3.320 10.200 3.880 ;
        RECT  9.160 3.200 9.440 3.880 ;
        RECT  8.310 3.260 9.160 3.880 ;
        RECT  8.030 3.200 8.310 3.880 ;
        RECT  6.620 3.320 8.030 3.880 ;
        RECT  6.340 3.200 6.620 3.880 ;
        RECT  5.580 3.320 6.340 3.880 ;
        RECT  5.300 3.200 5.580 3.880 ;
        RECT  3.740 3.320 5.300 3.880 ;
        RECT  3.460 3.200 3.740 3.880 ;
        RECT  1.960 3.260 3.460 3.880 ;
        RECT  1.620 2.860 1.960 3.880 ;
        RECT  0.480 3.320 1.620 3.880 ;
        RECT  0.200 2.190 0.480 3.880 ;
        RECT  0.000 3.320 0.200 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.150 0.540 13.310 3.000 ;
        RECT  13.060 0.540 13.150 1.050 ;
        RECT  13.120 1.680 13.150 3.000 ;
        RECT  12.370 0.540 13.060 0.700 ;
        RECT  12.880 1.210 12.990 1.490 ;
        RECT  12.720 0.860 12.880 2.600 ;
        RECT  11.860 0.860 12.720 1.020 ;
        RECT  10.990 2.440 12.720 2.600 ;
        RECT  12.400 1.240 12.560 2.260 ;
        RECT  11.340 1.240 12.400 1.400 ;
        RECT  11.470 2.100 12.400 2.260 ;
        RECT  12.210 0.440 12.370 0.700 ;
        RECT  12.080 1.560 12.240 1.940 ;
        RECT  6.090 0.440 12.210 0.600 ;
        RECT  10.640 2.820 12.160 3.100 ;
        RECT  10.080 1.560 12.080 1.720 ;
        RECT  11.580 0.760 11.860 1.020 ;
        RECT  10.760 0.760 11.580 0.920 ;
        RECT  11.190 1.940 11.470 2.260 ;
        RECT  11.060 1.080 11.340 1.400 ;
        RECT  9.960 1.940 11.190 2.100 ;
        RECT  10.400 1.240 11.060 1.400 ;
        RECT  10.710 2.260 10.990 2.600 ;
        RECT  10.600 0.760 10.760 1.040 ;
        RECT  7.990 2.820 10.640 2.980 ;
        RECT  10.240 0.760 10.400 1.400 ;
        RECT  9.680 0.760 10.240 0.920 ;
        RECT  9.920 1.080 10.080 1.720 ;
        RECT  9.680 1.940 9.960 2.660 ;
        RECT  9.230 1.080 9.920 1.240 ;
        RECT  9.480 1.440 9.760 1.660 ;
        RECT  8.990 2.350 9.680 2.510 ;
        RECT  8.720 1.500 9.480 1.660 ;
        RECT  9.070 0.760 9.230 1.240 ;
        RECT  6.420 0.760 9.070 0.920 ;
        RECT  8.560 1.080 8.720 2.240 ;
        RECT  8.400 1.080 8.560 1.300 ;
        RECT  7.190 1.960 8.560 2.240 ;
        RECT  7.220 1.080 8.400 1.240 ;
        RECT  7.030 1.570 8.400 1.730 ;
        RECT  7.830 2.500 7.990 2.980 ;
        RECT  7.030 2.500 7.830 2.660 ;
        RECT  6.940 2.940 7.670 3.100 ;
        RECT  6.870 1.230 7.030 2.660 ;
        RECT  6.780 2.880 6.940 3.100 ;
        RECT  6.860 1.230 6.870 1.390 ;
        RECT  3.280 2.500 6.870 2.660 ;
        RECT  6.580 1.110 6.860 1.390 ;
        RECT  2.960 2.880 6.780 3.040 ;
        RECT  6.420 1.550 6.710 1.830 ;
        RECT  6.260 0.760 6.420 2.220 ;
        RECT  5.820 1.000 6.260 1.280 ;
        RECT  6.100 2.060 6.260 2.220 ;
        RECT  5.820 2.060 6.100 2.280 ;
        RECT  5.930 0.440 6.090 0.680 ;
        RECT  4.920 0.520 5.930 0.680 ;
        RECT  5.620 1.620 5.900 1.900 ;
        RECT  4.700 2.060 5.820 2.220 ;
        RECT  5.580 1.620 5.620 1.880 ;
        RECT  5.420 0.840 5.580 1.880 ;
        RECT  5.320 0.840 5.420 1.120 ;
        RECT  4.260 1.720 5.420 1.880 ;
        RECT  4.760 0.520 4.920 1.080 ;
        RECT  3.650 0.920 4.760 1.080 ;
        RECT  4.420 2.060 4.700 2.280 ;
        RECT  4.220 0.480 4.500 0.760 ;
        RECT  3.980 1.600 4.260 1.880 ;
        RECT  3.280 0.600 4.220 0.760 ;
        RECT  3.440 0.920 3.650 1.250 ;
        RECT  3.120 0.600 3.280 2.660 ;
        RECT  2.800 0.500 2.960 3.040 ;
        RECT  2.680 0.500 2.800 0.720 ;
        RECT  1.440 2.490 2.800 2.650 ;
        RECT  2.500 0.920 2.640 2.330 ;
        RECT  2.480 0.630 2.500 2.330 ;
        RECT  2.220 0.630 2.480 1.080 ;
        RECT  1.880 2.050 2.480 2.330 ;
        RECT  1.600 1.720 1.880 2.330 ;
        RECT  1.320 0.520 1.440 1.290 ;
        RECT  1.320 2.040 1.440 3.160 ;
        RECT  1.160 0.520 1.320 3.160 ;
        RECT  0.840 0.440 1.000 3.160 ;
        RECT  0.680 0.440 0.840 1.080 ;
        RECT  0.680 1.950 0.840 3.160 ;
    END
END EDFFHQX4TR

MACRO EDFFHQX2TR
    CLASS CORE ;
    FOREIGN EDFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 0.440 10.720 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.450 1.640 1.960 ;
        RECT  1.280 0.540 1.440 1.960 ;
        RECT  0.680 0.540 1.280 0.700 ;
        RECT  0.520 0.470 0.680 0.700 ;
        RECT  0.370 0.470 0.520 0.630 ;
        END
        ANTENNAGATEAREA 0.1512 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.800 1.960 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.040 3.820 1.630 ;
        RECT  3.440 1.470 3.600 1.960 ;
        RECT  3.280 1.640 3.440 1.960 ;
        END
        ANTENNAGATEAREA 0.216 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.230 -0.280 10.800 0.280 ;
        RECT  9.950 -0.280 10.230 0.760 ;
        RECT  9.090 -0.280 9.950 0.300 ;
        RECT  3.240 -0.280 9.090 0.280 ;
        RECT  2.960 -0.280 3.240 0.400 ;
        RECT  1.370 -0.280 2.960 0.280 ;
        RECT  1.090 -0.280 1.370 0.380 ;
        RECT  0.000 -0.280 1.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.230 3.320 10.800 3.880 ;
        RECT  8.900 2.800 10.230 3.880 ;
        RECT  7.300 3.320 8.900 3.880 ;
        RECT  7.020 3.260 7.300 3.880 ;
        RECT  5.440 3.320 7.020 3.880 ;
        RECT  5.160 3.200 5.440 3.880 ;
        RECT  3.500 3.320 5.160 3.880 ;
        RECT  3.220 3.200 3.500 3.880 ;
        RECT  1.640 3.260 3.220 3.880 ;
        RECT  1.360 3.200 1.640 3.880 ;
        RECT  0.000 3.320 1.360 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.070 1.040 10.230 2.050 ;
        RECT  9.640 1.040 10.070 1.200 ;
        RECT  9.640 1.890 10.070 2.050 ;
        RECT  9.630 1.360 9.910 1.640 ;
        RECT  9.360 0.920 9.640 1.200 ;
        RECT  9.360 1.890 9.640 2.210 ;
        RECT  8.830 1.360 9.630 1.520 ;
        RECT  9.150 0.920 9.360 1.080 ;
        RECT  9.210 1.890 9.360 2.050 ;
        RECT  8.990 1.770 9.210 2.050 ;
        RECT  8.990 0.460 9.150 1.080 ;
        RECT  8.340 0.460 8.990 0.620 ;
        RECT  8.670 0.780 8.830 2.460 ;
        RECT  8.180 0.780 8.670 1.000 ;
        RECT  8.020 2.300 8.670 2.460 ;
        RECT  8.230 1.190 8.510 2.130 ;
        RECT  8.230 2.940 8.510 3.160 ;
        RECT  8.180 0.440 8.340 0.620 ;
        RECT  8.020 1.190 8.230 1.410 ;
        RECT  6.750 2.940 8.230 3.100 ;
        RECT  3.680 0.440 8.180 0.600 ;
        RECT  7.860 0.760 8.020 1.410 ;
        RECT  5.240 0.760 7.860 0.920 ;
        RECT  7.700 1.800 7.820 2.720 ;
        RECT  7.540 1.080 7.700 2.720 ;
        RECT  7.400 1.080 7.540 1.240 ;
        RECT  6.910 2.360 7.540 2.640 ;
        RECT  6.960 1.560 7.380 1.720 ;
        RECT  6.800 1.140 6.960 2.190 ;
        RECT  6.120 1.140 6.800 1.320 ;
        RECT  6.120 2.030 6.800 2.190 ;
        RECT  6.590 2.560 6.750 3.100 ;
        RECT  5.960 1.680 6.640 1.840 ;
        RECT  5.960 2.560 6.590 2.720 ;
        RECT  6.210 2.880 6.430 3.160 ;
        RECT  2.520 2.880 6.210 3.040 ;
        RECT  5.800 1.300 5.960 2.720 ;
        RECT  5.680 1.300 5.800 1.460 ;
        RECT  2.840 2.560 5.800 2.720 ;
        RECT  5.400 1.180 5.680 1.460 ;
        RECT  5.240 1.620 5.640 1.900 ;
        RECT  5.080 0.760 5.240 2.280 ;
        RECT  4.610 0.760 5.080 1.060 ;
        RECT  4.300 2.000 5.080 2.280 ;
        RECT  4.140 1.330 4.920 1.610 ;
        RECT  4.140 0.770 4.320 0.990 ;
        RECT  3.980 0.770 4.140 1.970 ;
        RECT  3.760 1.810 3.980 1.970 ;
        RECT  3.520 0.440 3.680 0.720 ;
        RECT  3.440 0.560 3.520 0.720 ;
        RECT  3.280 0.560 3.440 1.310 ;
        RECT  3.000 1.150 3.280 1.430 ;
        RECT  2.900 0.710 3.120 0.990 ;
        RECT  2.840 0.830 2.900 0.990 ;
        RECT  2.680 0.830 2.840 2.720 ;
        RECT  2.360 0.550 2.520 3.040 ;
        RECT  1.680 0.550 2.360 0.830 ;
        RECT  2.240 2.520 2.360 3.040 ;
        RECT  0.420 2.880 2.240 3.040 ;
        RECT  2.080 1.350 2.200 1.630 ;
        RECT  2.080 2.020 2.200 2.300 ;
        RECT  1.920 1.010 2.080 2.720 ;
        RECT  1.600 1.010 1.920 1.290 ;
        RECT  0.680 2.560 1.920 2.720 ;
        RECT  0.960 0.860 1.120 2.400 ;
        RECT  0.570 0.860 0.960 1.080 ;
        RECT  0.840 2.120 0.960 2.400 ;
        RECT  0.520 2.170 0.680 2.720 ;
        RECT  0.400 2.170 0.520 2.450 ;
        RECT  0.360 2.880 0.420 3.140 ;
        RECT  0.240 0.790 0.370 1.070 ;
        RECT  0.240 2.610 0.360 3.140 ;
        RECT  0.080 0.790 0.240 3.140 ;
    END
END EDFFHQX2TR

MACRO EDFFHQX1TR
    CLASS CORE ;
    FOREIGN EDFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 0.440 10.720 2.950 ;
        END
        ANTENNADIFFAREA 1.92 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.450 1.640 1.960 ;
        RECT  1.280 0.540 1.440 1.960 ;
        RECT  0.680 0.540 1.280 0.700 ;
        RECT  0.520 0.470 0.680 0.700 ;
        RECT  0.370 0.470 0.520 0.630 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.800 1.960 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.040 3.820 1.630 ;
        RECT  3.440 1.470 3.600 1.960 ;
        RECT  3.280 1.640 3.440 1.960 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.230 -0.280 10.800 0.280 ;
        RECT  9.420 -0.280 10.230 0.760 ;
        RECT  1.370 -0.280 9.420 0.280 ;
        RECT  1.090 -0.280 1.370 0.380 ;
        RECT  0.000 -0.280 1.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.230 3.320 10.800 3.880 ;
        RECT  8.900 2.640 10.230 3.880 ;
        RECT  7.300 3.320 8.900 3.880 ;
        RECT  7.020 3.260 7.300 3.880 ;
        RECT  5.440 3.320 7.020 3.880 ;
        RECT  5.160 3.200 5.440 3.880 ;
        RECT  3.500 3.320 5.160 3.880 ;
        RECT  3.220 3.200 3.500 3.880 ;
        RECT  1.640 3.260 3.220 3.880 ;
        RECT  1.360 3.200 1.640 3.880 ;
        RECT  0.000 3.320 1.360 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.070 1.040 10.230 2.050 ;
        RECT  9.640 1.040 10.070 1.200 ;
        RECT  9.640 1.890 10.070 2.050 ;
        RECT  9.630 1.360 9.910 1.640 ;
        RECT  9.360 0.920 9.640 1.200 ;
        RECT  9.360 1.890 9.640 2.210 ;
        RECT  8.830 1.360 9.630 1.520 ;
        RECT  9.150 0.920 9.360 1.080 ;
        RECT  9.210 1.890 9.360 2.050 ;
        RECT  8.990 1.770 9.210 2.050 ;
        RECT  8.990 0.460 9.150 1.080 ;
        RECT  8.340 0.460 8.990 0.620 ;
        RECT  8.670 0.780 8.830 2.460 ;
        RECT  8.180 0.780 8.670 1.000 ;
        RECT  8.020 2.300 8.670 2.460 ;
        RECT  8.230 1.190 8.510 2.130 ;
        RECT  8.230 2.940 8.510 3.160 ;
        RECT  8.180 0.440 8.340 0.620 ;
        RECT  8.020 1.190 8.230 1.410 ;
        RECT  6.750 2.940 8.230 3.100 ;
        RECT  3.680 0.440 8.180 0.600 ;
        RECT  7.860 0.760 8.020 1.410 ;
        RECT  5.240 0.760 7.860 0.920 ;
        RECT  7.700 1.800 7.820 2.720 ;
        RECT  7.540 1.080 7.700 2.720 ;
        RECT  7.400 1.080 7.540 1.240 ;
        RECT  6.910 2.360 7.540 2.640 ;
        RECT  6.960 1.560 7.380 1.720 ;
        RECT  6.800 1.140 6.960 2.190 ;
        RECT  6.120 1.140 6.800 1.320 ;
        RECT  6.120 2.030 6.800 2.190 ;
        RECT  6.590 2.560 6.750 3.100 ;
        RECT  5.960 1.680 6.640 1.840 ;
        RECT  5.960 2.560 6.590 2.720 ;
        RECT  5.820 2.880 6.040 3.160 ;
        RECT  5.800 1.300 5.960 2.720 ;
        RECT  2.520 2.880 5.820 3.040 ;
        RECT  5.680 1.300 5.800 1.460 ;
        RECT  2.840 2.560 5.800 2.720 ;
        RECT  5.400 1.180 5.680 1.460 ;
        RECT  5.240 1.620 5.640 1.900 ;
        RECT  5.080 0.760 5.240 2.280 ;
        RECT  4.610 0.760 5.080 1.070 ;
        RECT  4.300 2.000 5.080 2.280 ;
        RECT  4.140 1.330 4.920 1.610 ;
        RECT  4.140 0.770 4.320 0.990 ;
        RECT  3.980 0.770 4.140 1.970 ;
        RECT  3.760 1.810 3.980 1.970 ;
        RECT  3.520 0.440 3.680 0.720 ;
        RECT  3.440 0.560 3.520 0.720 ;
        RECT  3.280 0.560 3.440 1.310 ;
        RECT  3.000 1.150 3.280 1.430 ;
        RECT  2.900 0.710 3.120 0.990 ;
        RECT  2.840 0.830 2.900 0.990 ;
        RECT  2.680 0.830 2.840 2.720 ;
        RECT  2.360 0.550 2.520 3.040 ;
        RECT  1.680 0.550 2.360 0.830 ;
        RECT  2.240 2.520 2.360 3.040 ;
        RECT  0.360 2.880 2.240 3.040 ;
        RECT  2.080 1.350 2.200 1.630 ;
        RECT  2.080 2.020 2.200 2.300 ;
        RECT  1.920 1.010 2.080 2.720 ;
        RECT  1.600 1.010 1.920 1.290 ;
        RECT  0.680 2.560 1.920 2.720 ;
        RECT  0.960 0.860 1.120 2.400 ;
        RECT  0.570 0.860 0.960 1.080 ;
        RECT  0.840 2.180 0.960 2.400 ;
        RECT  0.520 2.170 0.680 2.720 ;
        RECT  0.400 2.170 0.520 2.390 ;
        RECT  0.240 0.800 0.370 1.080 ;
        RECT  0.240 2.600 0.360 3.040 ;
        RECT  0.080 0.800 0.240 3.040 ;
    END
END EDFFHQX1TR

MACRO EDFFXLTR
    CLASS CORE ;
    FOREIGN EDFFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.030 9.520 2.760 ;
        RECT  9.230 1.030 9.280 1.310 ;
        RECT  9.200 2.280 9.280 2.760 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.910 0.680 9.070 2.010 ;
        RECT  8.480 0.680 8.910 0.840 ;
        RECT  8.880 1.850 8.910 2.010 ;
        RECT  8.720 1.850 8.880 2.820 ;
        RECT  8.160 2.440 8.720 2.820 ;
        RECT  8.200 0.560 8.480 0.840 ;
        END
        ANTENNADIFFAREA 1.046 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.330 2.770 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.840 2.250 2.120 ;
        RECT  1.970 1.590 2.130 2.120 ;
        RECT  1.960 1.590 1.970 1.750 ;
        RECT  1.800 1.240 1.960 1.750 ;
        RECT  1.640 1.240 1.800 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.160 1.690 ;
        RECT  4.680 1.530 4.880 1.690 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.940 -0.280 9.600 0.280 ;
        RECT  8.660 -0.280 8.940 0.400 ;
        RECT  7.920 -0.280 8.660 0.280 ;
        RECT  7.640 -0.280 7.920 0.400 ;
        RECT  6.340 -0.280 7.640 0.340 ;
        RECT  6.060 -0.280 6.340 0.660 ;
        RECT  4.820 -0.280 6.060 0.280 ;
        RECT  4.540 -0.280 4.820 0.760 ;
        RECT  3.780 -0.280 4.540 0.280 ;
        RECT  3.500 -0.280 3.780 0.990 ;
        RECT  1.710 -0.280 3.500 0.280 ;
        RECT  1.430 -0.280 1.710 0.400 ;
        RECT  0.370 -0.280 1.430 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.900 3.320 9.600 3.880 ;
        RECT  8.620 3.200 8.900 3.880 ;
        RECT  7.920 3.320 8.620 3.880 ;
        RECT  7.640 2.420 7.920 3.880 ;
        RECT  5.410 3.260 7.640 3.880 ;
        RECT  3.210 3.320 5.410 3.880 ;
        RECT  1.690 3.260 3.210 3.880 ;
        RECT  1.410 3.200 1.690 3.880 ;
        RECT  0.370 3.320 1.410 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.640 1.410 8.750 1.690 ;
        RECT  8.560 1.050 8.640 1.690 ;
        RECT  8.400 1.050 8.560 2.220 ;
        RECT  8.200 1.050 8.400 1.340 ;
        RECT  7.420 1.980 8.400 2.220 ;
        RECT  7.960 1.500 8.240 1.780 ;
        RECT  7.130 1.620 7.960 1.780 ;
        RECT  7.220 1.980 7.420 3.100 ;
        RECT  7.120 0.700 7.400 0.980 ;
        RECT  4.120 2.940 7.220 3.100 ;
        RECT  6.980 1.140 7.130 1.780 ;
        RECT  6.400 0.820 7.120 0.980 ;
        RECT  6.840 1.140 6.980 2.660 ;
        RECT  6.820 1.140 6.840 2.780 ;
        RECT  6.560 2.500 6.820 2.780 ;
        RECT  6.400 2.060 6.620 2.340 ;
        RECT  6.240 0.820 6.400 2.780 ;
        RECT  5.900 0.820 6.240 0.980 ;
        RECT  4.740 2.560 6.240 2.780 ;
        RECT  5.920 1.220 6.080 2.400 ;
        RECT  5.620 1.220 5.920 1.380 ;
        RECT  5.220 2.240 5.920 2.400 ;
        RECT  5.740 0.440 5.900 0.980 ;
        RECT  5.480 1.740 5.760 2.020 ;
        RECT  5.140 0.440 5.740 0.600 ;
        RECT  5.580 1.100 5.620 1.380 ;
        RECT  5.340 0.760 5.580 1.380 ;
        RECT  4.460 1.860 5.480 2.020 ;
        RECT  5.300 0.760 5.340 0.980 ;
        RECT  4.940 2.180 5.220 2.400 ;
        RECT  4.980 0.440 5.140 1.080 ;
        RECT  4.720 0.920 4.980 1.080 ;
        RECT  4.460 2.430 4.740 2.780 ;
        RECT  4.500 0.920 4.720 1.370 ;
        RECT  4.340 1.860 4.460 2.250 ;
        RECT  2.710 2.430 4.460 2.650 ;
        RECT  4.180 0.630 4.340 2.250 ;
        RECT  4.060 0.630 4.180 1.310 ;
        RECT  3.960 2.810 4.120 3.100 ;
        RECT  3.650 1.150 4.060 1.310 ;
        RECT  3.800 1.520 4.020 1.800 ;
        RECT  0.770 2.810 3.960 3.030 ;
        RECT  3.090 1.640 3.800 1.800 ;
        RECT  3.370 1.150 3.650 1.430 ;
        RECT  3.030 1.640 3.090 2.270 ;
        RECT  2.870 0.440 3.030 2.270 ;
        RECT  2.620 0.440 2.870 0.720 ;
        RECT  2.550 1.350 2.710 2.650 ;
        RECT  2.410 1.350 2.550 1.630 ;
        RECT  2.170 2.370 2.390 2.650 ;
        RECT  2.090 0.440 2.370 0.850 ;
        RECT  0.810 2.490 2.170 2.650 ;
        RECT  0.830 0.690 2.090 0.850 ;
        RECT  1.450 2.040 1.810 2.320 ;
        RECT  1.290 1.280 1.450 2.320 ;
        RECT  1.170 1.280 1.290 1.560 ;
        RECT  0.810 1.280 1.170 1.440 ;
        RECT  0.550 0.570 0.830 0.850 ;
        RECT  0.650 1.030 0.810 2.190 ;
        RECT  0.530 2.370 0.810 2.650 ;
        RECT  0.530 1.030 0.650 1.360 ;
        RECT  0.530 1.910 0.650 2.190 ;
    END
END EDFFXLTR

MACRO EDFFX4TR
    CLASS CORE ;
    FOREIGN EDFFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.900 1.040 11.920 1.760 ;
        RECT  11.820 1.040 11.900 2.940 ;
        RECT  11.680 0.570 11.820 2.940 ;
        RECT  11.540 0.570 11.680 1.210 ;
        RECT  11.600 1.940 11.680 2.940 ;
        END
        ANTENNADIFFAREA 4.134 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.770 0.530 10.780 1.640 ;
        RECT  10.480 0.530 10.770 2.330 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.160 0.370 2.370 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.630 1.170 1.810 ;
        RECT  0.790 1.630 1.130 1.960 ;
        RECT  0.670 1.640 0.790 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.580 4.440 1.960 ;
        END
        ANTENNAGATEAREA 0.1032 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.270 -0.280 12.400 0.280 ;
        RECT  12.080 -0.280 12.270 1.240 ;
        RECT  11.300 -0.280 12.080 0.280 ;
        RECT  11.020 -0.280 11.300 1.190 ;
        RECT  10.270 -0.280 11.020 0.280 ;
        RECT  9.990 -0.280 10.270 0.480 ;
        RECT  9.370 -0.280 9.990 0.280 ;
        RECT  9.090 -0.280 9.370 0.440 ;
        RECT  8.040 -0.280 9.090 0.280 ;
        RECT  7.760 -0.280 8.040 0.430 ;
        RECT  6.320 -0.280 7.760 0.280 ;
        RECT  6.040 -0.280 6.320 0.880 ;
        RECT  4.580 -0.280 6.040 0.280 ;
        RECT  4.140 -0.280 4.580 0.620 ;
        RECT  1.810 -0.280 4.140 0.280 ;
        RECT  1.530 -0.280 1.810 0.740 ;
        RECT  0.440 -0.280 1.530 0.280 ;
        RECT  0.160 -0.280 0.440 0.380 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.260 3.320 12.400 3.880 ;
        RECT  12.070 2.120 12.260 3.880 ;
        RECT  11.300 3.320 12.070 3.880 ;
        RECT  11.020 2.930 11.300 3.880 ;
        RECT  10.240 3.320 11.020 3.880 ;
        RECT  9.960 3.130 10.240 3.880 ;
        RECT  8.730 3.320 9.960 3.880 ;
        RECT  8.040 3.240 8.730 3.880 ;
        RECT  6.390 3.320 8.040 3.880 ;
        RECT  5.780 3.240 6.390 3.880 ;
        RECT  4.850 3.320 5.780 3.880 ;
        RECT  3.850 3.240 4.850 3.880 ;
        RECT  1.780 3.320 3.850 3.880 ;
        RECT  1.500 2.850 1.780 3.880 ;
        RECT  0.380 3.320 1.500 3.880 ;
        RECT  0.100 3.200 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.370 1.500 11.500 1.780 ;
        RECT  11.340 1.500 11.370 2.750 ;
        RECT  11.200 1.510 11.340 2.750 ;
        RECT  10.060 2.590 11.200 2.750 ;
        RECT  10.010 2.580 10.060 2.750 ;
        RECT  9.850 1.010 10.010 2.750 ;
        RECT  9.620 1.010 9.850 1.290 ;
        RECT  9.720 2.580 9.850 2.750 ;
        RECT  9.440 2.580 9.720 2.860 ;
        RECT  9.210 1.680 9.670 1.990 ;
        RECT  9.280 2.700 9.440 2.860 ;
        RECT  9.120 2.700 9.280 3.080 ;
        RECT  9.050 1.100 9.210 2.280 ;
        RECT  9.000 2.880 9.120 3.080 ;
        RECT  8.570 1.100 9.050 1.260 ;
        RECT  8.700 2.120 9.050 2.280 ;
        RECT  3.500 2.880 9.000 3.040 ;
        RECT  8.570 1.470 8.730 1.960 ;
        RECT  8.530 2.120 8.700 2.700 ;
        RECT  8.350 1.070 8.570 1.260 ;
        RECT  8.270 1.800 8.570 1.960 ;
        RECT  7.130 2.540 8.530 2.700 ;
        RECT  7.690 1.070 8.350 1.230 ;
        RECT  8.110 1.800 8.270 2.300 ;
        RECT  7.340 1.480 8.150 1.640 ;
        RECT  7.230 2.140 8.110 2.300 ;
        RECT  7.530 0.700 7.690 1.230 ;
        RECT  7.160 0.700 7.530 0.860 ;
        RECT  7.180 1.090 7.340 1.640 ;
        RECT  6.960 2.080 7.230 2.360 ;
        RECT  6.750 1.090 7.180 1.250 ;
        RECT  6.880 0.580 7.160 0.860 ;
        RECT  6.950 2.080 6.960 2.720 ;
        RECT  6.800 2.200 6.950 2.720 ;
        RECT  4.460 2.560 6.800 2.720 ;
        RECT  6.630 1.080 6.750 1.250 ;
        RECT  6.470 1.080 6.630 2.340 ;
        RECT  5.660 1.080 6.470 1.240 ;
        RECT  5.740 2.180 6.470 2.340 ;
        RECT  6.140 1.740 6.300 2.020 ;
        RECT  5.460 1.800 6.140 1.960 ;
        RECT  5.500 0.440 5.660 1.240 ;
        RECT  4.850 0.440 5.500 0.600 ;
        RECT  5.450 1.800 5.460 2.330 ;
        RECT  5.300 1.400 5.450 2.330 ;
        RECT  5.290 1.200 5.300 2.330 ;
        RECT  5.140 1.200 5.290 1.560 ;
        RECT  3.820 2.170 5.290 2.330 ;
        RECT  4.990 1.200 5.140 1.360 ;
        RECT  4.800 1.730 5.120 1.890 ;
        RECT  4.640 0.880 4.800 1.890 ;
        RECT  3.320 0.880 4.640 1.040 ;
        RECT  4.180 2.520 4.460 2.720 ;
        RECT  3.750 1.230 4.240 1.390 ;
        RECT  3.500 2.560 4.180 2.720 ;
        RECT  3.660 2.050 3.820 2.330 ;
        RECT  3.590 1.230 3.750 1.540 ;
        RECT  3.340 1.380 3.590 1.540 ;
        RECT  3.340 2.220 3.500 2.720 ;
        RECT  3.340 2.880 3.500 3.160 ;
        RECT  3.180 1.380 3.340 2.380 ;
        RECT  2.200 3.000 3.340 3.160 ;
        RECT  3.200 0.600 3.320 1.040 ;
        RECT  3.040 0.600 3.200 1.150 ;
        RECT  2.710 1.380 3.180 1.540 ;
        RECT  3.120 2.220 3.180 2.380 ;
        RECT  2.940 2.600 3.180 2.760 ;
        RECT  2.540 0.990 3.040 1.150 ;
        RECT  2.780 1.880 2.940 2.760 ;
        RECT  2.540 1.880 2.780 2.040 ;
        RECT  2.160 0.660 2.720 0.820 ;
        RECT  2.440 2.530 2.600 2.830 ;
        RECT  2.380 0.990 2.540 2.040 ;
        RECT  0.900 2.530 2.440 2.690 ;
        RECT  2.000 0.660 2.160 1.090 ;
        RECT  1.730 1.260 2.010 1.540 ;
        RECT  1.280 0.930 2.000 1.090 ;
        RECT  1.640 1.270 1.730 1.540 ;
        RECT  1.480 1.270 1.640 2.280 ;
        RECT  0.910 1.270 1.480 1.430 ;
        RECT  0.580 2.120 1.480 2.280 ;
        RECT  1.120 0.620 1.280 1.090 ;
        RECT  0.630 0.620 1.120 0.780 ;
        RECT  0.720 1.030 0.910 1.430 ;
        RECT  0.680 2.530 0.900 2.820 ;
        RECT  0.630 1.030 0.720 1.320 ;
        RECT  0.630 2.540 0.680 2.820 ;
    END
END EDFFX4TR

MACRO EDFFX2TR
    CLASS CORE ;
    FOREIGN EDFFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 0.590 9.520 3.020 ;
        RECT  9.260 2.210 9.280 3.020 ;
        END
        ANTENNADIFFAREA 3.392 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.010 0.790 9.120 2.010 ;
        RECT  8.960 0.790 9.010 2.730 ;
        RECT  8.430 0.790 8.960 0.950 ;
        RECT  8.850 1.850 8.960 2.730 ;
        RECT  8.810 2.440 8.850 2.730 ;
        RECT  8.480 2.440 8.810 2.870 ;
        RECT  8.160 2.590 8.480 2.870 ;
        RECT  8.150 0.560 8.430 0.950 ;
        END
        ANTENNADIFFAREA 2.256 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.180 1.840 2.280 2.120 ;
        RECT  2.000 1.590 2.180 2.120 ;
        RECT  1.960 1.590 2.000 1.750 ;
        RECT  1.800 1.240 1.960 1.750 ;
        RECT  1.640 1.240 1.800 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.240 5.160 1.560 ;
        RECT  4.880 1.240 5.040 1.690 ;
        RECT  4.680 1.530 4.880 1.690 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.030 -0.280 9.600 0.280 ;
        RECT  8.750 -0.280 9.030 0.620 ;
        RECT  7.910 -0.280 8.750 0.280 ;
        RECT  7.630 -0.280 7.910 0.400 ;
        RECT  6.340 -0.280 7.630 0.340 ;
        RECT  6.120 -0.280 6.340 0.660 ;
        RECT  4.820 -0.280 6.120 0.280 ;
        RECT  4.540 -0.280 4.820 0.760 ;
        RECT  3.780 -0.280 4.540 0.280 ;
        RECT  3.500 -0.280 3.780 0.990 ;
        RECT  1.710 -0.280 3.500 0.280 ;
        RECT  1.430 -0.280 1.710 0.400 ;
        RECT  0.370 -0.280 1.430 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.960 3.320 9.600 3.880 ;
        RECT  8.680 3.200 8.960 3.880 ;
        RECT  7.920 3.320 8.680 3.880 ;
        RECT  7.640 2.560 7.920 3.880 ;
        RECT  5.570 3.260 7.640 3.880 ;
        RECT  4.100 3.320 5.570 3.880 ;
        RECT  3.720 3.200 4.100 3.880 ;
        RECT  1.690 3.260 3.720 3.880 ;
        RECT  1.410 3.200 1.690 3.880 ;
        RECT  0.370 3.320 1.410 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.720 1.410 8.770 1.690 ;
        RECT  8.640 1.110 8.720 1.690 ;
        RECT  8.480 1.110 8.640 2.220 ;
        RECT  8.230 1.110 8.480 1.340 ;
        RECT  7.420 1.980 8.480 2.220 ;
        RECT  7.960 1.500 8.240 1.780 ;
        RECT  7.130 1.620 7.960 1.780 ;
        RECT  7.220 1.980 7.420 3.100 ;
        RECT  7.110 0.700 7.390 0.980 ;
        RECT  4.420 2.940 7.220 3.100 ;
        RECT  6.980 1.140 7.130 1.780 ;
        RECT  6.500 0.820 7.110 0.980 ;
        RECT  6.820 1.140 6.980 2.780 ;
        RECT  6.660 2.500 6.820 2.780 ;
        RECT  6.500 2.060 6.620 2.340 ;
        RECT  6.340 0.820 6.500 2.780 ;
        RECT  5.960 0.820 6.340 0.980 ;
        RECT  4.740 2.560 6.340 2.780 ;
        RECT  6.020 1.220 6.180 2.400 ;
        RECT  5.630 1.220 6.020 1.380 ;
        RECT  5.320 2.240 6.020 2.400 ;
        RECT  5.800 0.440 5.960 0.980 ;
        RECT  5.640 1.740 5.860 2.020 ;
        RECT  5.140 0.440 5.800 0.600 ;
        RECT  4.400 1.860 5.640 2.020 ;
        RECT  5.580 1.100 5.630 1.380 ;
        RECT  5.410 0.760 5.580 1.380 ;
        RECT  5.300 0.760 5.410 0.980 ;
        RECT  5.040 2.180 5.320 2.400 ;
        RECT  4.980 0.440 5.140 1.080 ;
        RECT  4.720 0.920 4.980 1.080 ;
        RECT  4.580 2.430 4.740 2.780 ;
        RECT  4.500 0.920 4.720 1.370 ;
        RECT  2.740 2.430 4.580 2.650 ;
        RECT  4.260 2.810 4.420 3.100 ;
        RECT  4.340 1.860 4.400 2.270 ;
        RECT  4.180 0.630 4.340 2.270 ;
        RECT  0.770 2.810 4.260 3.030 ;
        RECT  4.060 0.630 4.180 1.310 ;
        RECT  3.650 1.150 4.060 1.310 ;
        RECT  3.800 1.520 4.020 1.800 ;
        RECT  3.120 1.640 3.800 1.800 ;
        RECT  3.370 1.150 3.650 1.430 ;
        RECT  3.100 1.640 3.120 2.270 ;
        RECT  2.900 0.440 3.100 2.270 ;
        RECT  2.620 0.440 2.900 0.720 ;
        RECT  2.580 1.350 2.740 2.650 ;
        RECT  2.410 1.350 2.580 1.630 ;
        RECT  2.160 0.440 2.440 0.850 ;
        RECT  2.200 2.370 2.420 2.650 ;
        RECT  0.810 2.490 2.200 2.650 ;
        RECT  0.830 0.690 2.160 0.850 ;
        RECT  1.450 2.040 1.840 2.320 ;
        RECT  1.290 1.280 1.450 2.320 ;
        RECT  1.170 1.280 1.290 1.560 ;
        RECT  0.810 1.280 1.170 1.440 ;
        RECT  0.550 0.570 0.830 0.850 ;
        RECT  0.650 1.030 0.810 2.190 ;
        RECT  0.530 2.370 0.810 2.650 ;
        RECT  0.530 1.030 0.650 1.360 ;
        RECT  0.530 1.910 0.650 2.190 ;
    END
END EDFFX2TR

MACRO EDFFX1TR
    CLASS CORE ;
    FOREIGN EDFFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.030 9.520 3.020 ;
        RECT  9.230 1.030 9.280 1.310 ;
        RECT  9.200 2.650 9.280 3.020 ;
        END
        ANTENNADIFFAREA 1.967 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.910 0.680 9.070 2.010 ;
        RECT  8.440 0.680 8.910 0.840 ;
        RECT  8.880 1.850 8.910 2.010 ;
        RECT  8.720 1.850 8.880 2.870 ;
        RECT  8.440 2.440 8.720 2.870 ;
        RECT  8.160 0.560 8.440 0.840 ;
        RECT  8.160 2.590 8.440 2.870 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.580 0.340 2.760 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.840 2.250 2.120 ;
        RECT  1.970 1.590 2.130 2.120 ;
        RECT  1.960 1.590 1.970 1.750 ;
        RECT  1.800 1.240 1.960 1.750 ;
        RECT  1.640 1.240 1.800 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.160 1.690 ;
        RECT  4.680 1.530 4.880 1.690 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.020 -0.280 9.600 0.280 ;
        RECT  8.740 -0.280 9.020 0.400 ;
        RECT  7.920 -0.280 8.740 0.280 ;
        RECT  7.640 -0.280 7.920 0.790 ;
        RECT  6.340 -0.280 7.640 0.340 ;
        RECT  6.060 -0.280 6.340 0.660 ;
        RECT  4.820 -0.280 6.060 0.280 ;
        RECT  4.540 -0.280 4.820 0.760 ;
        RECT  3.780 -0.280 4.540 0.280 ;
        RECT  3.500 -0.280 3.780 0.990 ;
        RECT  1.710 -0.280 3.500 0.280 ;
        RECT  1.430 -0.280 1.710 0.400 ;
        RECT  0.370 -0.280 1.430 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.900 3.320 9.600 3.880 ;
        RECT  8.620 3.200 8.900 3.880 ;
        RECT  7.920 3.320 8.620 3.880 ;
        RECT  7.640 2.560 7.920 3.880 ;
        RECT  5.570 3.260 7.640 3.880 ;
        RECT  3.080 3.320 5.570 3.880 ;
        RECT  1.690 3.260 3.080 3.880 ;
        RECT  1.410 3.200 1.690 3.880 ;
        RECT  0.370 3.320 1.410 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.640 1.410 8.750 1.690 ;
        RECT  8.560 1.050 8.640 1.690 ;
        RECT  8.400 1.050 8.560 2.220 ;
        RECT  8.240 1.050 8.400 1.340 ;
        RECT  7.420 1.980 8.400 2.220 ;
        RECT  7.960 1.500 8.240 1.780 ;
        RECT  7.130 1.620 7.960 1.780 ;
        RECT  7.220 1.980 7.420 3.100 ;
        RECT  7.120 0.700 7.400 0.980 ;
        RECT  5.320 2.940 7.220 3.100 ;
        RECT  6.980 1.140 7.130 1.780 ;
        RECT  6.460 0.820 7.120 0.980 ;
        RECT  6.840 1.140 6.980 2.660 ;
        RECT  6.820 1.140 6.840 2.780 ;
        RECT  6.620 2.500 6.820 2.780 ;
        RECT  6.460 2.060 6.620 2.340 ;
        RECT  6.300 0.820 6.460 2.780 ;
        RECT  5.900 0.820 6.300 0.980 ;
        RECT  4.820 2.560 6.300 2.780 ;
        RECT  5.980 1.220 6.140 2.400 ;
        RECT  5.620 1.220 5.980 1.380 ;
        RECT  5.310 2.240 5.980 2.400 ;
        RECT  5.740 0.440 5.900 0.980 ;
        RECT  5.480 1.740 5.820 2.020 ;
        RECT  5.140 0.440 5.740 0.600 ;
        RECT  5.580 1.100 5.620 1.380 ;
        RECT  5.340 0.760 5.580 1.380 ;
        RECT  4.460 1.860 5.480 2.020 ;
        RECT  5.300 0.760 5.340 0.980 ;
        RECT  5.160 2.940 5.320 3.160 ;
        RECT  5.030 2.180 5.310 2.400 ;
        RECT  4.120 3.000 5.160 3.160 ;
        RECT  4.980 0.440 5.140 1.080 ;
        RECT  4.720 0.920 4.980 1.080 ;
        RECT  4.810 2.430 4.820 2.780 ;
        RECT  4.530 2.430 4.810 2.840 ;
        RECT  4.500 0.920 4.720 1.370 ;
        RECT  2.710 2.430 4.530 2.650 ;
        RECT  4.340 1.860 4.460 2.250 ;
        RECT  4.180 0.630 4.340 2.250 ;
        RECT  4.060 0.630 4.180 1.310 ;
        RECT  3.960 2.810 4.120 3.160 ;
        RECT  3.650 1.150 4.060 1.310 ;
        RECT  3.800 1.520 4.020 1.800 ;
        RECT  0.770 2.810 3.960 3.030 ;
        RECT  3.090 1.640 3.800 1.800 ;
        RECT  3.370 1.150 3.650 1.430 ;
        RECT  3.030 1.640 3.090 2.270 ;
        RECT  2.870 0.440 3.030 2.270 ;
        RECT  2.620 0.440 2.870 0.720 ;
        RECT  2.550 1.350 2.710 2.650 ;
        RECT  2.410 1.350 2.550 1.630 ;
        RECT  2.170 2.370 2.390 2.650 ;
        RECT  2.090 0.440 2.370 0.850 ;
        RECT  0.810 2.490 2.170 2.650 ;
        RECT  0.830 0.690 2.090 0.850 ;
        RECT  1.450 2.040 1.810 2.320 ;
        RECT  1.290 1.280 1.450 2.320 ;
        RECT  1.170 1.280 1.290 1.560 ;
        RECT  0.810 1.280 1.170 1.440 ;
        RECT  0.550 0.570 0.830 0.850 ;
        RECT  0.650 1.030 0.810 2.190 ;
        RECT  0.530 2.370 0.810 2.650 ;
        RECT  0.530 1.030 0.650 1.360 ;
        RECT  0.530 1.910 0.650 2.190 ;
    END
END EDFFX1TR

MACRO DLY4X4TR
    CLASS CORE ;
    FOREIGN DLY4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.040 4.290 2.150 ;
        RECT  4.020 1.040 4.050 1.310 ;
        RECT  3.820 1.910 4.050 2.150 ;
        RECT  3.740 0.500 4.020 1.310 ;
        RECT  3.550 1.910 3.820 3.160 ;
        RECT  3.280 2.240 3.550 2.960 ;
        END
        ANTENNADIFFAREA 3.85 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.280 4.400 0.280 ;
        RECT  3.180 -0.280 3.460 1.310 ;
        RECT  0.900 -0.280 3.180 0.280 ;
        RECT  0.620 -0.280 0.900 0.420 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.400 3.880 ;
        RECT  4.030 2.390 4.310 3.880 ;
        RECT  3.310 3.320 4.030 3.880 ;
        RECT  3.030 3.200 3.310 3.880 ;
        RECT  0.860 3.320 3.030 3.880 ;
        RECT  0.580 3.190 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 1.470 3.680 1.750 ;
        RECT  2.860 1.230 3.020 2.150 ;
        RECT  2.330 1.230 2.860 1.390 ;
        RECT  2.360 1.990 2.860 2.150 ;
        RECT  2.440 1.550 2.700 1.830 ;
        RECT  1.900 1.550 2.440 1.710 ;
        RECT  2.080 1.990 2.360 2.710 ;
        RECT  2.080 1.030 2.330 1.390 ;
        RECT  1.620 1.030 1.900 2.710 ;
        RECT  1.080 1.360 1.220 1.640 ;
        RECT  0.920 0.920 1.080 2.070 ;
        RECT  0.370 0.920 0.920 1.080 ;
        RECT  0.370 1.910 0.920 2.070 ;
        RECT  0.090 0.790 0.370 1.080 ;
        RECT  0.090 1.910 0.370 2.700 ;
    END
END DLY4X4TR

MACRO DLY4X1TR
    CLASS CORE ;
    FOREIGN DLY4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.240 3.920 2.360 ;
        RECT  3.800 1.240 3.830 2.550 ;
        RECT  3.640 1.000 3.800 2.550 ;
        RECT  3.560 1.000 3.640 1.280 ;
        RECT  3.390 1.910 3.640 2.550 ;
        END
        ANTENNADIFFAREA 1.636 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.280 4.000 0.280 ;
        RECT  3.000 -0.280 3.280 0.340 ;
        RECT  0.900 -0.280 3.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.410 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 3.320 4.000 3.880 ;
        RECT  3.000 3.200 3.280 3.880 ;
        RECT  0.900 3.320 3.000 3.880 ;
        RECT  0.620 3.170 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 1.390 3.420 1.670 ;
        RECT  2.760 1.150 2.920 2.070 ;
        RECT  2.320 1.150 2.760 1.310 ;
        RECT  2.320 1.910 2.760 2.070 ;
        RECT  2.320 1.470 2.600 1.750 ;
        RECT  2.040 1.030 2.320 1.310 ;
        RECT  1.860 1.470 2.320 1.630 ;
        RECT  2.040 1.910 2.320 2.710 ;
        RECT  1.700 1.030 1.860 2.710 ;
        RECT  1.580 1.030 1.700 1.310 ;
        RECT  1.580 1.910 1.700 2.710 ;
        RECT  1.100 1.580 1.220 1.860 ;
        RECT  0.940 1.580 1.100 2.070 ;
        RECT  0.380 1.910 0.940 2.070 ;
        RECT  0.240 1.910 0.380 2.710 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.080 1.030 0.240 2.710 ;
    END
END DLY4X1TR

MACRO DLY3X4TR
    CLASS CORE ;
    FOREIGN DLY3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.040 4.290 2.150 ;
        RECT  4.020 1.040 4.050 1.310 ;
        RECT  3.820 1.910 4.050 2.150 ;
        RECT  3.740 0.500 4.020 1.310 ;
        RECT  3.550 1.910 3.820 3.160 ;
        RECT  3.280 2.240 3.550 2.960 ;
        END
        ANTENNADIFFAREA 3.85 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.280 4.400 0.280 ;
        RECT  3.180 -0.280 3.460 1.310 ;
        RECT  0.940 -0.280 3.180 0.280 ;
        RECT  0.660 -0.280 0.940 0.420 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.400 3.880 ;
        RECT  4.030 2.390 4.310 3.880 ;
        RECT  3.310 3.320 4.030 3.880 ;
        RECT  3.030 3.200 3.310 3.880 ;
        RECT  0.940 3.320 3.030 3.880 ;
        RECT  0.660 2.290 0.940 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 1.470 3.680 1.750 ;
        RECT  2.860 1.230 3.020 2.150 ;
        RECT  2.330 1.230 2.860 1.390 ;
        RECT  2.360 1.990 2.860 2.150 ;
        RECT  2.440 1.550 2.700 1.830 ;
        RECT  1.900 1.550 2.440 1.710 ;
        RECT  2.080 1.990 2.360 2.710 ;
        RECT  2.080 1.030 2.330 1.390 ;
        RECT  1.620 1.030 1.900 2.710 ;
        RECT  1.080 1.360 1.250 1.640 ;
        RECT  0.920 0.920 1.080 2.070 ;
        RECT  0.370 0.920 0.920 1.080 ;
        RECT  0.370 1.910 0.920 2.070 ;
        RECT  0.090 0.790 0.370 1.080 ;
        RECT  0.090 1.910 0.370 2.700 ;
    END
END DLY3X4TR

MACRO DLY3X1TR
    CLASS CORE ;
    FOREIGN DLY3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.000 3.920 2.360 ;
        RECT  3.640 1.000 3.830 2.550 ;
        RECT  3.560 1.000 3.640 1.280 ;
        RECT  3.510 1.910 3.640 2.550 ;
        END
        ANTENNADIFFAREA 1.636 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.280 4.000 0.280 ;
        RECT  3.000 -0.280 3.280 0.830 ;
        RECT  0.900 -0.280 3.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.810 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 3.320 4.000 3.880 ;
        RECT  3.000 2.370 3.280 3.880 ;
        RECT  0.900 3.320 3.000 3.880 ;
        RECT  0.620 2.370 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 1.390 3.420 1.670 ;
        RECT  2.760 1.150 2.920 2.070 ;
        RECT  2.320 1.150 2.760 1.310 ;
        RECT  2.320 1.910 2.760 2.070 ;
        RECT  2.320 1.470 2.600 1.750 ;
        RECT  2.040 1.030 2.320 1.310 ;
        RECT  1.860 1.470 2.320 1.630 ;
        RECT  2.040 1.910 2.320 2.630 ;
        RECT  1.700 1.030 1.860 2.630 ;
        RECT  1.580 1.030 1.700 1.310 ;
        RECT  1.580 1.910 1.700 2.630 ;
        RECT  1.100 1.580 1.220 1.860 ;
        RECT  0.940 1.580 1.100 2.070 ;
        RECT  0.380 1.910 0.940 2.070 ;
        RECT  0.240 1.910 0.380 2.630 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.080 1.030 0.240 2.630 ;
    END
END DLY3X1TR

MACRO DLY2X4TR
    CLASS CORE ;
    FOREIGN DLY2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.040 4.290 2.150 ;
        RECT  4.020 1.040 4.050 1.310 ;
        RECT  3.820 1.910 4.050 2.150 ;
        RECT  3.740 0.500 4.020 1.310 ;
        RECT  3.550 1.910 3.820 3.160 ;
        RECT  3.280 2.240 3.550 2.960 ;
        END
        ANTENNADIFFAREA 3.85 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.280 4.400 0.280 ;
        RECT  3.180 -0.280 3.460 1.310 ;
        RECT  0.940 -0.280 3.180 0.280 ;
        RECT  0.660 -0.280 0.940 0.420 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.400 3.880 ;
        RECT  4.030 2.390 4.310 3.880 ;
        RECT  3.310 3.320 4.030 3.880 ;
        RECT  3.120 3.200 3.310 3.880 ;
        RECT  2.880 2.380 3.120 3.880 ;
        RECT  0.940 3.320 2.880 3.880 ;
        RECT  0.660 2.340 0.940 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 1.470 3.680 1.750 ;
        RECT  2.860 1.230 3.020 2.150 ;
        RECT  2.330 1.230 2.860 1.390 ;
        RECT  2.360 1.990 2.860 2.150 ;
        RECT  2.440 1.550 2.700 1.830 ;
        RECT  1.720 1.550 2.440 1.710 ;
        RECT  2.080 1.990 2.360 2.710 ;
        RECT  2.080 1.030 2.330 1.390 ;
        RECT  1.440 1.030 1.720 2.710 ;
        RECT  1.080 1.360 1.250 1.640 ;
        RECT  0.920 0.920 1.080 2.070 ;
        RECT  0.370 0.920 0.920 1.080 ;
        RECT  0.370 1.910 0.920 2.070 ;
        RECT  0.090 0.790 0.370 1.080 ;
        RECT  0.090 1.910 0.370 2.700 ;
    END
END DLY2X4TR

MACRO DLY2X1TR
    CLASS CORE ;
    FOREIGN DLY2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.240 3.920 2.360 ;
        RECT  3.800 1.240 3.830 2.550 ;
        RECT  3.640 1.000 3.800 2.550 ;
        RECT  3.560 1.000 3.640 1.280 ;
        RECT  3.450 1.910 3.640 2.550 ;
        END
        ANTENNADIFFAREA 1.636 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.280 4.000 0.280 ;
        RECT  3.000 -0.280 3.280 0.910 ;
        RECT  0.940 -0.280 3.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.860 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 3.320 4.000 3.880 ;
        RECT  3.000 2.330 3.280 3.880 ;
        RECT  0.900 3.320 3.000 3.880 ;
        RECT  0.620 2.350 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 1.390 3.420 1.670 ;
        RECT  2.760 1.150 2.920 2.070 ;
        RECT  2.320 1.150 2.760 1.310 ;
        RECT  2.320 1.910 2.760 2.070 ;
        RECT  2.320 1.470 2.600 1.750 ;
        RECT  2.040 1.030 2.320 1.310 ;
        RECT  1.860 1.470 2.320 1.630 ;
        RECT  2.040 1.910 2.320 2.630 ;
        RECT  1.700 1.030 1.860 2.630 ;
        RECT  1.580 1.030 1.700 1.310 ;
        RECT  1.580 1.910 1.700 2.630 ;
        RECT  1.100 1.580 1.220 1.860 ;
        RECT  0.940 1.580 1.100 2.070 ;
        RECT  0.380 1.910 0.940 2.070 ;
        RECT  0.240 1.910 0.380 2.630 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.080 1.030 0.240 2.630 ;
    END
END DLY2X1TR

MACRO DLY1X4TR
    CLASS CORE ;
    FOREIGN DLY1X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.040 4.290 2.150 ;
        RECT  4.020 1.040 4.050 1.310 ;
        RECT  3.820 1.910 4.050 2.150 ;
        RECT  3.740 0.500 4.020 1.310 ;
        RECT  3.550 1.910 3.820 3.160 ;
        RECT  3.280 2.240 3.550 2.960 ;
        END
        ANTENNADIFFAREA 3.85 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.280 4.400 0.280 ;
        RECT  3.180 -0.280 3.460 1.310 ;
        RECT  0.940 -0.280 3.180 0.280 ;
        RECT  0.660 -0.280 0.940 0.420 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.400 3.880 ;
        RECT  4.030 2.390 4.310 3.880 ;
        RECT  3.310 3.320 4.030 3.880 ;
        RECT  3.120 3.200 3.310 3.880 ;
        RECT  2.880 2.380 3.120 3.880 ;
        RECT  0.940 3.320 2.880 3.880 ;
        RECT  0.660 2.340 0.940 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 1.470 3.680 1.750 ;
        RECT  2.860 1.230 3.020 2.150 ;
        RECT  2.630 1.230 2.860 1.390 ;
        RECT  2.640 1.990 2.860 2.150 ;
        RECT  2.440 1.550 2.700 1.830 ;
        RECT  2.340 1.990 2.640 2.710 ;
        RECT  2.340 1.030 2.630 1.390 ;
        RECT  1.560 1.550 2.440 1.710 ;
        RECT  1.280 1.030 1.560 2.710 ;
        RECT  1.080 1.360 1.120 1.640 ;
        RECT  0.920 0.920 1.080 2.070 ;
        RECT  0.370 0.920 0.920 1.080 ;
        RECT  0.370 1.910 0.920 2.070 ;
        RECT  0.090 0.790 0.370 1.080 ;
        RECT  0.090 1.910 0.370 2.700 ;
    END
END DLY1X4TR

MACRO DLY1X1TR
    CLASS CORE ;
    FOREIGN DLY1X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.240 3.920 2.360 ;
        RECT  3.800 1.240 3.830 2.550 ;
        RECT  3.640 1.000 3.800 2.550 ;
        RECT  3.560 1.000 3.640 1.280 ;
        RECT  3.480 1.910 3.640 2.550 ;
        END
        ANTENNADIFFAREA 1.636 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.280 4.000 0.280 ;
        RECT  3.000 -0.280 3.280 0.910 ;
        RECT  0.940 -0.280 3.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.860 ;
        RECT  0.000 -0.280 0.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 3.320 4.000 3.880 ;
        RECT  3.000 2.330 3.280 3.880 ;
        RECT  0.900 3.320 3.000 3.880 ;
        RECT  0.620 2.350 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 1.390 3.420 1.670 ;
        RECT  2.990 1.150 3.150 2.070 ;
        RECT  2.550 1.150 2.990 1.310 ;
        RECT  2.550 1.910 2.990 2.070 ;
        RECT  2.550 1.470 2.830 1.750 ;
        RECT  2.270 1.030 2.550 1.310 ;
        RECT  1.640 1.470 2.550 1.630 ;
        RECT  2.270 1.910 2.550 2.630 ;
        RECT  1.480 1.030 1.640 2.630 ;
        RECT  1.360 1.030 1.480 1.310 ;
        RECT  1.360 1.910 1.480 2.630 ;
        RECT  1.010 1.580 1.200 2.070 ;
        RECT  0.380 1.910 1.010 2.070 ;
        RECT  0.240 1.910 0.380 2.630 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.080 1.030 0.240 2.630 ;
    END
END DLY1X1TR

MACRO DFFTRXLTR
    CLASS CORE ;
    FOREIGN DFFTRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.220 1.520 1.700 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.840 8.320 2.250 ;
        END
        ANTENNADIFFAREA 1.1 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.030 7.520 2.270 ;
        RECT  6.980 1.030 7.280 1.310 ;
        RECT  6.800 1.910 7.280 2.270 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.220 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.760 -0.280 8.400 0.280 ;
        RECT  7.480 -0.280 7.760 0.400 ;
        RECT  6.500 -0.280 7.480 0.280 ;
        RECT  6.020 -0.280 6.500 0.670 ;
        RECT  4.420 -0.280 6.020 0.340 ;
        RECT  4.140 -0.280 4.420 0.990 ;
        RECT  2.520 -0.280 4.140 0.340 ;
        RECT  2.240 -0.280 2.520 0.400 ;
        RECT  1.620 -0.280 2.240 0.280 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  0.730 -0.280 1.340 0.340 ;
        RECT  0.000 -0.280 0.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.760 3.320 8.400 3.880 ;
        RECT  7.290 3.260 7.760 3.880 ;
        RECT  6.380 3.320 7.290 3.880 ;
        RECT  6.080 2.850 6.380 3.880 ;
        RECT  4.000 3.260 6.080 3.880 ;
        RECT  3.720 2.400 4.000 3.880 ;
        RECT  2.520 3.260 3.720 3.880 ;
        RECT  2.240 3.210 2.520 3.880 ;
        RECT  1.400 3.320 2.240 3.880 ;
        RECT  1.120 3.210 1.400 3.880 ;
        RECT  0.470 3.260 1.120 3.880 ;
        RECT  0.000 3.320 0.470 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.760 0.710 7.920 3.090 ;
        RECT  7.060 0.710 7.760 0.870 ;
        RECT  6.900 2.930 7.760 3.090 ;
        RECT  6.740 1.560 7.120 1.720 ;
        RECT  6.780 0.450 7.060 0.870 ;
        RECT  6.620 2.930 6.900 3.150 ;
        RECT  6.640 1.030 6.740 1.720 ;
        RECT  6.480 1.030 6.640 2.620 ;
        RECT  6.460 1.030 6.480 1.720 ;
        RECT  6.300 2.340 6.480 2.620 ;
        RECT  5.780 1.560 6.460 1.720 ;
        RECT  5.340 1.900 6.320 2.180 ;
        RECT  5.340 0.580 5.540 0.820 ;
        RECT  5.220 2.710 5.500 2.990 ;
        RECT  5.260 0.580 5.340 2.180 ;
        RECT  5.180 0.580 5.260 2.500 ;
        RECT  4.400 2.710 5.220 2.870 ;
        RECT  5.100 1.900 5.180 2.500 ;
        RECT  4.980 2.220 5.100 2.500 ;
        RECT  4.820 0.730 4.940 1.010 ;
        RECT  4.780 0.730 4.820 1.310 ;
        RECT  4.660 0.730 4.780 2.540 ;
        RECT  4.560 1.150 4.660 2.540 ;
        RECT  4.300 1.150 4.560 1.310 ;
        RECT  4.240 1.590 4.400 2.870 ;
        RECT  4.020 1.150 4.300 1.430 ;
        RECT  3.860 1.590 4.240 1.750 ;
        RECT  3.540 1.910 4.080 2.190 ;
        RECT  3.780 0.620 3.860 1.750 ;
        RECT  3.700 0.500 3.780 1.750 ;
        RECT  3.100 0.500 3.700 0.780 ;
        RECT  3.420 0.940 3.540 2.190 ;
        RECT  3.260 0.940 3.420 2.680 ;
        RECT  2.960 2.440 3.260 2.680 ;
        RECT  2.940 0.500 3.100 2.280 ;
        RECT  2.800 2.440 2.960 3.050 ;
        RECT  2.800 0.780 2.940 1.060 ;
        RECT  2.800 1.910 2.940 2.280 ;
        RECT  0.680 2.120 2.800 2.280 ;
        RECT  0.370 2.890 2.800 3.050 ;
        RECT  2.640 1.220 2.780 1.500 ;
        RECT  2.480 0.900 2.640 1.940 ;
        RECT  2.080 0.900 2.480 1.060 ;
        RECT  1.680 1.720 2.480 1.940 ;
        RECT  1.800 0.780 2.080 1.060 ;
        RECT  0.600 2.460 1.920 2.730 ;
        RECT  0.800 0.900 1.800 1.060 ;
        RECT  0.640 0.500 0.800 1.060 ;
        RECT  0.400 1.980 0.680 2.280 ;
        RECT  0.440 0.500 0.640 0.780 ;
        RECT  0.240 0.940 0.480 1.220 ;
        RECT  0.240 2.440 0.370 3.050 ;
        RECT  0.210 0.940 0.240 3.050 ;
        RECT  0.080 0.940 0.210 2.720 ;
    END
END DFFTRXLTR

MACRO DFFTRX4TR
    CLASS CORE ;
    FOREIGN DFFTRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.220 1.520 1.700 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.630 1.040 8.720 2.370 ;
        RECT  8.480 0.520 8.630 3.110 ;
        RECT  8.410 0.520 8.480 1.200 ;
        RECT  8.410 2.090 8.480 3.110 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.090 7.920 2.430 ;
        RECT  7.390 1.090 7.680 1.310 ;
        RECT  7.440 2.150 7.680 2.430 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.220 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 -0.280 9.200 0.280 ;
        RECT  8.880 -0.280 9.110 1.070 ;
        RECT  8.150 -0.280 8.880 0.280 ;
        RECT  7.870 -0.280 8.150 0.610 ;
        RECT  7.190 -0.280 7.870 0.280 ;
        RECT  6.910 -0.280 7.190 0.610 ;
        RECT  6.130 -0.280 6.910 0.280 ;
        RECT  5.850 -0.280 6.130 0.400 ;
        RECT  4.300 -0.280 5.850 0.340 ;
        RECT  4.020 -0.280 4.300 0.990 ;
        RECT  2.520 -0.280 4.020 0.340 ;
        RECT  2.240 -0.280 2.520 0.400 ;
        RECT  1.620 -0.280 2.240 0.280 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  0.730 -0.280 1.340 0.340 ;
        RECT  0.000 -0.280 0.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 3.320 9.200 3.880 ;
        RECT  8.890 2.050 9.110 3.880 ;
        RECT  8.830 2.600 8.890 3.880 ;
        RECT  8.150 3.320 8.830 3.880 ;
        RECT  7.870 2.930 8.150 3.880 ;
        RECT  7.190 3.320 7.870 3.880 ;
        RECT  6.910 2.930 7.190 3.880 ;
        RECT  5.970 3.320 6.910 3.880 ;
        RECT  5.690 3.200 5.970 3.880 ;
        RECT  4.000 3.320 5.690 3.880 ;
        RECT  3.720 2.400 4.000 3.880 ;
        RECT  2.520 3.260 3.720 3.880 ;
        RECT  2.240 3.230 2.520 3.880 ;
        RECT  1.400 3.320 2.240 3.880 ;
        RECT  1.120 3.230 1.400 3.880 ;
        RECT  0.470 3.260 1.120 3.880 ;
        RECT  0.000 3.320 0.470 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.240 1.360 8.320 1.640 ;
        RECT  8.080 0.770 8.240 2.750 ;
        RECT  6.710 0.770 8.080 0.930 ;
        RECT  6.670 2.590 8.080 2.750 ;
        RECT  7.040 1.520 7.520 1.680 ;
        RECT  6.880 1.090 7.040 2.430 ;
        RECT  5.960 1.090 6.880 1.250 ;
        RECT  6.300 2.190 6.880 2.430 ;
        RECT  6.430 0.450 6.710 0.930 ;
        RECT  6.510 2.590 6.670 3.150 ;
        RECT  6.390 2.910 6.510 3.150 ;
        RECT  6.120 1.740 6.400 2.030 ;
        RECT  5.300 1.870 6.120 2.030 ;
        RECT  5.680 1.090 5.960 1.680 ;
        RECT  5.140 2.710 5.420 3.160 ;
        RECT  5.040 0.920 5.300 2.300 ;
        RECT  4.400 2.710 5.140 2.870 ;
        RECT  4.720 0.730 4.860 1.010 ;
        RECT  4.560 0.730 4.720 2.540 ;
        RECT  4.180 1.150 4.560 1.310 ;
        RECT  4.240 1.590 4.400 2.870 ;
        RECT  3.680 1.590 4.240 1.750 ;
        RECT  3.900 1.150 4.180 1.430 ;
        RECT  3.420 1.910 4.080 2.190 ;
        RECT  3.520 0.500 3.680 1.750 ;
        RECT  3.040 0.500 3.520 0.740 ;
        RECT  3.360 1.910 3.420 2.680 ;
        RECT  3.200 1.030 3.360 2.680 ;
        RECT  2.960 2.440 3.200 2.680 ;
        RECT  2.880 0.500 3.040 2.280 ;
        RECT  2.800 2.440 2.960 3.070 ;
        RECT  2.800 0.500 2.880 0.850 ;
        RECT  2.800 1.910 2.880 2.280 ;
        RECT  0.680 2.120 2.800 2.280 ;
        RECT  0.370 2.910 2.800 3.070 ;
        RECT  2.640 1.220 2.720 1.500 ;
        RECT  2.480 0.900 2.640 1.940 ;
        RECT  2.080 0.900 2.480 1.060 ;
        RECT  1.680 1.720 2.480 1.940 ;
        RECT  1.800 0.780 2.080 1.060 ;
        RECT  0.600 2.460 1.920 2.750 ;
        RECT  0.800 0.900 1.800 1.060 ;
        RECT  0.640 0.500 0.800 1.060 ;
        RECT  0.400 1.980 0.680 2.280 ;
        RECT  0.440 0.500 0.640 0.780 ;
        RECT  0.240 0.940 0.480 1.220 ;
        RECT  0.240 2.440 0.370 3.070 ;
        RECT  0.210 0.940 0.240 3.070 ;
        RECT  0.080 0.940 0.210 2.720 ;
    END
END DFFTRX4TR

MACRO DFFTRX2TR
    CLASS CORE ;
    FOREIGN DFFTRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.220 1.520 1.700 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.500 8.320 2.890 ;
        END
        ANTENNADIFFAREA 3.804 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.090 7.520 2.270 ;
        RECT  7.040 1.090 7.280 1.310 ;
        RECT  7.040 1.910 7.280 2.270 ;
        END
        ANTENNADIFFAREA 3.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.220 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 -0.280 8.400 0.280 ;
        RECT  7.520 -0.280 7.800 0.610 ;
        RECT  6.400 -0.280 7.520 0.280 ;
        RECT  5.920 -0.280 6.400 0.400 ;
        RECT  4.300 -0.280 5.920 0.340 ;
        RECT  4.020 -0.280 4.300 0.990 ;
        RECT  2.520 -0.280 4.020 0.340 ;
        RECT  2.240 -0.280 2.520 0.400 ;
        RECT  1.620 -0.280 2.240 0.280 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  0.730 -0.280 1.340 0.340 ;
        RECT  0.000 -0.280 0.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 3.320 8.400 3.880 ;
        RECT  7.520 2.990 7.800 3.880 ;
        RECT  6.370 3.320 7.520 3.880 ;
        RECT  6.090 2.850 6.370 3.880 ;
        RECT  4.000 3.260 6.090 3.880 ;
        RECT  3.720 2.400 4.000 3.880 ;
        RECT  2.520 3.260 3.720 3.880 ;
        RECT  2.240 3.210 2.520 3.880 ;
        RECT  1.400 3.320 2.240 3.880 ;
        RECT  1.120 3.210 1.400 3.880 ;
        RECT  0.470 3.260 1.120 3.880 ;
        RECT  0.000 3.320 0.470 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.760 0.770 7.920 2.810 ;
        RECT  6.960 0.770 7.760 0.930 ;
        RECT  6.920 2.650 7.760 2.810 ;
        RECT  6.640 1.560 7.120 1.720 ;
        RECT  6.680 0.450 6.960 0.930 ;
        RECT  6.760 2.650 6.920 3.150 ;
        RECT  6.580 2.910 6.760 3.150 ;
        RECT  6.600 1.090 6.640 1.720 ;
        RECT  6.440 1.090 6.600 2.600 ;
        RECT  6.360 1.090 6.440 1.720 ;
        RECT  6.300 2.340 6.440 2.600 ;
        RECT  5.680 1.560 6.360 1.720 ;
        RECT  5.320 1.900 6.280 2.180 ;
        RECT  5.220 2.710 5.500 2.990 ;
        RECT  5.260 0.920 5.320 2.180 ;
        RECT  5.040 0.920 5.260 2.500 ;
        RECT  4.400 2.710 5.220 2.870 ;
        RECT  4.980 2.220 5.040 2.500 ;
        RECT  4.720 0.730 4.860 1.010 ;
        RECT  4.560 0.730 4.720 2.540 ;
        RECT  4.180 1.150 4.560 1.310 ;
        RECT  4.240 1.590 4.400 2.870 ;
        RECT  3.680 1.590 4.240 1.750 ;
        RECT  3.900 1.150 4.180 1.430 ;
        RECT  3.420 1.910 4.080 2.190 ;
        RECT  3.520 0.500 3.680 1.750 ;
        RECT  3.040 0.500 3.520 0.780 ;
        RECT  3.360 1.910 3.420 2.680 ;
        RECT  3.200 1.030 3.360 2.680 ;
        RECT  2.960 2.440 3.200 2.680 ;
        RECT  2.940 0.500 3.040 2.280 ;
        RECT  2.800 2.440 2.960 3.050 ;
        RECT  2.880 0.570 2.940 2.280 ;
        RECT  2.800 0.570 2.880 0.850 ;
        RECT  2.800 1.910 2.880 2.280 ;
        RECT  0.680 2.120 2.800 2.280 ;
        RECT  0.370 2.890 2.800 3.050 ;
        RECT  2.640 1.220 2.720 1.500 ;
        RECT  2.480 0.900 2.640 1.940 ;
        RECT  2.080 0.900 2.480 1.060 ;
        RECT  1.680 1.720 2.480 1.940 ;
        RECT  1.800 0.780 2.080 1.060 ;
        RECT  0.600 2.460 1.920 2.730 ;
        RECT  0.800 0.900 1.800 1.060 ;
        RECT  0.640 0.500 0.800 1.060 ;
        RECT  0.400 1.980 0.680 2.280 ;
        RECT  0.440 0.500 0.640 0.780 ;
        RECT  0.240 0.940 0.480 1.220 ;
        RECT  0.240 2.440 0.370 3.050 ;
        RECT  0.210 0.940 0.240 3.050 ;
        RECT  0.080 0.940 0.210 2.720 ;
    END
END DFFTRX2TR

MACRO DFFTRX1TR
    CLASS CORE ;
    FOREIGN DFFTRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.220 1.520 1.700 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.840 8.320 2.250 ;
        END
        ANTENNADIFFAREA 1.98 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.030 7.520 2.270 ;
        RECT  6.980 1.030 7.280 1.310 ;
        RECT  6.800 1.910 7.280 2.270 ;
        END
        ANTENNADIFFAREA 1.852 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.220 2.320 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.760 -0.280 8.400 0.280 ;
        RECT  7.480 -0.280 7.760 0.400 ;
        RECT  6.500 -0.280 7.480 0.280 ;
        RECT  6.020 -0.280 6.500 0.670 ;
        RECT  4.420 -0.280 6.020 0.340 ;
        RECT  4.140 -0.280 4.420 0.990 ;
        RECT  2.520 -0.280 4.140 0.340 ;
        RECT  2.240 -0.280 2.520 0.400 ;
        RECT  1.620 -0.280 2.240 0.280 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  0.730 -0.280 1.340 0.340 ;
        RECT  0.000 -0.280 0.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.760 3.320 8.400 3.880 ;
        RECT  7.290 3.260 7.760 3.880 ;
        RECT  6.390 3.320 7.290 3.880 ;
        RECT  6.070 2.850 6.390 3.880 ;
        RECT  4.000 3.260 6.070 3.880 ;
        RECT  3.720 2.400 4.000 3.880 ;
        RECT  2.520 3.260 3.720 3.880 ;
        RECT  2.240 3.210 2.520 3.880 ;
        RECT  1.400 3.320 2.240 3.880 ;
        RECT  1.120 3.210 1.400 3.880 ;
        RECT  0.470 3.260 1.120 3.880 ;
        RECT  0.000 3.320 0.470 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.760 0.710 7.920 3.090 ;
        RECT  7.060 0.710 7.760 0.870 ;
        RECT  6.900 2.930 7.760 3.090 ;
        RECT  6.740 1.560 7.120 1.720 ;
        RECT  6.780 0.450 7.060 0.870 ;
        RECT  6.620 2.930 6.900 3.150 ;
        RECT  6.640 1.030 6.740 1.720 ;
        RECT  6.480 1.030 6.640 2.620 ;
        RECT  6.460 1.030 6.480 1.720 ;
        RECT  6.300 2.340 6.480 2.620 ;
        RECT  5.780 1.560 6.460 1.720 ;
        RECT  5.340 1.900 6.320 2.180 ;
        RECT  5.340 0.580 5.540 0.820 ;
        RECT  5.220 2.710 5.500 2.990 ;
        RECT  5.260 0.580 5.340 2.180 ;
        RECT  5.180 0.580 5.260 2.500 ;
        RECT  4.400 2.710 5.220 2.870 ;
        RECT  5.100 1.900 5.180 2.500 ;
        RECT  4.980 2.220 5.100 2.500 ;
        RECT  4.820 0.730 4.940 1.010 ;
        RECT  4.780 0.730 4.820 1.310 ;
        RECT  4.660 0.730 4.780 2.540 ;
        RECT  4.560 1.150 4.660 2.540 ;
        RECT  4.300 1.150 4.560 1.310 ;
        RECT  4.240 1.590 4.400 2.870 ;
        RECT  4.020 1.150 4.300 1.430 ;
        RECT  3.860 1.590 4.240 1.750 ;
        RECT  3.540 1.910 4.080 2.190 ;
        RECT  3.780 0.620 3.860 1.750 ;
        RECT  3.700 0.500 3.780 1.750 ;
        RECT  3.100 0.500 3.700 0.780 ;
        RECT  3.420 0.940 3.540 2.190 ;
        RECT  3.260 0.940 3.420 2.680 ;
        RECT  2.960 2.440 3.260 2.680 ;
        RECT  2.940 0.500 3.100 2.280 ;
        RECT  2.800 2.440 2.960 3.050 ;
        RECT  2.800 0.780 2.940 1.060 ;
        RECT  2.800 1.910 2.940 2.280 ;
        RECT  0.680 2.120 2.800 2.280 ;
        RECT  0.370 2.890 2.800 3.050 ;
        RECT  2.640 1.220 2.780 1.500 ;
        RECT  2.480 0.900 2.640 1.940 ;
        RECT  2.080 0.900 2.480 1.060 ;
        RECT  1.680 1.720 2.480 1.940 ;
        RECT  1.800 0.780 2.080 1.060 ;
        RECT  0.600 2.460 1.920 2.730 ;
        RECT  0.800 0.900 1.800 1.060 ;
        RECT  0.640 0.500 0.800 1.060 ;
        RECT  0.400 1.980 0.680 2.280 ;
        RECT  0.440 0.500 0.640 0.780 ;
        RECT  0.240 0.940 0.480 1.220 ;
        RECT  0.240 2.440 0.370 3.050 ;
        RECT  0.210 0.940 0.240 3.050 ;
        RECT  0.080 0.940 0.210 2.720 ;
    END
END DFFTRX1TR

MACRO DFFSRHQX8TR
    CLASS CORE ;
    FOREIGN DFFSRHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.640 4.960 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.260 1.640 11.520 2.210 ;
        RECT  10.150 1.640 11.260 1.800 ;
        RECT  9.990 1.640 10.150 1.940 ;
        RECT  9.870 1.780 9.990 1.940 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.740 0.470 15.020 3.110 ;
        RECT  14.030 1.440 14.740 2.160 ;
        RECT  13.760 0.470 14.030 3.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.240 3.920 1.600 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.890 1.560 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.500 -0.280 15.600 0.280 ;
        RECT  15.220 -0.280 15.500 1.170 ;
        RECT  14.540 -0.280 15.220 0.280 ;
        RECT  14.260 -0.280 14.540 1.150 ;
        RECT  13.510 -0.280 14.260 0.280 ;
        RECT  13.230 -0.280 13.510 0.610 ;
        RECT  12.010 -0.280 13.230 0.280 ;
        RECT  11.730 -0.280 12.010 0.340 ;
        RECT  8.950 -0.280 11.730 0.280 ;
        RECT  8.670 -0.280 8.950 0.320 ;
        RECT  7.050 -0.280 8.670 0.280 ;
        RECT  6.770 -0.280 7.050 0.340 ;
        RECT  5.020 -0.280 6.770 0.280 ;
        RECT  4.740 -0.280 5.020 0.340 ;
        RECT  2.990 -0.280 4.740 0.280 ;
        RECT  2.710 -0.280 2.990 0.340 ;
        RECT  1.190 -0.280 2.710 0.280 ;
        RECT  0.910 -0.280 1.190 0.340 ;
        RECT  0.000 -0.280 0.910 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.500 3.320 15.600 3.880 ;
        RECT  15.220 2.000 15.500 3.880 ;
        RECT  14.540 3.320 15.220 3.880 ;
        RECT  14.260 2.420 14.540 3.880 ;
        RECT  13.540 3.320 14.260 3.880 ;
        RECT  12.990 2.920 13.540 3.880 ;
        RECT  11.690 3.320 12.990 3.880 ;
        RECT  11.410 3.260 11.690 3.880 ;
        RECT  9.230 3.320 11.410 3.880 ;
        RECT  8.950 3.260 9.230 3.880 ;
        RECT  8.190 3.320 8.950 3.880 ;
        RECT  7.910 3.260 8.190 3.880 ;
        RECT  6.550 3.320 7.910 3.880 ;
        RECT  6.390 2.580 6.550 3.880 ;
        RECT  4.840 3.320 6.390 3.880 ;
        RECT  4.560 3.260 4.840 3.880 ;
        RECT  3.350 3.320 4.560 3.880 ;
        RECT  3.070 3.260 3.350 3.880 ;
        RECT  2.430 3.320 3.070 3.880 ;
        RECT  2.150 3.260 2.430 3.880 ;
        RECT  0.830 3.320 2.150 3.880 ;
        RECT  0.550 3.260 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.300 0.770 13.460 2.540 ;
        RECT  12.590 0.770 13.300 0.930 ;
        RECT  12.800 2.380 13.300 2.540 ;
        RECT  12.930 1.090 13.110 2.220 ;
        RECT  12.830 1.090 12.930 1.730 ;
        RECT  12.630 1.570 12.830 1.730 ;
        RECT  12.640 2.380 12.800 2.850 ;
        RECT  10.780 2.690 12.640 2.850 ;
        RECT  12.430 0.770 12.590 1.050 ;
        RECT  12.280 1.210 12.440 2.530 ;
        RECT  10.190 0.890 12.430 1.050 ;
        RECT  11.100 2.370 12.280 2.530 ;
        RECT  11.860 1.210 12.020 2.210 ;
        RECT  10.030 1.210 11.860 1.370 ;
        RECT  10.940 1.980 11.100 2.530 ;
        RECT  10.830 1.980 10.940 2.260 ;
        RECT  9.710 2.100 10.830 2.260 ;
        RECT  10.620 2.420 10.780 3.160 ;
        RECT  10.030 0.440 10.680 0.600 ;
        RECT  9.810 2.420 10.300 2.700 ;
        RECT  9.550 3.000 10.150 3.160 ;
        RECT  9.870 0.440 10.030 1.370 ;
        RECT  9.270 0.440 9.870 0.600 ;
        RECT  7.950 2.420 9.810 2.580 ;
        RECT  9.550 0.760 9.710 2.260 ;
        RECT  9.430 0.760 9.550 0.960 ;
        RECT  9.110 2.100 9.550 2.260 ;
        RECT  9.390 2.920 9.550 3.160 ;
        RECT  7.630 0.800 9.430 0.960 ;
        RECT  7.950 1.120 9.390 1.280 ;
        RECT  6.930 2.920 9.390 3.080 ;
        RECT  9.110 0.440 9.270 0.640 ;
        RECT  7.370 0.480 9.110 0.640 ;
        RECT  7.790 1.120 7.950 2.580 ;
        RECT  7.770 1.740 7.790 2.020 ;
        RECT  7.470 0.800 7.630 0.980 ;
        RECT  7.470 1.300 7.630 1.580 ;
        RECT  4.460 0.820 7.470 0.980 ;
        RECT  7.350 1.420 7.470 1.580 ;
        RECT  7.210 0.480 7.370 0.660 ;
        RECT  7.190 1.420 7.350 2.690 ;
        RECT  2.970 0.500 7.210 0.660 ;
        RECT  6.260 1.420 7.190 1.580 ;
        RECT  6.770 2.260 6.930 3.080 ;
        RECT  5.980 2.260 6.770 2.420 ;
        RECT  6.100 1.140 6.260 1.580 ;
        RECT  5.280 1.140 6.100 1.300 ;
        RECT  5.820 1.820 5.980 3.160 ;
        RECT  5.600 1.820 5.820 1.980 ;
        RECT  5.160 3.000 5.820 3.160 ;
        RECT  5.440 1.700 5.600 1.980 ;
        RECT  5.480 2.680 5.600 2.840 ;
        RECT  5.280 2.280 5.540 2.440 ;
        RECT  5.320 2.620 5.480 2.840 ;
        RECT  3.810 2.620 5.320 2.780 ;
        RECT  5.120 1.140 5.280 2.440 ;
        RECT  5.000 2.940 5.160 3.160 ;
        RECT  1.570 2.940 5.000 3.100 ;
        RECT  4.240 2.300 4.500 2.460 ;
        RECT  4.240 0.820 4.460 1.250 ;
        RECT  4.080 0.820 4.240 2.460 ;
        RECT  3.650 1.910 3.810 2.780 ;
        RECT  3.290 1.910 3.650 2.070 ;
        RECT  3.290 0.920 3.510 1.080 ;
        RECT  3.130 0.920 3.290 2.070 ;
        RECT  2.810 0.500 2.970 2.740 ;
        RECT  2.190 0.710 2.810 0.870 ;
        RECT  2.730 1.680 2.810 2.740 ;
        RECT  1.710 1.680 2.730 1.840 ;
        RECT  2.030 1.360 2.650 1.520 ;
        RECT  1.870 0.550 2.030 1.520 ;
        RECT  0.610 0.550 1.870 0.710 ;
        RECT  1.390 0.870 1.710 1.030 ;
        RECT  1.550 1.560 1.710 1.840 ;
        RECT  1.410 2.000 1.570 3.100 ;
        RECT  1.390 2.000 1.410 2.160 ;
        RECT  1.230 0.870 1.390 2.160 ;
        RECT  0.310 0.550 0.610 0.870 ;
        RECT  0.150 0.550 0.310 3.000 ;
    END
END DFFSRHQX8TR

MACRO DFFSRHQX4TR
    CLASS CORE ;
    FOREIGN DFFSRHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.640 4.960 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.260 1.640 11.520 2.210 ;
        RECT  10.150 1.640 11.260 1.800 ;
        RECT  9.990 1.640 10.150 1.940 ;
        RECT  9.870 1.780 9.990 1.940 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.180 1.440 14.320 2.160 ;
        RECT  14.170 1.440 14.180 3.160 ;
        RECT  13.820 0.470 14.170 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.240 3.920 1.600 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.890 1.560 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.670 -0.280 14.800 0.280 ;
        RECT  14.400 -0.280 14.670 1.150 ;
        RECT  13.620 -0.280 14.400 0.280 ;
        RECT  13.340 -0.280 13.620 0.340 ;
        RECT  12.160 -0.280 13.340 0.280 ;
        RECT  11.850 -0.280 12.160 0.730 ;
        RECT  8.950 -0.280 11.850 0.280 ;
        RECT  8.670 -0.280 8.950 0.320 ;
        RECT  7.050 -0.280 8.670 0.280 ;
        RECT  6.770 -0.280 7.050 0.340 ;
        RECT  5.020 -0.280 6.770 0.280 ;
        RECT  4.740 -0.280 5.020 0.340 ;
        RECT  2.990 -0.280 4.740 0.280 ;
        RECT  2.710 -0.280 2.990 0.340 ;
        RECT  1.190 -0.280 2.710 0.280 ;
        RECT  0.910 -0.280 1.190 0.340 ;
        RECT  0.000 -0.280 0.910 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.700 3.320 14.800 3.880 ;
        RECT  14.480 1.910 14.700 3.880 ;
        RECT  13.660 3.320 14.480 3.880 ;
        RECT  13.030 2.920 13.660 3.880 ;
        RECT  11.690 3.320 13.030 3.880 ;
        RECT  11.410 3.260 11.690 3.880 ;
        RECT  9.230 3.320 11.410 3.880 ;
        RECT  8.950 3.260 9.230 3.880 ;
        RECT  8.190 3.320 8.950 3.880 ;
        RECT  7.910 3.260 8.190 3.880 ;
        RECT  6.550 3.320 7.910 3.880 ;
        RECT  6.390 2.580 6.550 3.880 ;
        RECT  4.840 3.320 6.390 3.880 ;
        RECT  4.560 3.260 4.840 3.880 ;
        RECT  3.350 3.320 4.560 3.880 ;
        RECT  3.070 3.260 3.350 3.880 ;
        RECT  2.430 3.320 3.070 3.880 ;
        RECT  2.150 3.260 2.430 3.880 ;
        RECT  0.830 3.320 2.150 3.880 ;
        RECT  0.550 3.260 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.530 1.470 13.640 1.750 ;
        RECT  13.370 0.770 13.530 2.540 ;
        RECT  12.690 0.770 13.370 0.930 ;
        RECT  12.800 2.380 13.370 2.540 ;
        RECT  13.050 1.090 13.210 2.220 ;
        RECT  12.930 1.090 13.050 1.250 ;
        RECT  12.660 1.670 13.050 1.830 ;
        RECT  12.640 2.380 12.800 2.850 ;
        RECT  12.530 0.770 12.690 1.050 ;
        RECT  10.780 2.690 12.640 2.850 ;
        RECT  10.190 0.890 12.530 1.050 ;
        RECT  12.480 1.210 12.490 1.490 ;
        RECT  12.320 1.210 12.480 2.530 ;
        RECT  11.100 2.370 12.320 2.530 ;
        RECT  11.920 1.210 12.080 2.210 ;
        RECT  10.030 1.210 11.920 1.370 ;
        RECT  10.940 1.980 11.100 2.530 ;
        RECT  10.830 1.980 10.940 2.260 ;
        RECT  9.710 2.100 10.830 2.260 ;
        RECT  10.620 2.420 10.780 3.160 ;
        RECT  10.030 0.440 10.680 0.600 ;
        RECT  9.810 2.420 10.300 2.700 ;
        RECT  9.550 3.000 10.150 3.160 ;
        RECT  9.870 0.440 10.030 1.370 ;
        RECT  9.270 0.440 9.870 0.600 ;
        RECT  7.950 2.420 9.810 2.580 ;
        RECT  9.550 0.760 9.710 2.260 ;
        RECT  9.430 0.760 9.550 0.960 ;
        RECT  9.110 2.100 9.550 2.260 ;
        RECT  9.390 2.920 9.550 3.160 ;
        RECT  7.630 0.800 9.430 0.960 ;
        RECT  7.950 1.120 9.390 1.280 ;
        RECT  6.930 2.920 9.390 3.080 ;
        RECT  9.110 0.440 9.270 0.640 ;
        RECT  7.370 0.480 9.110 0.640 ;
        RECT  7.790 1.120 7.950 2.580 ;
        RECT  7.770 1.740 7.790 2.020 ;
        RECT  7.470 0.800 7.630 0.980 ;
        RECT  7.470 1.300 7.630 1.580 ;
        RECT  4.460 0.820 7.470 0.980 ;
        RECT  7.350 1.420 7.470 1.580 ;
        RECT  7.210 0.480 7.370 0.660 ;
        RECT  7.190 1.420 7.350 2.690 ;
        RECT  2.970 0.500 7.210 0.660 ;
        RECT  6.260 1.420 7.190 1.580 ;
        RECT  6.770 2.260 6.930 3.080 ;
        RECT  5.980 2.260 6.770 2.420 ;
        RECT  6.100 1.140 6.260 1.580 ;
        RECT  5.280 1.140 6.100 1.300 ;
        RECT  5.820 1.820 5.980 3.160 ;
        RECT  5.600 1.820 5.820 1.980 ;
        RECT  5.160 3.000 5.820 3.160 ;
        RECT  5.440 1.700 5.600 1.980 ;
        RECT  5.480 2.680 5.600 2.840 ;
        RECT  5.280 2.280 5.540 2.440 ;
        RECT  5.320 2.620 5.480 2.840 ;
        RECT  3.810 2.620 5.320 2.780 ;
        RECT  5.120 1.140 5.280 2.440 ;
        RECT  5.000 2.940 5.160 3.160 ;
        RECT  1.570 2.940 5.000 3.100 ;
        RECT  4.240 2.300 4.500 2.460 ;
        RECT  4.240 0.820 4.460 1.250 ;
        RECT  4.080 0.820 4.240 2.460 ;
        RECT  3.650 1.910 3.810 2.780 ;
        RECT  3.290 1.910 3.650 2.070 ;
        RECT  3.290 0.920 3.510 1.080 ;
        RECT  3.130 0.920 3.290 2.070 ;
        RECT  2.810 0.500 2.970 2.740 ;
        RECT  2.190 0.710 2.810 0.870 ;
        RECT  2.730 1.680 2.810 2.740 ;
        RECT  1.710 1.680 2.730 1.840 ;
        RECT  2.030 1.360 2.650 1.520 ;
        RECT  1.870 0.550 2.030 1.520 ;
        RECT  0.610 0.550 1.870 0.710 ;
        RECT  1.390 0.870 1.710 1.030 ;
        RECT  1.550 1.560 1.710 1.840 ;
        RECT  1.410 2.000 1.570 3.100 ;
        RECT  1.390 2.000 1.410 2.160 ;
        RECT  1.230 0.870 1.390 2.160 ;
        RECT  0.310 0.550 0.610 0.870 ;
        RECT  0.150 0.550 0.310 3.000 ;
    END
END DFFSRHQX4TR

MACRO DFFSRHQX2TR
    CLASS CORE ;
    FOREIGN DFFSRHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.220 3.210 1.710 ;
        END
        ANTENNAGATEAREA 0.192 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.760 1.640 9.390 1.870 ;
        RECT  8.440 1.640 8.760 2.120 ;
        RECT  7.720 1.900 8.440 2.120 ;
        END
        ANTENNAGATEAREA 0.216 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.680 0.440 11.920 3.150 ;
        RECT  10.670 2.670 11.680 2.830 ;
        RECT  10.510 2.670 10.670 3.160 ;
        RECT  10.390 2.880 10.510 3.160 ;
        END
        ANTENNADIFFAREA 3.958 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.100 2.400 1.560 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.220 0.760 1.600 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.430 -0.280 12.000 0.280 ;
        RECT  11.150 -0.280 11.430 0.800 ;
        RECT  11.110 -0.280 11.150 0.400 ;
        RECT  9.950 -0.280 11.110 0.280 ;
        RECT  9.670 -0.280 9.950 0.400 ;
        RECT  5.930 -0.280 9.670 0.280 ;
        RECT  5.650 -0.280 5.930 0.340 ;
        RECT  3.730 -0.280 5.650 0.280 ;
        RECT  0.890 -0.280 3.730 0.340 ;
        RECT  0.610 -0.280 0.890 0.360 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.230 3.320 12.000 3.880 ;
        RECT  10.950 2.990 11.230 3.880 ;
        RECT  9.630 3.320 10.950 3.880 ;
        RECT  9.350 3.200 9.630 3.880 ;
        RECT  7.440 3.320 9.350 3.880 ;
        RECT  7.160 3.260 7.440 3.880 ;
        RECT  6.420 3.320 7.160 3.880 ;
        RECT  2.270 3.260 6.420 3.880 ;
        RECT  1.990 3.200 2.270 3.880 ;
        RECT  0.770 3.260 1.990 3.880 ;
        RECT  0.490 2.800 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.150 1.370 11.310 1.590 ;
        RECT  10.990 1.370 11.150 2.510 ;
        RECT  10.830 0.570 10.990 1.590 ;
        RECT  9.630 2.350 10.990 2.510 ;
        RECT  10.510 0.570 10.830 0.730 ;
        RECT  10.630 1.830 10.830 2.110 ;
        RECT  10.630 0.890 10.670 1.230 ;
        RECT  10.350 0.890 10.630 2.110 ;
        RECT  10.230 0.450 10.510 0.730 ;
        RECT  9.750 0.890 10.350 1.050 ;
        RECT  8.750 0.570 10.230 0.730 ;
        RECT  10.030 1.210 10.190 2.190 ;
        RECT  9.910 1.210 10.030 1.430 ;
        RECT  9.080 2.030 10.030 2.190 ;
        RECT  9.710 1.590 9.870 1.870 ;
        RECT  9.470 0.890 9.750 1.110 ;
        RECT  9.550 1.320 9.710 1.870 ;
        RECT  9.400 2.350 9.630 2.570 ;
        RECT  8.840 1.320 9.550 1.480 ;
        RECT  9.240 2.350 9.400 3.020 ;
        RECT  8.790 2.860 9.240 3.020 ;
        RECT  8.920 2.030 9.080 2.700 ;
        RECT  8.710 2.280 8.920 2.700 ;
        RECT  8.310 1.260 8.840 1.480 ;
        RECT  8.510 2.860 8.790 3.140 ;
        RECT  8.470 0.570 8.750 0.930 ;
        RECT  7.560 2.280 8.710 2.440 ;
        RECT  8.150 0.440 8.310 1.480 ;
        RECT  8.080 2.600 8.300 3.160 ;
        RECT  6.250 0.440 8.150 0.600 ;
        RECT  6.990 2.600 8.080 2.760 ;
        RECT  7.830 0.760 7.990 1.740 ;
        RECT  7.640 2.940 7.920 3.160 ;
        RECT  6.410 0.760 7.830 0.980 ;
        RECT  7.560 1.580 7.830 1.740 ;
        RECT  6.990 1.140 7.670 1.420 ;
        RECT  4.810 2.940 7.640 3.100 ;
        RECT  7.400 1.580 7.560 2.440 ;
        RECT  7.280 1.940 7.400 2.440 ;
        RECT  6.830 1.140 6.990 2.760 ;
        RECT  6.110 1.140 6.830 1.420 ;
        RECT  6.660 2.480 6.830 2.760 ;
        RECT  6.550 1.810 6.670 2.090 ;
        RECT  6.230 2.480 6.660 2.640 ;
        RECT  6.390 1.580 6.550 2.090 ;
        RECT  3.530 0.820 6.410 0.980 ;
        RECT  5.790 1.580 6.390 1.740 ;
        RECT  6.090 0.440 6.250 0.660 ;
        RECT  6.070 1.900 6.230 2.640 ;
        RECT  1.860 0.500 6.090 0.660 ;
        RECT  5.950 1.900 6.070 2.120 ;
        RECT  5.630 1.140 5.790 2.780 ;
        RECT  3.850 1.140 5.630 1.420 ;
        RECT  5.310 2.500 5.630 2.780 ;
        RECT  4.810 2.060 5.470 2.340 ;
        RECT  4.650 1.740 4.810 3.100 ;
        RECT  4.290 1.740 4.650 1.900 ;
        RECT  2.590 2.940 4.650 3.100 ;
        RECT  3.850 2.060 4.410 2.340 ;
        RECT  4.010 1.620 4.290 1.900 ;
        RECT  2.750 2.500 4.200 2.780 ;
        RECT  3.690 1.140 3.850 2.340 ;
        RECT  3.370 0.820 3.530 2.240 ;
        RECT  3.050 0.820 3.370 1.060 ;
        RECT  2.750 2.080 3.370 2.240 ;
        RECT  2.720 0.820 2.870 1.040 ;
        RECT  2.570 2.500 2.750 2.660 ;
        RECT  2.570 0.820 2.720 1.910 ;
        RECT  2.430 2.820 2.590 3.100 ;
        RECT  2.560 0.820 2.570 2.660 ;
        RECT  2.410 1.730 2.560 2.660 ;
        RECT  1.690 2.820 2.430 2.980 ;
        RECT  1.860 1.750 2.030 2.320 ;
        RECT  1.750 0.500 1.860 2.320 ;
        RECT  1.700 0.500 1.750 1.960 ;
        RECT  1.640 0.500 1.700 0.930 ;
        RECT  1.250 1.680 1.700 1.960 ;
        RECT  1.530 2.500 1.690 2.980 ;
        RECT  1.410 2.500 1.530 2.780 ;
        RECT  1.190 0.550 1.470 0.780 ;
        RECT  1.090 2.500 1.410 2.660 ;
        RECT  1.090 0.950 1.330 1.110 ;
        RECT  0.310 0.620 1.190 0.780 ;
        RECT  0.930 0.950 1.090 2.660 ;
        RECT  0.150 0.620 0.310 2.200 ;
        RECT  0.090 0.970 0.150 1.250 ;
        RECT  0.090 1.920 0.150 2.200 ;
    END
END DFFSRHQX2TR

MACRO DFFSRHQX1TR
    CLASS CORE ;
    FOREIGN DFFSRHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.240 3.200 1.800 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.840 1.640 9.120 1.980 ;
        RECT  8.400 1.800 8.840 1.960 ;
        RECT  8.120 1.700 8.400 1.980 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.240 0.840 11.600 2.650 ;
        END
        ANTENNADIFFAREA 1.952 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.200 2.400 1.640 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.890 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.080 -0.280 12.000 0.280 ;
        RECT  10.800 -0.280 11.080 0.400 ;
        RECT  9.760 -0.280 10.800 0.280 ;
        RECT  9.480 -0.280 9.760 0.360 ;
        RECT  0.930 -0.280 9.480 0.280 ;
        RECT  0.650 -0.280 0.930 0.400 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.040 3.320 12.000 3.880 ;
        RECT  10.360 3.040 11.040 3.880 ;
        RECT  9.440 3.320 10.360 3.880 ;
        RECT  9.160 3.200 9.440 3.880 ;
        RECT  7.320 3.320 9.160 3.880 ;
        RECT  7.040 3.260 7.320 3.880 ;
        RECT  6.340 3.320 7.040 3.880 ;
        RECT  5.080 3.260 6.340 3.880 ;
        RECT  3.850 3.320 5.080 3.880 ;
        RECT  3.570 3.200 3.850 3.880 ;
        RECT  2.390 3.320 3.570 3.880 ;
        RECT  2.110 3.200 2.390 3.880 ;
        RECT  0.810 3.260 2.110 3.880 ;
        RECT  0.530 2.800 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.960 1.310 11.080 1.590 ;
        RECT  10.800 0.560 10.960 2.760 ;
        RECT  10.320 0.560 10.800 0.720 ;
        RECT  9.120 2.480 10.800 2.760 ;
        RECT  10.520 1.910 10.640 2.190 ;
        RECT  10.360 1.030 10.520 2.190 ;
        RECT  10.240 1.030 10.360 1.310 ;
        RECT  10.160 1.470 10.360 1.750 ;
        RECT  10.040 0.440 10.320 0.720 ;
        RECT  9.880 0.880 10.080 1.160 ;
        RECT  8.720 0.520 10.040 0.720 ;
        RECT  9.880 1.810 10.000 2.090 ;
        RECT  9.720 0.880 9.880 2.320 ;
        RECT  8.800 2.160 9.720 2.320 ;
        RECT  9.440 1.720 9.560 2.000 ;
        RECT  9.280 0.960 9.440 2.000 ;
        RECT  8.280 0.960 9.280 1.120 ;
        RECT  8.960 2.480 9.120 3.040 ;
        RECT  8.570 2.880 8.960 3.040 ;
        RECT  8.520 2.160 8.800 2.720 ;
        RECT  8.440 0.520 8.720 0.800 ;
        RECT  8.290 2.880 8.570 3.150 ;
        RECT  7.960 2.160 8.520 2.320 ;
        RECT  8.120 0.440 8.280 1.120 ;
        RECT  1.820 0.440 8.120 0.600 ;
        RECT  6.980 2.500 8.090 2.780 ;
        RECT  7.800 0.760 7.960 2.320 ;
        RECT  3.520 0.760 7.800 0.920 ;
        RECT  7.440 2.160 7.800 2.320 ;
        RECT  7.640 3.000 7.760 3.160 ;
        RECT  6.980 1.090 7.640 1.310 ;
        RECT  7.480 2.940 7.640 3.160 ;
        RECT  4.920 2.940 7.480 3.100 ;
        RECT  7.160 1.940 7.440 2.320 ;
        RECT  6.820 1.090 6.980 2.780 ;
        RECT  5.940 1.090 6.820 1.310 ;
        RECT  6.220 2.500 6.820 2.780 ;
        RECT  6.540 2.020 6.660 2.300 ;
        RECT  6.380 1.590 6.540 2.300 ;
        RECT  5.780 1.590 6.380 1.750 ;
        RECT  5.940 2.020 6.220 2.780 ;
        RECT  5.620 1.590 5.780 2.630 ;
        RECT  5.240 1.590 5.620 1.750 ;
        RECT  5.300 2.350 5.620 2.630 ;
        RECT  4.920 1.910 5.460 2.190 ;
        RECT  5.080 1.080 5.240 1.750 ;
        RECT  3.840 1.080 5.080 1.300 ;
        RECT  4.760 1.460 4.920 3.100 ;
        RECT  4.000 1.460 4.760 1.680 ;
        RECT  4.170 2.940 4.760 3.100 ;
        RECT  4.380 2.500 4.600 2.780 ;
        RECT  3.840 1.910 4.400 2.190 ;
        RECT  3.090 2.500 4.380 2.660 ;
        RECT  4.010 2.880 4.170 3.100 ;
        RECT  3.410 2.880 4.010 3.040 ;
        RECT  3.680 1.080 3.840 2.190 ;
        RECT  3.360 0.760 3.520 2.340 ;
        RECT  3.250 2.880 3.410 3.130 ;
        RECT  3.000 0.760 3.360 1.040 ;
        RECT  3.000 2.060 3.360 2.340 ;
        RECT  2.710 2.970 3.250 3.130 ;
        RECT  2.870 2.500 3.090 2.810 ;
        RECT  2.720 2.500 2.870 2.660 ;
        RECT  2.720 0.760 2.820 1.040 ;
        RECT  2.560 0.760 2.720 2.660 ;
        RECT  2.550 2.820 2.710 3.130 ;
        RECT  1.730 2.820 2.550 2.980 ;
        RECT  1.910 2.120 2.190 2.450 ;
        RECT  1.820 2.120 1.910 2.280 ;
        RECT  1.660 0.440 1.820 2.280 ;
        RECT  1.570 2.440 1.730 2.980 ;
        RECT  1.540 0.440 1.660 0.940 ;
        RECT  1.250 1.740 1.660 2.020 ;
        RECT  1.450 2.440 1.570 2.720 ;
        RECT  1.090 2.440 1.450 2.600 ;
        RECT  1.100 0.440 1.380 0.720 ;
        RECT  1.090 1.030 1.370 1.310 ;
        RECT  0.310 0.560 1.100 0.720 ;
        RECT  0.930 1.030 1.090 2.600 ;
        RECT  0.150 0.560 0.310 2.300 ;
        RECT  0.090 1.030 0.150 1.310 ;
        RECT  0.090 2.020 0.150 2.300 ;
    END
END DFFSRHQX1TR

MACRO DFFSRXLTR
    CLASS CORE ;
    FOREIGN DFFSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 2.780 7.560 3.160 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.580 3.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.370 2.040 9.520 2.670 ;
        RECT  9.210 0.620 9.370 2.670 ;
        RECT  8.750 0.620 9.210 0.780 ;
        RECT  8.750 2.510 9.210 2.670 ;
        END
        ANTENNADIFFAREA 1.0895 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.200 1.240 10.320 2.360 ;
        RECT  10.160 1.030 10.200 2.360 ;
        RECT  10.000 1.030 10.160 2.370 ;
        RECT  9.920 1.030 10.000 1.310 ;
        END
        ANTENNADIFFAREA 1.199 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.930 0.360 2.370 ;
        RECT  0.080 1.240 0.320 2.370 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.410 2.760 1.690 ;
        RECT  2.040 1.240 2.360 1.690 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.630 -0.280 10.400 0.280 ;
        RECT  9.330 -0.280 9.630 0.360 ;
        RECT  8.410 -0.280 9.330 0.280 ;
        RECT  7.710 -0.280 8.410 0.800 ;
        RECT  3.480 -0.280 7.710 0.280 ;
        RECT  3.200 -0.280 3.480 0.290 ;
        RECT  2.140 -0.280 3.200 0.280 ;
        RECT  1.860 -0.280 2.140 0.290 ;
        RECT  0.370 -0.280 1.860 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.320 10.400 3.880 ;
        RECT  9.290 3.250 9.580 3.880 ;
        RECT  8.470 3.320 9.290 3.880 ;
        RECT  8.190 3.260 8.470 3.880 ;
        RECT  6.340 3.320 8.190 3.880 ;
        RECT  5.620 3.260 6.340 3.880 ;
        RECT  4.290 3.320 5.620 3.880 ;
        RECT  3.490 2.880 4.290 3.880 ;
        RECT  2.020 3.320 3.490 3.880 ;
        RECT  1.740 3.260 2.020 3.880 ;
        RECT  0.360 3.320 1.740 3.880 ;
        RECT  0.130 2.610 0.360 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.680 1.550 9.840 3.060 ;
        RECT  9.530 1.550 9.680 1.840 ;
        RECT  8.420 2.900 9.680 3.060 ;
        RECT  8.980 1.480 9.050 1.780 ;
        RECT  8.820 1.060 8.980 2.220 ;
        RECT  8.710 1.060 8.820 1.340 ;
        RECT  8.690 2.000 8.820 2.220 ;
        RECT  8.420 1.520 8.650 1.800 ;
        RECT  8.260 1.150 8.420 3.060 ;
        RECT  8.030 1.150 8.260 1.310 ;
        RECT  7.960 1.940 8.260 2.100 ;
        RECT  7.880 1.470 8.100 1.750 ;
        RECT  7.750 1.030 8.030 1.310 ;
        RECT  7.720 1.940 7.960 2.220 ;
        RECT  7.510 1.470 7.880 1.630 ;
        RECT  7.680 1.800 7.720 2.220 ;
        RECT  7.560 1.800 7.680 2.100 ;
        RECT  7.190 1.800 7.560 1.960 ;
        RECT  7.230 0.440 7.510 0.720 ;
        RECT  7.350 1.360 7.510 1.630 ;
        RECT  7.120 2.120 7.400 2.400 ;
        RECT  6.430 1.360 7.350 1.520 ;
        RECT  5.060 0.440 7.230 0.600 ;
        RECT  6.910 1.680 7.190 1.960 ;
        RECT  6.920 2.240 7.120 2.400 ;
        RECT  6.760 2.240 6.920 3.100 ;
        RECT  6.590 0.770 6.870 1.000 ;
        RECT  4.620 2.880 6.760 3.100 ;
        RECT  6.600 1.680 6.720 1.960 ;
        RECT  6.440 1.680 6.600 2.720 ;
        RECT  5.900 0.770 6.590 0.930 ;
        RECT  2.580 2.560 6.440 2.720 ;
        RECT  6.280 1.090 6.430 1.520 ;
        RECT  6.060 1.090 6.280 2.290 ;
        RECT  5.740 0.770 5.900 2.400 ;
        RECT  5.420 1.480 5.740 1.760 ;
        RECT  4.900 2.240 5.740 2.400 ;
        RECT  5.300 0.950 5.580 1.320 ;
        RECT  5.260 1.920 5.460 2.080 ;
        RECT  5.260 1.160 5.300 1.320 ;
        RECT  5.100 1.160 5.260 2.080 ;
        RECT  4.680 1.160 5.100 1.320 ;
        RECT  4.840 0.440 5.060 1.000 ;
        RECT  4.740 1.480 4.900 2.400 ;
        RECT  4.360 1.480 4.740 1.640 ;
        RECT  4.520 0.450 4.680 1.320 ;
        RECT  4.040 1.800 4.580 2.080 ;
        RECT  1.810 0.450 4.520 0.610 ;
        RECT  4.200 0.770 4.360 1.640 ;
        RECT  3.080 0.770 4.200 0.930 ;
        RECT  3.880 1.090 4.040 2.400 ;
        RECT  3.760 1.090 3.880 1.310 ;
        RECT  3.760 2.120 3.880 2.400 ;
        RECT  2.990 2.940 3.270 3.160 ;
        RECT  3.040 0.770 3.080 2.010 ;
        RECT  2.920 0.770 3.040 2.270 ;
        RECT  1.260 2.940 2.990 3.100 ;
        RECT  2.760 0.970 2.920 1.250 ;
        RECT  2.760 1.850 2.920 2.270 ;
        RECT  1.280 1.850 2.760 2.130 ;
        RECT  2.210 0.800 2.580 1.080 ;
        RECT  1.580 2.560 2.580 2.780 ;
        RECT  1.490 0.920 2.210 1.080 ;
        RECT  1.530 0.450 1.810 0.760 ;
        RECT  1.420 2.290 1.580 2.780 ;
        RECT  1.330 0.920 1.490 1.690 ;
        RECT  1.120 2.290 1.420 2.450 ;
        RECT  1.130 1.410 1.330 1.690 ;
        RECT  1.100 2.610 1.260 3.100 ;
        RECT  0.890 0.970 1.170 1.250 ;
        RECT  1.120 1.530 1.130 1.690 ;
        RECT  0.960 1.530 1.120 2.450 ;
        RECT  0.680 2.610 1.100 2.890 ;
        RECT  0.840 2.170 0.960 2.450 ;
        RECT  0.680 1.090 0.890 1.250 ;
        RECT  0.520 1.090 0.680 2.890 ;
    END
END DFFSRXLTR

MACRO DFFSRX4TR
    CLASS CORE ;
    FOREIGN DFFSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.880 2.440 7.120 2.870 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.580 3.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.010 0.630 10.320 3.160 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.970 1.090 9.250 2.380 ;
        RECT  8.880 1.440 8.970 2.380 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.490 2.800 1.650 ;
        RECT  2.080 1.240 2.320 1.650 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 -0.280 10.800 0.280 ;
        RECT  10.480 -0.280 10.710 1.270 ;
        RECT  9.750 -0.280 10.480 0.280 ;
        RECT  9.470 -0.280 9.750 0.610 ;
        RECT  8.770 -0.280 9.470 0.280 ;
        RECT  8.490 -0.280 8.770 0.610 ;
        RECT  7.730 -0.280 8.490 0.280 ;
        RECT  7.450 -0.280 7.730 0.400 ;
        RECT  4.060 -0.280 7.450 0.280 ;
        RECT  2.970 -0.280 4.060 0.370 ;
        RECT  1.260 -0.280 2.970 0.280 ;
        RECT  1.040 -0.280 1.260 0.730 ;
        RECT  0.440 -0.280 1.040 0.280 ;
        RECT  0.090 -0.280 0.440 0.840 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 3.320 10.800 3.880 ;
        RECT  10.480 2.100 10.710 3.880 ;
        RECT  9.750 3.320 10.480 3.880 ;
        RECT  9.470 2.970 9.750 3.880 ;
        RECT  8.770 3.320 9.470 3.880 ;
        RECT  8.490 2.970 8.770 3.880 ;
        RECT  7.630 3.320 8.490 3.880 ;
        RECT  7.350 3.200 7.630 3.880 ;
        RECT  6.180 3.320 7.350 3.880 ;
        RECT  5.460 3.260 6.180 3.880 ;
        RECT  4.140 3.320 5.460 3.880 ;
        RECT  3.210 3.000 4.140 3.880 ;
        RECT  1.930 3.320 3.210 3.880 ;
        RECT  1.710 2.830 1.930 3.880 ;
        RECT  0.370 3.320 1.710 3.880 ;
        RECT  0.090 3.260 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.790 1.430 9.850 1.710 ;
        RECT  9.630 0.770 9.790 2.710 ;
        RECT  8.290 0.770 9.630 0.930 ;
        RECT  8.250 2.550 9.630 2.710 ;
        RECT  8.190 1.580 8.430 1.860 ;
        RECT  8.010 0.530 8.290 0.930 ;
        RECT  7.970 2.550 8.250 3.150 ;
        RECT  8.030 1.110 8.190 2.190 ;
        RECT  7.750 2.030 8.030 2.310 ;
        RECT  7.690 1.300 7.850 1.860 ;
        RECT  7.530 2.030 7.750 2.190 ;
        RECT  6.140 1.300 7.690 1.460 ;
        RECT  7.370 1.700 7.530 2.190 ;
        RECT  6.990 1.700 7.370 1.860 ;
        RECT  7.090 0.440 7.250 1.130 ;
        RECT  4.800 0.440 7.090 0.600 ;
        RECT  6.720 2.020 7.070 2.180 ;
        RECT  6.710 1.620 6.990 1.860 ;
        RECT  6.560 2.020 6.720 3.100 ;
        RECT  6.390 0.760 6.670 1.140 ;
        RECT  4.500 2.940 6.560 3.100 ;
        RECT  5.600 0.760 6.390 0.920 ;
        RECT  6.280 1.640 6.380 1.860 ;
        RECT  6.120 1.640 6.280 2.780 ;
        RECT  5.960 1.080 6.140 1.460 ;
        RECT  2.570 2.620 6.120 2.780 ;
        RECT  5.860 1.080 5.960 2.200 ;
        RECT  5.800 1.300 5.860 2.200 ;
        RECT  5.600 1.610 5.640 2.460 ;
        RECT  5.480 0.760 5.600 2.460 ;
        RECT  5.440 0.760 5.480 1.770 ;
        RECT  4.700 2.300 5.480 2.460 ;
        RECT  5.220 1.610 5.440 1.770 ;
        RECT  5.060 1.980 5.300 2.140 ;
        RECT  5.120 0.900 5.280 1.450 ;
        RECT  5.060 1.290 5.120 1.450 ;
        RECT  4.900 1.290 5.060 2.140 ;
        RECT  4.480 1.290 4.900 1.450 ;
        RECT  4.640 0.440 4.800 1.130 ;
        RECT  4.540 1.680 4.700 2.460 ;
        RECT  4.160 1.680 4.540 1.840 ;
        RECT  4.320 0.530 4.480 1.450 ;
        RECT  3.920 2.000 4.380 2.160 ;
        RECT  2.960 0.530 4.320 0.690 ;
        RECT  4.000 0.850 4.160 1.840 ;
        RECT  3.280 0.850 4.000 1.010 ;
        RECT  3.840 2.000 3.920 2.340 ;
        RECT  3.680 1.170 3.840 2.340 ;
        RECT  3.530 1.170 3.680 1.330 ;
        RECT  3.640 2.120 3.680 2.340 ;
        RECT  3.120 0.850 3.280 1.250 ;
        RECT  2.960 1.090 3.120 2.270 ;
        RECT  2.250 3.000 3.050 3.160 ;
        RECT  2.800 0.530 2.960 0.930 ;
        RECT  2.480 1.090 2.960 1.250 ;
        RECT  2.730 1.810 2.960 2.270 ;
        RECT  1.900 0.770 2.800 0.930 ;
        RECT  2.060 1.810 2.730 1.970 ;
        RECT  1.580 0.450 2.640 0.610 ;
        RECT  2.410 2.190 2.570 2.820 ;
        RECT  1.320 2.190 2.410 2.350 ;
        RECT  2.090 2.510 2.250 3.160 ;
        RECT  1.150 2.510 2.090 2.670 ;
        RECT  1.740 0.770 1.900 2.030 ;
        RECT  1.480 1.870 1.740 2.030 ;
        RECT  1.420 0.450 1.580 1.630 ;
        RECT  1.320 1.470 1.420 1.630 ;
        RECT  1.160 1.470 1.320 2.350 ;
        RECT  1.000 0.960 1.260 1.240 ;
        RECT  1.000 2.510 1.150 2.780 ;
        RECT  0.840 0.960 1.000 2.780 ;
    END
END DFFSRX4TR

MACRO DFFSRX2TR
    CLASS CORE ;
    FOREIGN DFFSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 2.760 7.560 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.640 3.700 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.440 1.640 9.520 1.960 ;
        RECT  9.420 1.630 9.440 2.660 ;
        RECT  9.280 0.500 9.420 2.660 ;
        RECT  9.260 0.500 9.280 1.960 ;
        RECT  8.890 2.500 9.280 2.660 ;
        RECT  9.000 0.500 9.260 0.660 ;
        END
        ANTENNADIFFAREA 2.928 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.220 1.240 10.320 2.360 ;
        RECT  10.180 0.490 10.220 2.360 ;
        RECT  10.020 0.490 10.180 3.100 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.360 2.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.410 2.760 1.690 ;
        RECT  2.200 1.240 2.360 1.690 ;
        RECT  2.040 1.240 2.200 1.560 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.760 -0.280 10.400 0.280 ;
        RECT  9.580 -0.280 9.760 1.140 ;
        RECT  8.570 -0.280 9.580 0.280 ;
        RECT  8.260 -0.280 8.570 0.560 ;
        RECT  7.980 -0.280 8.260 0.280 ;
        RECT  7.680 -0.280 7.980 0.700 ;
        RECT  3.460 -0.280 7.680 0.280 ;
        RECT  3.180 -0.280 3.460 0.290 ;
        RECT  2.100 -0.280 3.180 0.280 ;
        RECT  1.820 -0.280 2.100 0.290 ;
        RECT  0.370 -0.280 1.820 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.720 3.320 10.400 3.880 ;
        RECT  9.440 3.170 9.720 3.880 ;
        RECT  8.660 3.320 9.440 3.880 ;
        RECT  8.090 3.260 8.660 3.880 ;
        RECT  7.930 2.530 8.090 3.880 ;
        RECT  6.430 3.320 7.930 3.880 ;
        RECT  5.680 3.260 6.430 3.880 ;
        RECT  4.320 3.320 5.680 3.880 ;
        RECT  3.410 2.940 4.320 3.880 ;
        RECT  2.080 3.320 3.410 3.880 ;
        RECT  1.800 3.260 2.080 3.880 ;
        RECT  0.480 3.320 1.800 3.880 ;
        RECT  0.200 3.260 0.480 3.880 ;
        RECT  0.000 3.320 0.200 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.700 1.350 9.860 2.980 ;
        RECT  8.420 2.820 9.700 2.980 ;
        RECT  9.010 1.370 9.100 1.640 ;
        RECT  8.960 0.950 9.010 1.640 ;
        RECT  8.800 0.950 8.960 2.180 ;
        RECT  8.700 0.950 8.800 1.210 ;
        RECT  8.580 1.910 8.800 2.180 ;
        RECT  8.420 1.450 8.640 1.730 ;
        RECT  8.260 1.020 8.420 2.980 ;
        RECT  7.740 1.020 8.260 1.180 ;
        RECT  7.890 1.780 8.260 1.950 ;
        RECT  7.850 1.340 8.100 1.590 ;
        RECT  7.640 1.780 7.890 2.190 ;
        RECT  6.370 1.340 7.850 1.500 ;
        RECT  7.170 1.780 7.640 1.940 ;
        RECT  5.040 0.440 7.500 0.600 ;
        RECT  7.060 2.100 7.340 2.380 ;
        RECT  6.890 1.660 7.170 1.940 ;
        RECT  6.900 2.220 7.060 2.380 ;
        RECT  6.740 2.220 6.900 3.100 ;
        RECT  6.720 0.940 6.840 1.180 ;
        RECT  4.600 2.940 6.740 3.100 ;
        RECT  6.560 0.760 6.720 1.180 ;
        RECT  6.580 1.660 6.700 1.940 ;
        RECT  6.420 1.660 6.580 2.720 ;
        RECT  5.820 0.760 6.560 0.920 ;
        RECT  2.640 2.560 6.420 2.720 ;
        RECT  6.260 1.080 6.370 1.500 ;
        RECT  6.090 1.080 6.260 2.270 ;
        RECT  5.980 1.970 6.090 2.270 ;
        RECT  5.660 0.760 5.820 2.400 ;
        RECT  5.400 1.480 5.660 1.700 ;
        RECT  4.880 2.240 5.660 2.400 ;
        RECT  5.280 0.940 5.500 1.320 ;
        RECT  5.240 1.860 5.440 2.080 ;
        RECT  5.240 1.160 5.280 1.320 ;
        RECT  5.080 1.160 5.240 2.080 ;
        RECT  4.660 1.160 5.080 1.320 ;
        RECT  4.820 0.440 5.040 1.000 ;
        RECT  4.720 1.480 4.880 2.400 ;
        RECT  4.340 1.480 4.720 1.640 ;
        RECT  4.500 0.450 4.660 1.320 ;
        RECT  4.020 1.800 4.560 2.080 ;
        RECT  1.490 0.450 4.500 0.610 ;
        RECT  4.180 0.770 4.340 1.640 ;
        RECT  3.080 0.770 4.180 0.930 ;
        RECT  3.860 1.090 4.020 2.400 ;
        RECT  3.740 1.090 3.860 1.310 ;
        RECT  3.740 2.120 3.860 2.400 ;
        RECT  2.970 2.940 3.250 3.160 ;
        RECT  3.020 0.770 3.080 2.010 ;
        RECT  2.920 0.770 3.020 2.260 ;
        RECT  1.320 2.940 2.970 3.100 ;
        RECT  2.740 1.030 2.920 1.250 ;
        RECT  2.740 1.850 2.920 2.260 ;
        RECT  1.280 1.850 2.740 2.130 ;
        RECT  1.640 2.560 2.640 2.780 ;
        RECT  1.450 0.770 2.540 0.990 ;
        RECT  1.480 2.290 1.640 2.780 ;
        RECT  1.120 2.290 1.480 2.450 ;
        RECT  1.290 0.770 1.450 1.430 ;
        RECT  1.160 2.610 1.320 3.100 ;
        RECT  1.120 1.150 1.290 1.430 ;
        RECT  0.680 2.610 1.160 2.890 ;
        RECT  0.850 0.710 1.130 0.990 ;
        RECT  1.090 1.150 1.120 2.450 ;
        RECT  0.960 1.270 1.090 2.450 ;
        RECT  0.840 2.170 0.960 2.450 ;
        RECT  0.680 0.830 0.850 0.990 ;
        RECT  0.520 0.830 0.680 2.890 ;
    END
END DFFSRX2TR

MACRO DFFSRX1TR
    CLASS CORE ;
    FOREIGN DFFSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 2.780 7.560 3.160 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.580 3.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.370 2.040 9.520 2.730 ;
        RECT  9.210 0.620 9.370 2.730 ;
        RECT  8.750 0.620 9.210 0.780 ;
        RECT  8.750 2.570 9.210 2.730 ;
        END
        ANTENNADIFFAREA 1.875 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.160 1.240 10.320 2.360 ;
        RECT  10.000 1.030 10.160 2.450 ;
        RECT  9.880 1.030 10.000 1.310 ;
        END
        ANTENNADIFFAREA 2.204 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.930 0.360 2.370 ;
        RECT  0.080 1.240 0.320 2.370 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.410 2.760 1.690 ;
        RECT  2.040 1.240 2.360 1.690 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.620 -0.280 10.400 0.280 ;
        RECT  9.290 -0.280 9.620 0.360 ;
        RECT  8.410 -0.280 9.290 0.280 ;
        RECT  7.710 -0.280 8.410 0.800 ;
        RECT  3.480 -0.280 7.710 0.280 ;
        RECT  3.200 -0.280 3.480 0.290 ;
        RECT  2.140 -0.280 3.200 0.280 ;
        RECT  1.860 -0.280 2.140 0.290 ;
        RECT  0.370 -0.280 1.860 0.280 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.580 3.320 10.400 3.880 ;
        RECT  9.290 3.250 9.580 3.880 ;
        RECT  8.470 3.320 9.290 3.880 ;
        RECT  8.190 3.260 8.470 3.880 ;
        RECT  6.430 3.320 8.190 3.880 ;
        RECT  5.620 3.260 6.430 3.880 ;
        RECT  4.290 3.320 5.620 3.880 ;
        RECT  3.490 2.880 4.290 3.880 ;
        RECT  2.020 3.320 3.490 3.880 ;
        RECT  1.740 3.260 2.020 3.880 ;
        RECT  0.360 3.320 1.740 3.880 ;
        RECT  0.130 2.610 0.360 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.680 1.550 9.840 3.060 ;
        RECT  9.530 1.550 9.680 1.840 ;
        RECT  8.420 2.900 9.680 3.060 ;
        RECT  8.980 1.480 9.050 1.780 ;
        RECT  8.820 1.060 8.980 2.220 ;
        RECT  8.710 1.060 8.820 1.340 ;
        RECT  8.690 2.000 8.820 2.220 ;
        RECT  8.420 1.520 8.650 1.800 ;
        RECT  8.260 1.150 8.420 3.060 ;
        RECT  8.030 1.150 8.260 1.310 ;
        RECT  7.960 1.940 8.260 2.100 ;
        RECT  7.880 1.470 8.100 1.750 ;
        RECT  7.750 1.030 8.030 1.310 ;
        RECT  7.720 1.940 7.960 2.220 ;
        RECT  7.510 1.470 7.880 1.630 ;
        RECT  7.680 1.800 7.720 2.220 ;
        RECT  7.560 1.800 7.680 2.100 ;
        RECT  7.190 1.800 7.560 1.960 ;
        RECT  7.230 0.440 7.510 0.720 ;
        RECT  7.350 1.360 7.510 1.630 ;
        RECT  7.120 2.120 7.400 2.400 ;
        RECT  6.430 1.360 7.350 1.520 ;
        RECT  5.060 0.440 7.230 0.600 ;
        RECT  6.910 1.680 7.190 1.960 ;
        RECT  6.920 2.240 7.120 2.400 ;
        RECT  6.760 2.240 6.920 3.100 ;
        RECT  6.590 0.770 6.870 1.000 ;
        RECT  4.620 2.880 6.760 3.100 ;
        RECT  6.600 1.680 6.720 1.960 ;
        RECT  6.440 1.680 6.600 2.720 ;
        RECT  5.900 0.770 6.590 0.930 ;
        RECT  2.580 2.560 6.440 2.720 ;
        RECT  6.280 1.090 6.430 1.520 ;
        RECT  6.060 1.090 6.280 2.290 ;
        RECT  5.740 0.770 5.900 2.400 ;
        RECT  5.420 1.480 5.740 1.760 ;
        RECT  4.900 2.240 5.740 2.400 ;
        RECT  5.300 0.950 5.580 1.320 ;
        RECT  5.260 1.920 5.460 2.080 ;
        RECT  5.260 1.160 5.300 1.320 ;
        RECT  5.100 1.160 5.260 2.080 ;
        RECT  4.680 1.160 5.100 1.320 ;
        RECT  4.840 0.440 5.060 1.000 ;
        RECT  4.740 1.480 4.900 2.400 ;
        RECT  4.360 1.480 4.740 1.640 ;
        RECT  4.520 0.450 4.680 1.320 ;
        RECT  4.040 1.800 4.580 2.080 ;
        RECT  1.810 0.450 4.520 0.610 ;
        RECT  4.200 0.770 4.360 1.640 ;
        RECT  3.080 0.770 4.200 0.930 ;
        RECT  3.880 1.090 4.040 2.400 ;
        RECT  3.760 1.090 3.880 1.310 ;
        RECT  3.760 2.120 3.880 2.400 ;
        RECT  2.990 2.940 3.270 3.160 ;
        RECT  3.040 0.770 3.080 2.010 ;
        RECT  2.920 0.770 3.040 2.270 ;
        RECT  1.260 2.940 2.990 3.100 ;
        RECT  2.760 0.970 2.920 1.250 ;
        RECT  2.760 1.850 2.920 2.270 ;
        RECT  1.280 1.850 2.760 2.130 ;
        RECT  2.210 0.800 2.580 1.080 ;
        RECT  1.580 2.560 2.580 2.780 ;
        RECT  1.490 0.920 2.210 1.080 ;
        RECT  1.530 0.450 1.810 0.760 ;
        RECT  1.420 2.290 1.580 2.780 ;
        RECT  1.330 0.920 1.490 1.690 ;
        RECT  1.120 2.290 1.420 2.450 ;
        RECT  1.130 1.410 1.330 1.690 ;
        RECT  1.100 2.610 1.260 3.100 ;
        RECT  0.890 0.970 1.170 1.250 ;
        RECT  1.120 1.530 1.130 1.690 ;
        RECT  0.960 1.530 1.120 2.450 ;
        RECT  0.680 2.610 1.100 2.890 ;
        RECT  0.840 2.170 0.960 2.450 ;
        RECT  0.680 1.090 0.890 1.250 ;
        RECT  0.520 1.090 0.680 2.890 ;
    END
END DFFSRX1TR

MACRO DFFSHQX8TR
    CLASS CORE ;
    FOREIGN DFFSHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.340 1.640 6.720 2.080 ;
        END
        ANTENNAGATEAREA 0.3264 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.710 0.440 14.970 3.160 ;
        RECT  14.700 1.440 14.710 3.160 ;
        RECT  14.100 1.440 14.700 2.160 ;
        RECT  14.090 1.440 14.100 3.160 ;
        RECT  13.830 0.440 14.090 3.160 ;
        END
        ANTENNADIFFAREA 7.944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.580 3.330 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.510 1.670 1.960 ;
        RECT  0.850 1.510 1.240 1.790 ;
        END
        ANTENNAGATEAREA 0.4128 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.500 -0.280 15.600 0.280 ;
        RECT  15.220 -0.280 15.500 1.260 ;
        RECT  14.540 -0.280 15.220 0.280 ;
        RECT  14.260 -0.280 14.540 1.060 ;
        RECT  13.540 -0.280 14.260 0.280 ;
        RECT  13.260 -0.280 13.540 0.300 ;
        RECT  11.510 -0.280 13.260 0.280 ;
        RECT  11.510 1.180 12.070 1.460 ;
        RECT  11.230 -0.280 11.510 1.460 ;
        RECT  8.640 -0.280 11.230 0.280 ;
        RECT  8.360 -0.280 8.640 0.580 ;
        RECT  7.720 -0.280 8.360 0.280 ;
        RECT  7.440 -0.280 7.720 0.580 ;
        RECT  6.380 -0.280 7.440 0.280 ;
        RECT  6.100 -0.280 6.380 0.580 ;
        RECT  3.900 -0.280 6.100 0.280 ;
        RECT  3.620 -0.280 3.900 0.300 ;
        RECT  2.180 -0.280 3.620 0.280 ;
        RECT  2.020 -0.280 2.180 0.720 ;
        RECT  0.890 -0.280 2.020 0.340 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.450 3.320 15.600 3.880 ;
        RECT  15.220 1.880 15.450 3.880 ;
        RECT  14.540 3.320 15.220 3.880 ;
        RECT  14.260 2.350 14.540 3.880 ;
        RECT  13.440 3.320 14.260 3.880 ;
        RECT  13.160 3.200 13.440 3.880 ;
        RECT  11.070 3.320 13.160 3.880 ;
        RECT  10.790 3.200 11.070 3.880 ;
        RECT  8.540 3.320 10.790 3.880 ;
        RECT  8.260 2.960 8.540 3.880 ;
        RECT  6.620 3.260 8.260 3.880 ;
        RECT  6.000 3.320 6.620 3.880 ;
        RECT  5.720 3.260 6.000 3.880 ;
        RECT  4.210 3.320 5.720 3.880 ;
        RECT  3.930 3.200 4.210 3.880 ;
        RECT  3.170 3.320 3.930 3.880 ;
        RECT  2.890 3.200 3.170 3.880 ;
        RECT  1.150 3.320 2.890 3.880 ;
        RECT  0.870 3.200 1.150 3.880 ;
        RECT  0.260 3.260 0.870 3.880 ;
        RECT  0.000 3.320 0.260 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.510 0.460 13.670 3.040 ;
        RECT  11.790 0.460 13.510 0.620 ;
        RECT  12.350 2.880 13.510 3.040 ;
        RECT  13.160 1.710 13.320 2.720 ;
        RECT  13.060 1.710 13.160 1.970 ;
        RECT  10.730 2.560 13.160 2.720 ;
        RECT  12.900 0.780 13.060 1.970 ;
        RECT  12.570 2.240 12.980 2.400 ;
        RECT  12.740 0.780 12.900 0.940 ;
        RECT  12.410 1.180 12.570 2.400 ;
        RECT  11.430 1.840 12.410 2.000 ;
        RECT  12.070 2.880 12.350 3.160 ;
        RECT  11.050 2.200 12.030 2.360 ;
        RECT  11.210 1.720 11.430 2.000 ;
        RECT  10.890 0.440 11.050 2.360 ;
        RECT  9.400 0.440 10.890 0.600 ;
        RECT  10.570 0.760 10.730 2.720 ;
        RECT  10.520 0.760 10.570 1.890 ;
        RECT  9.730 0.760 10.520 0.920 ;
        RECT  9.930 1.730 10.520 1.890 ;
        RECT  10.130 2.050 10.410 3.160 ;
        RECT  10.150 1.080 10.270 1.300 ;
        RECT  9.990 1.080 10.150 1.570 ;
        RECT  9.550 3.000 10.130 3.160 ;
        RECT  9.160 1.410 9.990 1.570 ;
        RECT  9.710 1.730 9.930 2.840 ;
        RECT  9.570 0.760 9.730 1.250 ;
        RECT  9.390 1.970 9.550 3.160 ;
        RECT  9.240 0.440 9.400 0.900 ;
        RECT  9.150 1.970 9.390 2.190 ;
        RECT  6.780 0.740 9.240 0.900 ;
        RECT  9.110 2.880 9.230 3.160 ;
        RECT  9.150 1.070 9.160 1.570 ;
        RECT  8.940 1.070 9.150 2.190 ;
        RECT  8.950 2.610 9.110 3.160 ;
        RECT  8.000 2.610 8.950 2.770 ;
        RECT  7.840 1.070 8.940 1.230 ;
        RECT  7.040 2.030 8.940 2.190 ;
        RECT  7.680 1.500 8.530 1.660 ;
        RECT  7.840 2.610 8.000 3.040 ;
        RECT  2.480 2.880 7.840 3.040 ;
        RECT  7.520 1.150 7.680 1.660 ;
        RECT  7.300 2.510 7.620 2.720 ;
        RECT  6.060 1.150 7.520 1.320 ;
        RECT  6.060 2.560 7.300 2.720 ;
        RECT  6.880 1.710 7.040 2.190 ;
        RECT  6.620 0.740 6.780 0.990 ;
        RECT  4.630 0.830 6.620 0.990 ;
        RECT  5.900 1.150 6.060 2.720 ;
        RECT  4.840 1.150 5.900 1.310 ;
        RECT  4.860 2.560 5.900 2.720 ;
        RECT  2.500 0.500 5.740 0.660 ;
        RECT  5.580 1.470 5.740 2.270 ;
        RECT  4.630 1.470 5.580 1.630 ;
        RECT  4.420 2.110 5.580 2.270 ;
        RECT  4.100 1.790 5.160 1.950 ;
        RECT  4.470 0.830 4.630 1.630 ;
        RECT  3.100 0.830 4.470 0.990 ;
        RECT  4.260 2.110 4.420 2.720 ;
        RECT  2.230 2.560 4.260 2.720 ;
        RECT  3.940 1.790 4.100 2.390 ;
        RECT  2.560 2.210 3.940 2.390 ;
        RECT  2.660 0.880 2.820 1.420 ;
        RECT  2.560 1.260 2.660 1.420 ;
        RECT  2.400 1.260 2.560 2.390 ;
        RECT  2.340 0.500 2.500 1.100 ;
        RECT  1.510 2.880 2.480 3.110 ;
        RECT  0.690 0.940 2.340 1.100 ;
        RECT  2.070 1.580 2.230 2.720 ;
        RECT  1.990 1.580 2.070 1.920 ;
        RECT  1.670 2.120 1.900 2.600 ;
        RECT  0.310 0.560 1.810 0.720 ;
        RECT  1.070 2.120 1.670 2.280 ;
        RECT  1.350 2.440 1.510 3.110 ;
        RECT  0.690 2.440 1.350 2.600 ;
        RECT  0.850 1.950 1.070 2.280 ;
        RECT  0.530 0.940 0.690 2.600 ;
        RECT  0.150 0.560 0.310 2.690 ;
    END
END DFFSHQX8TR

MACRO DFFSHQX4TR
    CLASS CORE ;
    FOREIGN DFFSHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.170 1.640 7.520 2.080 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.120 1.440 14.320 2.160 ;
        RECT  13.840 0.440 14.120 3.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.690 1.580 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.510 1.670 1.960 ;
        RECT  0.850 1.510 1.240 1.790 ;
        END
        ANTENNAGATEAREA 0.4128 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.600 -0.280 14.800 0.280 ;
        RECT  14.320 -0.280 14.600 1.280 ;
        RECT  13.600 -0.280 14.320 0.280 ;
        RECT  13.320 -0.280 13.600 0.300 ;
        RECT  11.510 -0.280 13.320 0.280 ;
        RECT  11.790 0.960 12.070 1.240 ;
        RECT  11.510 0.960 11.790 1.120 ;
        RECT  11.350 -0.280 11.510 1.120 ;
        RECT  11.230 -0.280 11.350 0.690 ;
        RECT  9.190 -0.280 11.230 0.280 ;
        RECT  8.910 -0.280 9.190 0.660 ;
        RECT  8.150 -0.280 8.910 0.280 ;
        RECT  7.870 -0.280 8.150 0.660 ;
        RECT  7.590 -0.280 7.870 0.280 ;
        RECT  7.310 -0.280 7.590 0.560 ;
        RECT  6.490 -0.280 7.310 0.280 ;
        RECT  6.210 -0.280 6.490 0.640 ;
        RECT  3.580 -0.280 6.210 0.280 ;
        RECT  3.300 -0.280 3.580 0.360 ;
        RECT  2.120 -0.280 3.300 0.280 ;
        RECT  1.900 -0.280 2.120 0.990 ;
        RECT  0.890 -0.280 1.900 0.340 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.600 3.320 14.800 3.880 ;
        RECT  14.320 2.410 14.600 3.880 ;
        RECT  13.440 3.320 14.320 3.880 ;
        RECT  13.160 3.200 13.440 3.880 ;
        RECT  11.070 3.320 13.160 3.880 ;
        RECT  10.790 3.200 11.070 3.880 ;
        RECT  8.540 3.320 10.790 3.880 ;
        RECT  8.260 2.930 8.540 3.880 ;
        RECT  6.800 3.260 8.260 3.880 ;
        RECT  6.220 3.320 6.800 3.880 ;
        RECT  5.910 3.260 6.220 3.880 ;
        RECT  4.210 3.320 5.910 3.880 ;
        RECT  3.930 3.200 4.210 3.880 ;
        RECT  3.170 3.320 3.930 3.880 ;
        RECT  2.890 3.200 3.170 3.880 ;
        RECT  1.150 3.320 2.890 3.880 ;
        RECT  0.870 3.200 1.150 3.880 ;
        RECT  0.000 3.320 0.870 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.520 0.460 13.680 3.040 ;
        RECT  12.070 0.460 13.520 0.620 ;
        RECT  12.670 2.760 13.520 3.040 ;
        RECT  13.240 1.440 13.360 2.600 ;
        RECT  13.200 0.780 13.240 2.600 ;
        RECT  13.080 0.780 13.200 1.720 ;
        RECT  12.270 2.440 13.200 2.600 ;
        RECT  12.810 0.780 13.080 0.990 ;
        RECT  12.630 2.000 13.000 2.280 ;
        RECT  12.510 2.760 12.670 3.160 ;
        RECT  12.470 1.100 12.630 2.280 ;
        RECT  12.070 2.880 12.510 3.160 ;
        RECT  12.350 1.100 12.470 1.320 ;
        RECT  11.430 1.650 12.470 1.810 ;
        RECT  10.690 2.440 12.270 2.720 ;
        RECT  11.790 0.460 12.070 0.630 ;
        RECT  11.750 2.060 12.030 2.280 ;
        RECT  11.010 2.060 11.750 2.220 ;
        RECT  11.370 1.590 11.430 1.810 ;
        RECT  11.210 1.590 11.370 1.870 ;
        RECT  10.850 0.480 11.010 2.220 ;
        RECT  9.510 0.480 10.850 0.640 ;
        RECT  10.530 0.820 10.690 2.720 ;
        RECT  9.830 0.820 10.530 0.980 ;
        RECT  10.510 1.840 10.530 2.720 ;
        RECT  9.870 1.840 10.510 2.000 ;
        RECT  10.130 2.430 10.350 3.160 ;
        RECT  10.150 1.140 10.270 1.360 ;
        RECT  9.990 1.140 10.150 1.680 ;
        RECT  9.490 3.000 10.130 3.160 ;
        RECT  8.670 1.520 9.990 1.680 ;
        RECT  9.710 1.840 9.870 2.840 ;
        RECT  9.670 0.820 9.830 1.360 ;
        RECT  9.510 1.140 9.670 1.360 ;
        RECT  9.350 0.480 9.510 0.980 ;
        RECT  9.330 2.240 9.490 3.160 ;
        RECT  9.330 0.820 9.350 0.980 ;
        RECT  9.130 0.820 9.330 1.200 ;
        RECT  8.610 2.240 9.330 2.400 ;
        RECT  9.110 2.880 9.170 3.160 ;
        RECT  7.070 0.820 9.130 0.980 ;
        RECT  8.950 2.610 9.110 3.160 ;
        RECT  7.920 2.610 8.950 2.770 ;
        RECT  8.610 1.140 8.670 1.680 ;
        RECT  8.450 1.140 8.610 2.400 ;
        RECT  8.390 1.140 8.450 1.300 ;
        RECT  6.960 2.240 8.450 2.400 ;
        RECT  8.220 1.420 8.280 1.700 ;
        RECT  8.060 1.220 8.220 1.700 ;
        RECT  6.770 1.220 8.060 1.400 ;
        RECT  7.760 2.610 7.920 3.100 ;
        RECT  5.460 2.880 7.760 3.100 ;
        RECT  6.460 2.560 7.600 2.720 ;
        RECT  6.950 0.540 7.070 0.980 ;
        RECT  6.800 1.560 6.960 2.400 ;
        RECT  6.790 0.540 6.950 0.960 ;
        RECT  6.680 1.560 6.800 1.840 ;
        RECT  4.950 0.800 6.790 0.960 ;
        RECT  6.460 1.120 6.770 1.400 ;
        RECT  6.300 1.120 6.460 2.720 ;
        RECT  5.330 1.120 6.300 1.280 ;
        RECT  6.080 2.390 6.300 2.720 ;
        RECT  5.860 1.810 6.140 2.130 ;
        RECT  5.140 2.560 6.080 2.720 ;
        RECT  4.700 1.810 5.860 1.970 ;
        RECT  5.300 2.880 5.460 3.160 ;
        RECT  5.110 1.120 5.330 1.400 ;
        RECT  4.700 3.000 5.300 3.160 ;
        RECT  4.860 2.130 5.140 2.840 ;
        RECT  4.790 0.800 4.950 1.120 ;
        RECT  4.190 0.960 4.790 1.120 ;
        RECT  4.540 1.460 4.700 3.160 ;
        RECT  4.350 0.440 4.630 0.720 ;
        RECT  4.350 1.460 4.540 1.740 ;
        RECT  4.500 2.880 4.540 3.160 ;
        RECT  2.430 2.880 4.500 3.040 ;
        RECT  4.190 1.950 4.380 2.230 ;
        RECT  2.600 0.520 4.350 0.680 ;
        RECT  4.030 0.960 4.190 2.600 ;
        RECT  3.060 0.960 4.030 1.120 ;
        RECT  3.690 2.440 4.030 2.600 ;
        RECT  3.410 2.440 3.690 2.720 ;
        RECT  2.210 2.560 3.410 2.720 ;
        RECT  2.780 0.840 3.060 1.120 ;
        RECT  2.530 2.120 2.770 2.400 ;
        RECT  2.530 0.520 2.600 0.990 ;
        RECT  2.440 0.520 2.530 2.400 ;
        RECT  2.380 0.710 2.440 2.400 ;
        RECT  1.510 2.880 2.430 3.160 ;
        RECT  2.370 0.830 2.380 2.400 ;
        RECT  2.150 1.700 2.210 2.720 ;
        RECT  2.050 1.580 2.150 2.720 ;
        RECT  1.870 1.580 2.050 1.860 ;
        RECT  1.670 2.120 1.890 2.720 ;
        RECT  1.460 0.500 1.740 0.780 ;
        RECT  1.070 2.120 1.670 2.280 ;
        RECT  1.350 2.440 1.510 3.160 ;
        RECT  0.370 0.620 1.460 0.780 ;
        RECT  1.130 1.030 1.410 1.310 ;
        RECT  0.690 2.440 1.350 2.600 ;
        RECT  0.690 1.150 1.130 1.310 ;
        RECT  0.850 1.950 1.070 2.280 ;
        RECT  0.530 1.150 0.690 2.600 ;
        RECT  0.250 0.620 0.370 1.050 ;
        RECT  0.250 2.410 0.370 2.690 ;
        RECT  0.210 0.620 0.250 2.690 ;
        RECT  0.090 0.770 0.210 2.690 ;
    END
END DFFSHQX4TR

MACRO DFFSHQX2TR
    CLASS CORE ;
    FOREIGN DFFSHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.280 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.840 0.440 11.120 2.190 ;
        RECT  10.830 0.440 10.840 1.230 ;
        RECT  10.710 1.910 10.840 2.190 ;
        RECT  10.430 1.910 10.710 2.650 ;
        END
        ANTENNADIFFAREA 2.676 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.230 2.720 1.600 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.180 0.760 1.560 ;
        END
        ANTENNAGATEAREA 0.24 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.590 -0.280 11.200 0.280 ;
        RECT  10.310 -0.280 10.590 0.400 ;
        RECT  9.470 -0.280 10.310 0.280 ;
        RECT  9.190 -0.280 9.470 0.360 ;
        RECT  8.550 -0.280 9.190 0.340 ;
        RECT  8.270 -0.280 8.550 0.360 ;
        RECT  5.910 -0.280 8.270 0.280 ;
        RECT  5.630 -0.280 5.910 0.290 ;
        RECT  3.680 -0.280 5.630 0.280 ;
        RECT  3.400 -0.280 3.680 0.290 ;
        RECT  2.410 -0.280 3.400 0.280 ;
        RECT  2.130 -0.280 2.410 0.290 ;
        RECT  0.890 -0.280 2.130 0.280 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.110 3.320 11.200 3.880 ;
        RECT  10.190 3.200 11.110 3.880 ;
        RECT  9.910 2.800 10.190 3.880 ;
        RECT  7.310 3.320 9.910 3.880 ;
        RECT  7.030 3.200 7.310 3.880 ;
        RECT  6.270 3.320 7.030 3.880 ;
        RECT  5.990 3.200 6.270 3.880 ;
        RECT  5.200 3.320 5.990 3.880 ;
        RECT  4.920 3.200 5.200 3.880 ;
        RECT  3.670 3.320 4.920 3.880 ;
        RECT  3.450 3.200 3.670 3.880 ;
        RECT  2.200 3.320 3.450 3.880 ;
        RECT  1.920 3.200 2.200 3.880 ;
        RECT  0.760 3.260 1.920 3.880 ;
        RECT  0.480 2.800 0.760 3.880 ;
        RECT  0.000 3.320 0.480 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.350 1.470 10.680 1.750 ;
        RECT  10.190 0.580 10.350 1.750 ;
        RECT  9.990 0.580 10.190 0.740 ;
        RECT  10.110 1.470 10.190 1.750 ;
        RECT  9.950 1.470 10.110 2.430 ;
        RECT  9.670 0.920 10.030 1.200 ;
        RECT  9.710 0.440 9.990 0.740 ;
        RECT  8.710 2.270 9.950 2.430 ;
        RECT  9.670 1.830 9.790 2.110 ;
        RECT  7.390 0.520 9.710 0.740 ;
        RECT  9.510 0.920 9.670 2.110 ;
        RECT  8.030 0.920 9.510 1.140 ;
        RECT  9.310 1.430 9.510 1.710 ;
        RECT  9.030 1.360 9.150 1.640 ;
        RECT  8.870 1.360 9.030 1.900 ;
        RECT  7.150 1.740 8.870 1.900 ;
        RECT  7.470 1.300 8.710 1.580 ;
        RECT  8.590 2.270 8.710 3.160 ;
        RECT  8.430 2.060 8.590 3.160 ;
        RECT  7.430 2.060 8.430 2.280 ;
        RECT  7.950 2.440 8.230 3.160 ;
        RECT  6.830 2.440 7.950 2.600 ;
        RECT  7.260 2.760 7.540 3.040 ;
        RECT  7.310 0.900 7.470 1.580 ;
        RECT  7.230 0.900 7.310 1.060 ;
        RECT  5.780 2.880 7.260 3.040 ;
        RECT  6.950 0.440 7.230 1.060 ;
        RECT  6.990 1.220 7.150 1.900 ;
        RECT  6.790 1.220 6.990 1.380 ;
        RECT  6.230 0.440 6.950 0.600 ;
        RECT  6.670 1.540 6.830 2.720 ;
        RECT  6.630 0.770 6.790 1.380 ;
        RECT  6.470 1.540 6.670 1.700 ;
        RECT  5.860 2.440 6.670 2.720 ;
        RECT  3.480 0.770 6.630 0.930 ;
        RECT  6.230 1.860 6.510 2.160 ;
        RECT  6.310 1.090 6.470 1.700 ;
        RECT  6.190 1.090 6.310 1.310 ;
        RECT  6.070 0.440 6.230 0.610 ;
        RECT  6.150 1.860 6.230 2.020 ;
        RECT  5.990 1.520 6.150 2.020 ;
        RECT  1.890 0.450 6.070 0.610 ;
        RECT  5.390 1.520 5.990 1.680 ;
        RECT  5.830 2.180 5.860 2.720 ;
        RECT  5.700 1.840 5.830 2.720 ;
        RECT  5.500 2.880 5.780 3.160 ;
        RECT  5.550 1.840 5.700 2.340 ;
        RECT  5.390 2.500 5.540 2.720 ;
        RECT  4.470 2.880 5.500 3.040 ;
        RECT  5.230 1.090 5.390 2.720 ;
        RECT  3.800 1.090 5.230 1.310 ;
        RECT  4.310 1.800 4.470 3.040 ;
        RECT  4.240 1.800 4.310 1.960 ;
        RECT  3.280 2.880 4.310 3.040 ;
        RECT  3.960 1.680 4.240 1.960 ;
        RECT  3.870 2.500 4.150 2.720 ;
        RECT  3.800 2.120 4.030 2.340 ;
        RECT  2.960 2.500 3.870 2.660 ;
        RECT  3.640 1.090 3.800 2.340 ;
        RECT  3.320 0.770 3.480 2.340 ;
        RECT  3.000 0.770 3.320 1.120 ;
        RECT  2.790 2.120 3.320 2.340 ;
        RECT  3.120 2.880 3.280 3.120 ;
        RECT  2.520 2.960 3.120 3.120 ;
        RECT  2.680 2.500 2.960 2.800 ;
        RECT  2.210 0.790 2.810 1.070 ;
        RECT  2.360 2.500 2.680 2.660 ;
        RECT  2.360 2.820 2.520 3.120 ;
        RECT  2.210 1.760 2.360 2.660 ;
        RECT  1.690 2.820 2.360 2.980 ;
        RECT  2.200 0.790 2.210 2.660 ;
        RECT  2.050 0.790 2.200 1.920 ;
        RECT  1.890 2.080 2.040 2.360 ;
        RECT  1.730 0.450 1.890 2.360 ;
        RECT  1.610 0.650 1.730 0.930 ;
        RECT  1.240 1.690 1.730 1.970 ;
        RECT  1.530 2.540 1.690 2.980 ;
        RECT  1.410 2.540 1.530 2.820 ;
        RECT  1.170 0.440 1.450 0.720 ;
        RECT  1.080 2.540 1.410 2.700 ;
        RECT  1.080 0.880 1.290 1.160 ;
        RECT  0.320 0.560 1.170 0.720 ;
        RECT  0.920 0.880 1.080 2.700 ;
        RECT  0.160 0.560 0.320 2.300 ;
        RECT  0.090 0.840 0.160 1.120 ;
        RECT  0.100 2.020 0.160 2.300 ;
    END
END DFFSHQX2TR

MACRO DFFSHQX1TR
    CLASS CORE ;
    FOREIGN DFFSHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.060 1.640 3.220 1.960 ;
        RECT  2.880 1.600 3.060 1.960 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.650 0.840 9.920 2.650 ;
        END
        ANTENNADIFFAREA 1.92 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.240 2.720 1.560 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.740 -0.280 10.000 0.280 ;
        RECT  2.120 -0.280 3.740 0.340 ;
        RECT  0.930 -0.280 2.120 0.280 ;
        RECT  0.650 -0.280 0.930 0.400 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.390 3.320 10.000 3.880 ;
        RECT  8.450 2.770 9.390 3.880 ;
        RECT  6.410 3.320 8.450 3.880 ;
        RECT  5.100 3.260 6.410 3.880 ;
        RECT  3.860 3.320 5.100 3.880 ;
        RECT  3.580 3.200 3.860 3.880 ;
        RECT  2.400 3.320 3.580 3.880 ;
        RECT  2.120 3.200 2.400 3.880 ;
        RECT  0.810 3.260 2.120 3.880 ;
        RECT  0.530 2.800 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.310 1.300 9.430 1.580 ;
        RECT  9.150 0.440 9.310 2.510 ;
        RECT  7.390 0.440 9.150 0.660 ;
        RECT  7.430 2.350 9.150 2.510 ;
        RECT  8.830 1.030 8.950 1.310 ;
        RECT  8.830 1.910 8.950 2.190 ;
        RECT  8.670 1.030 8.830 2.190 ;
        RECT  8.290 1.350 8.670 1.630 ;
        RECT  8.230 0.820 8.510 1.100 ;
        RECT  8.130 0.940 8.230 1.100 ;
        RECT  8.010 0.940 8.130 1.820 ;
        RECT  7.970 0.940 8.010 2.190 ;
        RECT  7.850 1.540 7.970 2.190 ;
        RECT  7.310 2.030 7.850 2.190 ;
        RECT  6.570 2.940 7.760 3.160 ;
        RECT  7.470 0.820 7.690 1.870 ;
        RECT  7.230 0.820 7.470 0.980 ;
        RECT  7.150 2.350 7.430 2.630 ;
        RECT  7.150 1.140 7.310 2.190 ;
        RECT  7.070 0.440 7.230 0.980 ;
        RECT  6.910 1.140 7.150 1.300 ;
        RECT  4.060 0.440 7.070 0.600 ;
        RECT  6.830 1.460 6.990 2.500 ;
        RECT  6.750 0.760 6.910 1.300 ;
        RECT  6.590 1.460 6.830 1.620 ;
        RECT  6.240 2.220 6.830 2.500 ;
        RECT  4.380 0.760 6.750 0.920 ;
        RECT  6.450 1.780 6.670 2.060 ;
        RECT  6.310 1.080 6.590 1.620 ;
        RECT  4.940 2.940 6.570 3.100 ;
        RECT  5.800 1.780 6.450 1.940 ;
        RECT  6.080 2.100 6.240 2.500 ;
        RECT  5.960 2.100 6.080 2.380 ;
        RECT  5.640 1.140 5.800 2.780 ;
        RECT  4.940 1.140 5.640 1.300 ;
        RECT  5.320 2.500 5.640 2.780 ;
        RECT  4.940 2.060 5.480 2.340 ;
        RECT  4.660 1.080 4.940 1.300 ;
        RECT  4.780 1.520 4.940 3.100 ;
        RECT  4.300 1.520 4.780 1.680 ;
        RECT  4.180 2.940 4.780 3.100 ;
        RECT  3.860 1.140 4.660 1.300 ;
        RECT  4.400 2.500 4.620 2.780 ;
        RECT  3.860 1.910 4.420 2.190 ;
        RECT  3.100 2.500 4.400 2.660 ;
        RECT  4.220 0.760 4.380 0.980 ;
        RECT  4.020 1.460 4.300 1.680 ;
        RECT  3.540 0.820 4.220 0.980 ;
        RECT  4.020 2.880 4.180 3.100 ;
        RECT  3.900 0.440 4.060 0.660 ;
        RECT  3.420 2.880 4.020 3.040 ;
        RECT  1.840 0.500 3.900 0.660 ;
        RECT  3.700 1.140 3.860 2.190 ;
        RECT  3.380 0.820 3.540 2.280 ;
        RECT  3.260 2.880 3.420 3.130 ;
        RECT  3.020 0.820 3.380 1.040 ;
        RECT  3.020 2.120 3.380 2.280 ;
        RECT  2.720 2.970 3.260 3.130 ;
        RECT  2.880 2.500 3.100 2.810 ;
        RECT  2.510 2.500 2.880 2.660 ;
        RECT  2.270 0.820 2.840 1.040 ;
        RECT  2.560 2.820 2.720 3.130 ;
        RECT  1.730 2.820 2.560 2.980 ;
        RECT  2.350 1.740 2.510 2.660 ;
        RECT  2.270 1.740 2.350 1.900 ;
        RECT  2.110 0.820 2.270 1.900 ;
        RECT  1.910 2.060 2.190 2.340 ;
        RECT  1.840 2.060 1.910 2.220 ;
        RECT  1.680 0.500 1.840 2.220 ;
        RECT  1.570 2.380 1.730 2.980 ;
        RECT  1.560 0.500 1.680 0.960 ;
        RECT  1.250 1.760 1.680 2.040 ;
        RECT  1.450 2.380 1.570 2.660 ;
        RECT  1.090 2.380 1.450 2.540 ;
        RECT  1.120 0.440 1.400 0.720 ;
        RECT  1.090 1.030 1.370 1.310 ;
        RECT  0.310 0.560 1.120 0.720 ;
        RECT  0.930 1.030 1.090 2.540 ;
        RECT  0.150 0.560 0.310 2.320 ;
    END
END DFFSHQX1TR

MACRO DFFSXLTR
    CLASS CORE ;
    FOREIGN DFFSXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.240 6.080 1.640 ;
        RECT  5.520 1.480 5.680 3.160 ;
        RECT  4.760 2.940 5.520 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.030 1.030 8.320 2.360 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 1.030 7.270 1.310 ;
        RECT  7.050 1.030 7.210 2.760 ;
        RECT  6.880 2.350 7.050 2.760 ;
        END
        ANTENNADIFFAREA 1.014 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.370 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 2.060 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.380 -0.280 8.400 0.280 ;
        RECT  6.100 -0.280 6.380 0.700 ;
        RECT  1.890 -0.280 6.100 0.280 ;
        RECT  1.610 -0.280 1.890 0.330 ;
        RECT  0.370 -0.280 1.610 0.280 ;
        RECT  0.090 -0.280 0.370 0.330 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.940 3.320 8.400 3.880 ;
        RECT  7.570 3.260 7.940 3.880 ;
        RECT  6.190 3.320 7.570 3.880 ;
        RECT  5.910 2.400 6.190 3.880 ;
        RECT  4.600 3.320 5.910 3.880 ;
        RECT  4.380 2.850 4.600 3.880 ;
        RECT  2.940 3.320 4.380 3.880 ;
        RECT  2.660 2.990 2.940 3.880 ;
        RECT  1.890 3.320 2.660 3.880 ;
        RECT  1.610 2.990 1.890 3.880 ;
        RECT  0.310 3.260 1.610 3.880 ;
        RECT  0.150 2.770 0.310 3.880 ;
        RECT  0.000 3.320 0.150 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.750 1.620 7.870 1.900 ;
        RECT  7.590 0.710 7.750 3.080 ;
        RECT  7.080 0.710 7.590 0.870 ;
        RECT  7.570 1.620 7.590 1.900 ;
        RECT  6.870 2.920 7.590 3.080 ;
        RECT  6.800 0.440 7.080 0.870 ;
        RECT  6.710 1.030 6.890 2.190 ;
        RECT  6.590 2.920 6.870 3.130 ;
        RECT  6.590 1.030 6.710 1.310 ;
        RECT  5.840 1.910 6.710 2.190 ;
        RECT  6.430 1.470 6.490 1.750 ;
        RECT  6.270 0.920 6.430 1.750 ;
        RECT  5.360 0.920 6.270 1.080 ;
        RECT  5.520 0.440 5.800 0.760 ;
        RECT  3.020 0.440 5.520 0.600 ;
        RECT  5.200 0.760 5.360 2.780 ;
        RECT  4.660 0.760 5.200 0.920 ;
        RECT  4.880 2.380 5.200 2.780 ;
        RECT  4.820 1.200 5.040 2.220 ;
        RECT  4.660 2.380 4.880 2.540 ;
        RECT  4.620 1.200 4.820 1.360 ;
        RECT  4.380 1.910 4.660 2.540 ;
        RECT  4.220 1.080 4.620 1.360 ;
        RECT  3.480 0.760 4.380 0.920 ;
        RECT  4.060 1.080 4.220 3.160 ;
        RECT  3.640 1.080 4.060 1.300 ;
        RECT  3.500 3.000 4.060 3.160 ;
        RECT  3.680 1.460 3.900 2.590 ;
        RECT  3.480 1.460 3.680 1.620 ;
        RECT  3.220 2.220 3.500 3.160 ;
        RECT  3.320 0.760 3.480 1.620 ;
        RECT  2.540 1.450 3.320 1.610 ;
        RECT  3.050 1.780 3.270 2.060 ;
        RECT  3.100 2.990 3.220 3.160 ;
        RECT  2.890 1.780 3.050 2.830 ;
        RECT  2.860 0.440 3.020 1.290 ;
        RECT  2.450 2.670 2.890 2.830 ;
        RECT  2.740 1.010 2.860 1.290 ;
        RECT  1.070 2.330 2.730 2.490 ;
        RECT  2.380 1.030 2.540 1.610 ;
        RECT  2.380 1.910 2.500 2.130 ;
        RECT  0.750 0.550 2.450 0.830 ;
        RECT  2.170 2.670 2.450 2.890 ;
        RECT  2.220 1.030 2.380 2.130 ;
        RECT  1.770 1.320 2.220 1.480 ;
        RECT  1.370 2.670 2.170 2.830 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.090 2.670 1.370 2.900 ;
        RECT  0.750 2.670 1.090 2.830 ;
        RECT  0.910 0.990 1.070 2.490 ;
        RECT  0.590 0.550 0.750 2.830 ;
    END
END DFFSXLTR

MACRO DFFSX4TR
    CLASS CORE ;
    FOREIGN DFFSX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.240 5.920 1.640 ;
        RECT  5.620 1.480 5.680 1.640 ;
        RECT  5.460 1.480 5.620 3.160 ;
        RECT  4.800 2.940 5.460 3.160 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.880 1.090 9.120 2.210 ;
        RECT  8.750 1.090 8.880 1.250 ;
        RECT  8.750 1.930 8.880 2.210 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 0.770 9.440 2.560 ;
        RECT  8.070 0.770 9.280 0.930 ;
        RECT  8.320 2.400 9.280 2.560 ;
        RECT  8.080 1.840 8.320 2.560 ;
        RECT  8.070 1.930 8.080 2.560 ;
        RECT  7.790 0.570 8.070 1.250 ;
        RECT  7.790 1.930 8.070 3.010 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 2.070 1.960 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.510 -0.280 9.600 0.280 ;
        RECT  9.230 -0.280 9.510 0.610 ;
        RECT  8.550 -0.280 9.230 0.280 ;
        RECT  8.270 -0.280 8.550 0.610 ;
        RECT  7.820 -0.280 8.270 0.290 ;
        RECT  7.590 -0.280 7.820 0.280 ;
        RECT  7.320 -0.280 7.590 1.220 ;
        RECT  6.270 -0.280 7.320 0.280 ;
        RECT  5.990 -0.280 6.270 0.760 ;
        RECT  1.930 -0.280 5.990 0.280 ;
        RECT  1.650 -0.280 1.930 0.390 ;
        RECT  0.370 -0.280 1.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.400 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.510 3.320 9.600 3.880 ;
        RECT  9.230 2.720 9.510 3.880 ;
        RECT  8.550 3.320 9.230 3.880 ;
        RECT  8.270 2.720 8.550 3.880 ;
        RECT  7.590 3.320 8.270 3.880 ;
        RECT  7.310 2.970 7.590 3.880 ;
        RECT  6.080 3.320 7.310 3.880 ;
        RECT  5.800 2.800 6.080 3.880 ;
        RECT  4.640 3.320 5.800 3.880 ;
        RECT  4.420 2.850 4.640 3.880 ;
        RECT  2.980 3.320 4.420 3.880 ;
        RECT  2.700 3.000 2.980 3.880 ;
        RECT  1.930 3.320 2.700 3.880 ;
        RECT  1.650 3.000 1.930 3.880 ;
        RECT  0.370 3.260 1.650 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.250 1.410 8.670 1.660 ;
        RECT  7.110 1.380 7.250 2.780 ;
        RECT  7.090 1.030 7.110 2.780 ;
        RECT  6.830 1.030 7.090 1.660 ;
        RECT  7.030 2.620 7.090 2.780 ;
        RECT  6.750 2.620 7.030 3.130 ;
        RECT  6.670 0.540 6.750 0.820 ;
        RECT  6.510 0.540 6.670 2.460 ;
        RECT  6.470 0.540 6.510 0.820 ;
        RECT  6.030 2.300 6.510 2.460 ;
        RECT  6.240 1.360 6.350 1.640 ;
        RECT  6.080 0.920 6.240 1.640 ;
        RECT  5.300 0.920 6.080 1.080 ;
        RECT  5.780 1.910 6.030 2.460 ;
        RECT  5.460 0.440 5.740 0.760 ;
        RECT  2.910 0.440 5.460 0.600 ;
        RECT  5.140 0.760 5.300 2.780 ;
        RECT  4.700 0.760 5.140 0.920 ;
        RECT  4.920 2.380 5.140 2.780 ;
        RECT  4.820 1.200 4.980 2.220 ;
        RECT  4.580 2.380 4.920 2.540 ;
        RECT  4.660 1.200 4.820 1.360 ;
        RECT  4.260 1.080 4.660 1.360 ;
        RECT  4.420 1.910 4.580 2.540 ;
        RECT  3.290 0.760 4.420 0.920 ;
        RECT  4.100 1.080 4.260 3.160 ;
        RECT  3.590 1.080 4.100 1.300 ;
        RECT  3.540 3.000 4.100 3.160 ;
        RECT  3.720 1.460 3.940 2.590 ;
        RECT  3.290 1.460 3.720 1.620 ;
        RECT  3.320 2.220 3.540 3.160 ;
        RECT  3.160 1.780 3.350 2.060 ;
        RECT  3.140 3.000 3.320 3.160 ;
        RECT  3.130 0.760 3.290 1.620 ;
        RECT  3.000 1.780 3.160 2.840 ;
        RECT  2.490 1.460 3.130 1.620 ;
        RECT  2.510 2.680 3.000 2.840 ;
        RECT  2.750 0.440 2.910 1.290 ;
        RECT  2.530 2.300 2.810 2.520 ;
        RECT  2.690 1.010 2.750 1.290 ;
        RECT  2.390 1.910 2.540 2.130 ;
        RECT  1.170 2.300 2.530 2.460 ;
        RECT  2.230 2.680 2.510 2.910 ;
        RECT  2.390 1.030 2.490 1.620 ;
        RECT  2.170 0.450 2.450 0.830 ;
        RECT  2.230 1.030 2.390 2.130 ;
        RECT  2.210 1.030 2.230 1.480 ;
        RECT  1.410 2.680 2.230 2.840 ;
        RECT  1.770 1.320 2.210 1.480 ;
        RECT  0.730 0.550 2.170 0.830 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.130 2.680 1.410 2.900 ;
        RECT  1.070 2.180 1.170 2.460 ;
        RECT  0.730 2.680 1.130 2.840 ;
        RECT  0.910 0.990 1.070 2.460 ;
        RECT  0.570 0.550 0.730 2.840 ;
    END
END DFFSX4TR

MACRO DFFSX2TR
    CLASS CORE ;
    FOREIGN DFFSX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.240 5.920 1.640 ;
        RECT  5.520 1.240 5.680 3.160 ;
        RECT  4.760 2.940 5.520 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.610 8.320 3.140 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 1.030 7.270 2.760 ;
        RECT  7.050 1.030 7.110 1.310 ;
        RECT  6.880 2.440 7.110 2.760 ;
        END
        ANTENNADIFFAREA 3.046 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.370 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.640 2.060 1.960 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.370 -0.280 8.400 0.280 ;
        RECT  6.090 -0.280 6.370 0.680 ;
        RECT  1.890 -0.280 6.090 0.280 ;
        RECT  1.610 -0.280 1.890 0.330 ;
        RECT  0.370 -0.280 1.610 0.280 ;
        RECT  0.090 -0.280 0.370 0.330 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.790 3.320 8.400 3.880 ;
        RECT  7.510 3.260 7.790 3.880 ;
        RECT  6.170 3.320 7.510 3.880 ;
        RECT  5.890 2.460 6.170 3.880 ;
        RECT  4.600 3.320 5.890 3.880 ;
        RECT  4.380 2.850 4.600 3.880 ;
        RECT  2.940 3.320 4.380 3.880 ;
        RECT  2.660 2.990 2.940 3.880 ;
        RECT  1.890 3.320 2.660 3.880 ;
        RECT  1.610 2.990 1.890 3.880 ;
        RECT  0.360 3.260 1.610 3.880 ;
        RECT  0.090 2.770 0.360 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.800 1.470 7.920 1.750 ;
        RECT  7.640 0.650 7.800 3.080 ;
        RECT  6.930 0.650 7.640 0.810 ;
        RECT  6.870 2.920 7.640 3.080 ;
        RECT  6.650 0.440 6.930 0.810 ;
        RECT  6.710 0.970 6.890 2.190 ;
        RECT  6.590 2.920 6.870 3.130 ;
        RECT  6.400 0.970 6.710 1.250 ;
        RECT  5.840 1.910 6.710 2.190 ;
        RECT  6.240 1.470 6.490 1.750 ;
        RECT  6.080 0.920 6.240 1.750 ;
        RECT  5.360 0.920 6.080 1.080 ;
        RECT  5.330 0.440 5.610 0.740 ;
        RECT  5.200 0.920 5.360 2.780 ;
        RECT  2.930 0.440 5.330 0.600 ;
        RECT  4.850 0.920 5.200 1.080 ;
        RECT  4.880 2.380 5.200 2.780 ;
        RECT  4.820 1.240 5.040 2.220 ;
        RECT  4.660 2.380 4.880 2.540 ;
        RECT  4.690 0.760 4.850 1.080 ;
        RECT  4.470 1.240 4.820 1.400 ;
        RECT  4.570 0.760 4.690 0.920 ;
        RECT  4.380 1.910 4.660 2.540 ;
        RECT  4.220 1.080 4.470 1.400 ;
        RECT  3.390 0.760 4.290 0.920 ;
        RECT  4.060 1.080 4.220 3.160 ;
        RECT  3.550 1.080 4.060 1.300 ;
        RECT  3.500 3.000 4.060 3.160 ;
        RECT  3.680 1.460 3.900 2.590 ;
        RECT  3.390 1.460 3.680 1.620 ;
        RECT  3.220 2.220 3.500 3.160 ;
        RECT  3.320 0.760 3.390 1.620 ;
        RECT  3.230 0.760 3.320 1.610 ;
        RECT  3.050 1.780 3.270 2.060 ;
        RECT  2.450 1.450 3.230 1.610 ;
        RECT  3.100 2.990 3.220 3.160 ;
        RECT  2.890 1.780 3.050 2.830 ;
        RECT  2.770 0.440 2.930 1.290 ;
        RECT  2.450 2.670 2.890 2.830 ;
        RECT  2.650 1.010 2.770 1.290 ;
        RECT  1.070 2.330 2.730 2.490 ;
        RECT  2.380 1.910 2.500 2.130 ;
        RECT  2.380 1.030 2.450 1.610 ;
        RECT  2.170 2.670 2.450 2.890 ;
        RECT  0.750 0.550 2.410 0.830 ;
        RECT  2.220 1.030 2.380 2.130 ;
        RECT  2.130 1.030 2.220 1.480 ;
        RECT  1.370 2.670 2.170 2.830 ;
        RECT  1.770 1.320 2.130 1.480 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.090 2.670 1.370 2.900 ;
        RECT  0.750 2.670 1.090 2.830 ;
        RECT  0.910 0.990 1.070 2.490 ;
        RECT  0.590 0.550 0.750 2.830 ;
    END
END DFFSX2TR

MACRO DFFSX1TR
    CLASS CORE ;
    FOREIGN DFFSX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.240 6.080 1.640 ;
        RECT  5.520 1.240 5.680 3.160 ;
        RECT  4.760 2.940 5.520 3.160 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.030 1.030 8.320 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.270 1.090 7.330 1.250 ;
        RECT  7.050 1.090 7.270 2.760 ;
        RECT  6.880 2.440 7.050 2.760 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.370 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.640 2.060 1.980 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.380 -0.280 8.400 0.280 ;
        RECT  6.100 -0.280 6.380 0.700 ;
        RECT  1.890 -0.280 6.100 0.280 ;
        RECT  1.610 -0.280 1.890 0.330 ;
        RECT  0.370 -0.280 1.610 0.280 ;
        RECT  0.090 -0.280 0.370 0.330 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.940 3.320 8.400 3.880 ;
        RECT  7.570 3.260 7.940 3.880 ;
        RECT  6.210 3.320 7.570 3.880 ;
        RECT  5.930 2.800 6.210 3.880 ;
        RECT  4.600 3.320 5.930 3.880 ;
        RECT  4.380 2.850 4.600 3.880 ;
        RECT  2.940 3.320 4.380 3.880 ;
        RECT  2.660 2.990 2.940 3.880 ;
        RECT  1.890 3.320 2.660 3.880 ;
        RECT  1.610 2.990 1.890 3.880 ;
        RECT  0.370 3.260 1.610 3.880 ;
        RECT  0.090 2.770 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.690 0.710 7.870 3.080 ;
        RECT  7.080 0.710 7.690 0.870 ;
        RECT  6.870 2.920 7.690 3.080 ;
        RECT  6.800 0.440 7.080 0.870 ;
        RECT  6.710 1.030 6.890 2.190 ;
        RECT  6.590 2.920 6.870 3.130 ;
        RECT  6.590 1.030 6.710 1.310 ;
        RECT  5.840 1.910 6.710 2.190 ;
        RECT  6.430 1.470 6.490 1.750 ;
        RECT  6.270 0.920 6.430 1.750 ;
        RECT  5.360 0.920 6.270 1.080 ;
        RECT  5.520 0.440 5.800 0.760 ;
        RECT  3.020 0.440 5.520 0.600 ;
        RECT  5.200 0.760 5.360 2.780 ;
        RECT  4.660 0.760 5.200 0.920 ;
        RECT  4.880 2.380 5.200 2.780 ;
        RECT  4.820 1.200 5.040 2.220 ;
        RECT  4.660 2.380 4.880 2.540 ;
        RECT  4.620 1.200 4.820 1.360 ;
        RECT  4.380 1.910 4.660 2.540 ;
        RECT  4.220 1.080 4.620 1.360 ;
        RECT  3.480 0.760 4.380 0.920 ;
        RECT  4.060 1.080 4.220 3.160 ;
        RECT  3.640 1.080 4.060 1.300 ;
        RECT  3.500 3.000 4.060 3.160 ;
        RECT  3.680 1.460 3.900 2.590 ;
        RECT  3.480 1.460 3.680 1.620 ;
        RECT  3.220 2.220 3.500 3.160 ;
        RECT  3.320 0.760 3.480 1.620 ;
        RECT  2.540 1.450 3.320 1.610 ;
        RECT  3.050 1.780 3.270 2.060 ;
        RECT  3.100 2.990 3.220 3.160 ;
        RECT  2.890 1.780 3.050 2.830 ;
        RECT  2.860 0.440 3.020 1.290 ;
        RECT  2.450 2.670 2.890 2.830 ;
        RECT  2.740 1.010 2.860 1.290 ;
        RECT  1.070 2.330 2.730 2.490 ;
        RECT  2.380 1.030 2.540 1.610 ;
        RECT  2.380 1.910 2.500 2.130 ;
        RECT  0.750 0.550 2.450 0.830 ;
        RECT  2.170 2.670 2.450 2.890 ;
        RECT  2.220 1.030 2.380 2.130 ;
        RECT  1.770 1.320 2.220 1.480 ;
        RECT  1.370 2.670 2.170 2.830 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.090 2.670 1.370 2.900 ;
        RECT  0.750 2.670 1.090 2.830 ;
        RECT  0.910 0.990 1.070 2.490 ;
        RECT  0.590 0.550 0.750 2.830 ;
    END
END DFFSX1TR

MACRO DFFRHQX8TR
    CLASS CORE ;
    FOREIGN DFFRHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.880 1.640 10.040 1.920 ;
        RECT  7.920 1.640 9.880 1.800 ;
        RECT  7.760 1.270 7.920 1.800 ;
        RECT  7.720 1.640 7.760 1.800 ;
        RECT  7.280 1.640 7.720 2.000 ;
        RECT  6.680 1.640 7.280 1.800 ;
        RECT  6.520 1.260 6.680 1.800 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.150 0.630 13.440 3.090 ;
        RECT  12.470 1.440 13.150 2.160 ;
        RECT  12.190 0.470 12.470 3.160 ;
        END
        ANTENNADIFFAREA 7.992 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.240 2.320 1.640 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.840 1.730 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.910 -0.280 14.000 0.280 ;
        RECT  13.620 -0.280 13.910 1.160 ;
        RECT  12.950 -0.280 13.620 0.280 ;
        RECT  12.670 -0.280 12.950 1.150 ;
        RECT  11.950 -0.280 12.670 0.280 ;
        RECT  11.670 -0.280 11.950 0.800 ;
        RECT  10.860 -0.280 11.670 0.280 ;
        RECT  10.580 -0.280 10.860 0.340 ;
        RECT  8.220 -0.280 10.580 0.280 ;
        RECT  7.940 -0.280 8.220 0.340 ;
        RECT  6.540 -0.280 7.940 0.280 ;
        RECT  6.260 -0.280 6.540 0.340 ;
        RECT  5.440 -0.280 6.260 0.280 ;
        RECT  5.160 -0.280 5.440 0.340 ;
        RECT  3.760 -0.280 5.160 0.280 ;
        RECT  3.480 -0.280 3.760 0.800 ;
        RECT  2.580 -0.280 3.480 0.280 ;
        RECT  2.300 -0.280 2.580 0.340 ;
        RECT  0.890 -0.280 2.300 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.910 3.320 14.000 3.880 ;
        RECT  13.620 1.910 13.910 3.880 ;
        RECT  12.950 3.320 13.620 3.880 ;
        RECT  12.660 2.410 12.950 3.880 ;
        RECT  11.750 3.320 12.660 3.880 ;
        RECT  11.470 2.910 11.750 3.880 ;
        RECT  10.370 3.320 11.470 3.880 ;
        RECT  10.210 2.870 10.370 3.880 ;
        RECT  7.500 3.320 10.210 3.880 ;
        RECT  7.220 3.260 7.500 3.880 ;
        RECT  6.460 3.320 7.220 3.880 ;
        RECT  6.180 3.260 6.460 3.880 ;
        RECT  5.060 3.320 6.180 3.880 ;
        RECT  4.780 3.260 5.060 3.880 ;
        RECT  3.340 3.320 4.780 3.880 ;
        RECT  3.060 3.260 3.340 3.880 ;
        RECT  2.460 3.320 3.060 3.880 ;
        RECT  2.180 3.260 2.460 3.880 ;
        RECT  0.780 3.320 2.180 3.880 ;
        RECT  0.620 2.910 0.780 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.710 1.570 11.870 2.650 ;
        RECT  11.270 2.490 11.710 2.650 ;
        RECT  11.250 1.030 11.470 2.190 ;
        RECT  10.980 2.490 11.270 2.790 ;
        RECT  11.180 1.430 11.250 1.710 ;
        RECT  10.850 0.510 11.010 2.330 ;
        RECT  10.680 2.490 10.980 2.650 ;
        RECT  9.320 0.510 10.850 0.670 ;
        RECT  10.520 0.840 10.680 2.650 ;
        RECT  8.560 0.840 10.520 1.000 ;
        RECT  9.280 2.490 10.520 2.650 ;
        RECT  10.200 1.280 10.360 2.330 ;
        RECT  9.100 1.280 10.200 1.440 ;
        RECT  8.800 2.170 10.200 2.330 ;
        RECT  9.750 2.870 10.030 3.090 ;
        RECT  3.840 2.930 9.750 3.090 ;
        RECT  8.620 0.440 9.320 0.670 ;
        RECT  9.120 2.490 9.280 2.770 ;
        RECT  8.320 2.610 9.120 2.770 ;
        RECT  8.820 1.230 9.100 1.440 ;
        RECT  8.240 1.280 8.820 1.440 ;
        RECT  8.640 2.170 8.800 2.450 ;
        RECT  7.840 2.170 8.640 2.330 ;
        RECT  6.980 0.510 8.620 0.670 ;
        RECT  8.400 0.840 8.560 1.120 ;
        RECT  8.160 2.490 8.320 2.770 ;
        RECT  8.080 0.950 8.240 1.440 ;
        RECT  7.320 0.950 8.080 1.110 ;
        RECT  7.680 2.170 7.840 2.450 ;
        RECT  6.920 2.170 7.680 2.330 ;
        RECT  7.000 1.320 7.580 1.480 ;
        RECT  7.160 0.830 7.320 1.110 ;
        RECT  6.840 0.940 7.000 1.480 ;
        RECT  6.720 0.500 6.980 0.670 ;
        RECT  6.760 2.030 6.920 2.770 ;
        RECT  5.780 0.940 6.840 1.100 ;
        RECT  6.280 2.030 6.760 2.190 ;
        RECT  4.160 0.500 6.720 0.660 ;
        RECT  6.120 1.500 6.280 2.190 ;
        RECT  5.620 0.940 5.780 2.770 ;
        RECT  4.320 0.940 5.620 1.100 ;
        RECT  5.420 2.550 5.620 2.770 ;
        RECT  4.160 2.610 5.420 2.770 ;
        RECT  5.040 1.500 5.200 2.450 ;
        RECT  4.480 2.290 5.040 2.450 ;
        RECT  4.640 1.320 4.800 2.130 ;
        RECT  4.160 1.320 4.640 1.480 ;
        RECT  4.320 2.110 4.480 2.450 ;
        RECT  4.000 2.110 4.320 2.270 ;
        RECT  4.000 0.500 4.160 1.480 ;
        RECT  4.000 2.430 4.160 2.770 ;
        RECT  3.280 1.030 4.000 1.190 ;
        RECT  3.840 1.640 4.000 2.270 ;
        RECT  3.680 1.640 3.840 3.090 ;
        RECT  1.180 2.930 3.680 3.090 ;
        RECT  3.280 1.720 3.520 2.000 ;
        RECT  3.120 1.030 3.280 2.450 ;
        RECT  3.090 0.440 3.250 0.720 ;
        RECT  1.500 2.290 3.120 2.450 ;
        RECT  2.960 0.560 3.090 0.720 ;
        RECT  2.800 0.560 2.960 2.130 ;
        RECT  1.880 1.970 2.800 2.130 ;
        RECT  2.480 0.590 2.640 1.810 ;
        RECT  0.310 0.590 2.480 0.750 ;
        RECT  1.880 0.920 2.060 1.080 ;
        RECT  1.720 0.920 1.880 2.130 ;
        RECT  1.340 1.580 1.500 2.450 ;
        RECT  1.230 0.910 1.390 1.190 ;
        RECT  1.180 1.030 1.230 1.190 ;
        RECT  1.020 1.030 1.180 3.090 ;
        RECT  0.310 1.910 0.460 2.190 ;
        RECT  0.150 0.590 0.310 2.190 ;
    END
END DFFRHQX8TR

MACRO DFFRHQX4TR
    CLASS CORE ;
    FOREIGN DFFRHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.880 1.640 10.040 1.920 ;
        RECT  7.920 1.640 9.880 1.800 ;
        RECT  7.760 1.270 7.920 1.800 ;
        RECT  7.720 1.640 7.760 1.800 ;
        RECT  7.280 1.640 7.720 2.000 ;
        RECT  6.680 1.640 7.280 1.800 ;
        RECT  6.520 1.260 6.680 1.800 ;
        END
        ANTENNAGATEAREA 0.3888 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.240 0.470 12.520 3.160 ;
        RECT  12.080 1.440 12.240 2.160 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.240 2.320 1.640 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.840 1.730 ;
        END
        ANTENNAGATEAREA 0.348 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.940 -0.280 13.200 0.280 ;
        RECT  12.780 -0.280 12.940 1.310 ;
        RECT  12.000 -0.280 12.780 0.280 ;
        RECT  11.720 -0.280 12.000 0.800 ;
        RECT  10.860 -0.280 11.720 0.280 ;
        RECT  10.580 -0.280 10.860 0.340 ;
        RECT  8.220 -0.280 10.580 0.280 ;
        RECT  7.940 -0.280 8.220 0.340 ;
        RECT  6.540 -0.280 7.940 0.280 ;
        RECT  6.260 -0.280 6.540 0.340 ;
        RECT  5.440 -0.280 6.260 0.280 ;
        RECT  5.160 -0.280 5.440 0.340 ;
        RECT  3.760 -0.280 5.160 0.280 ;
        RECT  3.480 -0.280 3.760 0.800 ;
        RECT  2.580 -0.280 3.480 0.280 ;
        RECT  2.300 -0.280 2.580 0.340 ;
        RECT  0.890 -0.280 2.300 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.000 3.320 13.200 3.880 ;
        RECT  12.710 1.910 13.000 3.880 ;
        RECT  11.900 3.320 12.710 3.880 ;
        RECT  11.620 2.910 11.900 3.880 ;
        RECT  10.370 3.320 11.620 3.880 ;
        RECT  10.210 2.870 10.370 3.880 ;
        RECT  7.500 3.320 10.210 3.880 ;
        RECT  7.220 3.260 7.500 3.880 ;
        RECT  6.460 3.320 7.220 3.880 ;
        RECT  6.180 3.260 6.460 3.880 ;
        RECT  5.060 3.320 6.180 3.880 ;
        RECT  4.780 3.260 5.060 3.880 ;
        RECT  3.340 3.320 4.780 3.880 ;
        RECT  3.060 3.260 3.340 3.880 ;
        RECT  2.460 3.320 3.060 3.880 ;
        RECT  2.180 3.260 2.460 3.880 ;
        RECT  0.780 3.320 2.180 3.880 ;
        RECT  0.620 2.910 0.780 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.760 1.570 11.920 2.650 ;
        RECT  11.310 2.490 11.760 2.650 ;
        RECT  11.300 1.030 11.520 2.190 ;
        RECT  11.020 2.490 11.310 3.040 ;
        RECT  11.180 1.430 11.300 1.710 ;
        RECT  10.680 2.490 11.020 2.650 ;
        RECT  10.850 0.510 11.010 2.330 ;
        RECT  9.320 0.510 10.850 0.670 ;
        RECT  10.520 0.840 10.680 2.650 ;
        RECT  8.560 0.840 10.520 1.000 ;
        RECT  9.280 2.490 10.520 2.650 ;
        RECT  10.200 1.280 10.360 2.330 ;
        RECT  9.100 1.280 10.200 1.440 ;
        RECT  8.800 2.170 10.200 2.330 ;
        RECT  9.750 2.870 10.030 3.090 ;
        RECT  3.840 2.930 9.750 3.090 ;
        RECT  8.620 0.440 9.320 0.670 ;
        RECT  9.120 2.490 9.280 2.770 ;
        RECT  8.320 2.610 9.120 2.770 ;
        RECT  8.820 1.230 9.100 1.440 ;
        RECT  8.240 1.280 8.820 1.440 ;
        RECT  8.640 2.170 8.800 2.450 ;
        RECT  7.840 2.170 8.640 2.330 ;
        RECT  6.980 0.510 8.620 0.670 ;
        RECT  8.400 0.840 8.560 1.120 ;
        RECT  8.160 2.490 8.320 2.770 ;
        RECT  8.080 0.950 8.240 1.440 ;
        RECT  7.320 0.950 8.080 1.110 ;
        RECT  7.680 2.170 7.840 2.450 ;
        RECT  6.920 2.170 7.680 2.330 ;
        RECT  7.000 1.320 7.580 1.480 ;
        RECT  7.160 0.830 7.320 1.110 ;
        RECT  6.840 0.940 7.000 1.480 ;
        RECT  6.720 0.500 6.980 0.670 ;
        RECT  6.760 2.030 6.920 2.770 ;
        RECT  5.780 0.940 6.840 1.100 ;
        RECT  6.280 2.030 6.760 2.190 ;
        RECT  4.160 0.500 6.720 0.660 ;
        RECT  6.120 1.500 6.280 2.190 ;
        RECT  5.620 0.940 5.780 2.770 ;
        RECT  4.320 0.940 5.620 1.100 ;
        RECT  5.420 2.550 5.620 2.770 ;
        RECT  4.160 2.610 5.420 2.770 ;
        RECT  5.040 1.500 5.200 2.450 ;
        RECT  4.480 2.290 5.040 2.450 ;
        RECT  4.640 1.320 4.800 2.130 ;
        RECT  4.160 1.320 4.640 1.480 ;
        RECT  4.320 2.110 4.480 2.450 ;
        RECT  4.000 2.110 4.320 2.270 ;
        RECT  4.000 0.500 4.160 1.480 ;
        RECT  4.000 2.430 4.160 2.770 ;
        RECT  3.280 1.030 4.000 1.190 ;
        RECT  3.840 1.640 4.000 2.270 ;
        RECT  3.680 1.640 3.840 3.090 ;
        RECT  1.180 2.930 3.680 3.090 ;
        RECT  3.280 1.720 3.520 2.000 ;
        RECT  3.120 1.030 3.280 2.450 ;
        RECT  3.090 0.440 3.250 0.720 ;
        RECT  1.500 2.290 3.120 2.450 ;
        RECT  2.960 0.560 3.090 0.720 ;
        RECT  2.800 0.560 2.960 2.130 ;
        RECT  1.880 1.970 2.800 2.130 ;
        RECT  2.480 0.590 2.640 1.810 ;
        RECT  0.310 0.590 2.480 0.750 ;
        RECT  1.880 0.920 2.060 1.080 ;
        RECT  1.720 0.920 1.880 2.130 ;
        RECT  1.340 1.580 1.500 2.450 ;
        RECT  1.230 0.910 1.390 1.190 ;
        RECT  1.180 1.030 1.230 1.190 ;
        RECT  1.020 1.030 1.180 3.090 ;
        RECT  0.310 1.910 0.460 2.190 ;
        RECT  0.150 0.590 0.310 2.190 ;
    END
END DFFRHQX4TR

MACRO DFFRHQX2TR
    CLASS CORE ;
    FOREIGN DFFRHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.060 1.480 7.180 1.640 ;
        RECT  6.900 1.480 7.060 1.930 ;
        RECT  6.240 1.770 6.900 1.930 ;
        RECT  6.120 1.770 6.240 1.980 ;
        RECT  5.960 1.770 6.120 2.360 ;
        RECT  5.520 2.180 5.960 2.360 ;
        RECT  5.420 2.040 5.520 2.360 ;
        RECT  5.260 1.480 5.420 2.360 ;
        RECT  5.120 1.480 5.260 1.640 ;
        END
        ANTENNAGATEAREA 0.2376 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.800 2.040 9.920 3.160 ;
        RECT  9.640 0.440 9.800 3.160 ;
        END
        ANTENNADIFFAREA 3.885 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.240 2.730 1.560 ;
        END
        ANTENNAGATEAREA 0.0768 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.240 0.720 1.750 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.390 -0.280 10.000 0.280 ;
        RECT  9.100 -0.280 9.390 0.670 ;
        RECT  7.760 -0.280 9.100 0.280 ;
        RECT  7.480 -0.280 7.760 0.340 ;
        RECT  5.160 -0.280 7.480 0.280 ;
        RECT  4.880 -0.280 5.160 0.340 ;
        RECT  3.330 -0.280 4.880 0.280 ;
        RECT  2.530 -0.280 3.330 0.340 ;
        RECT  2.370 -0.280 2.530 1.080 ;
        RECT  0.000 -0.280 2.370 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.320 3.320 10.000 3.880 ;
        RECT  9.160 2.930 9.320 3.880 ;
        RECT  7.820 3.320 9.160 3.880 ;
        RECT  7.540 2.850 7.820 3.880 ;
        RECT  6.000 3.320 7.540 3.880 ;
        RECT  5.720 3.260 6.000 3.880 ;
        RECT  5.080 3.320 5.720 3.880 ;
        RECT  4.800 3.260 5.080 3.880 ;
        RECT  2.750 3.320 4.800 3.880 ;
        RECT  2.470 3.260 2.750 3.880 ;
        RECT  0.790 3.320 2.470 3.880 ;
        RECT  0.460 2.660 0.790 3.880 ;
        RECT  0.000 3.320 0.460 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.040 1.540 9.200 2.690 ;
        RECT  8.600 2.530 9.040 2.690 ;
        RECT  8.720 0.990 8.880 2.190 ;
        RECT  8.300 0.990 8.720 1.320 ;
        RECT  8.440 2.530 8.600 2.890 ;
        RECT  7.820 2.530 8.440 2.690 ;
        RECT  8.240 1.480 8.400 2.370 ;
        RECT  8.140 1.480 8.240 1.640 ;
        RECT  7.980 0.510 8.140 1.640 ;
        RECT  6.280 0.510 7.980 0.670 ;
        RECT  7.660 0.830 7.820 2.690 ;
        RECT  6.420 0.830 7.660 0.990 ;
        RECT  6.940 2.530 7.660 2.690 ;
        RECT  7.340 1.160 7.500 2.370 ;
        RECT  6.740 1.160 7.340 1.320 ;
        RECT  7.260 2.090 7.340 2.370 ;
        RECT  6.560 2.090 7.260 2.250 ;
        RECT  6.780 2.410 6.940 2.690 ;
        RECT  6.580 1.160 6.740 1.430 ;
        RECT  3.810 2.940 6.720 3.100 ;
        RECT  6.060 1.270 6.580 1.430 ;
        RECT  6.400 2.090 6.560 2.720 ;
        RECT  6.260 0.830 6.420 1.110 ;
        RECT  6.300 2.210 6.400 2.720 ;
        RECT  4.940 2.560 6.300 2.720 ;
        RECT  6.000 0.440 6.280 0.670 ;
        RECT  5.900 0.840 6.060 1.430 ;
        RECT  5.480 0.510 6.000 0.670 ;
        RECT  5.720 0.840 5.900 1.000 ;
        RECT  5.580 1.160 5.740 1.700 ;
        RECT  4.290 1.160 5.580 1.320 ;
        RECT  5.320 0.510 5.480 0.920 ;
        RECT  4.680 0.760 5.320 0.920 ;
        RECT  4.780 1.760 4.940 2.720 ;
        RECT  4.520 0.500 4.680 0.920 ;
        RECT  3.970 0.760 4.520 0.920 ;
        RECT  4.130 1.160 4.290 2.470 ;
        RECT  3.650 0.440 4.210 0.600 ;
        RECT  3.810 0.760 3.970 0.980 ;
        RECT  3.370 0.820 3.810 0.980 ;
        RECT  3.650 1.560 3.810 3.100 ;
        RECT  3.490 0.440 3.650 0.660 ;
        RECT  3.530 1.560 3.650 1.720 ;
        RECT  1.710 2.940 3.650 3.100 ;
        RECT  3.050 0.500 3.490 0.660 ;
        RECT  3.210 0.820 3.370 2.650 ;
        RECT  2.170 2.490 3.210 2.650 ;
        RECT  2.890 0.500 3.050 2.330 ;
        RECT  2.050 0.460 2.210 0.740 ;
        RECT  2.050 1.590 2.170 2.650 ;
        RECT  1.040 0.580 2.050 0.740 ;
        RECT  2.010 0.950 2.050 2.650 ;
        RECT  1.890 0.950 2.010 1.750 ;
        RECT  1.530 1.470 1.890 1.750 ;
        RECT  1.550 1.910 1.710 3.100 ;
        RECT  1.370 1.910 1.550 2.070 ;
        RECT  1.210 0.920 1.370 2.070 ;
        RECT  0.880 0.580 1.040 2.070 ;
        RECT  0.170 0.920 0.880 1.080 ;
        RECT  0.430 1.910 0.880 2.070 ;
        RECT  0.270 1.910 0.430 2.190 ;
    END
END DFFRHQX2TR

MACRO DFFRHQX1TR
    CLASS CORE ;
    FOREIGN DFFRHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.070 1.580 7.350 1.960 ;
        RECT  6.760 1.800 7.070 1.960 ;
        RECT  6.440 1.640 6.760 1.960 ;
        RECT  6.230 1.680 6.440 1.960 ;
        RECT  5.470 1.800 6.230 1.960 ;
        RECT  5.310 1.340 5.470 1.960 ;
        RECT  5.190 1.340 5.310 1.620 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.790 1.640 9.920 2.760 ;
        RECT  9.790 1.030 9.910 1.310 ;
        RECT  9.630 1.030 9.790 2.760 ;
        END
        ANTENNADIFFAREA 1.92 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.200 2.360 1.600 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.760 1.580 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.390 -0.280 10.000 0.280 ;
        RECT  9.110 -0.280 9.390 0.800 ;
        RECT  7.930 -0.280 9.110 0.340 ;
        RECT  7.650 -0.280 7.930 0.400 ;
        RECT  5.270 -0.280 7.650 0.340 ;
        RECT  4.990 -0.280 5.270 0.400 ;
        RECT  3.450 -0.280 4.990 0.340 ;
        RECT  2.080 -0.280 3.450 0.280 ;
        RECT  0.760 -0.280 2.080 0.340 ;
        RECT  0.000 -0.280 0.760 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.190 3.320 10.000 3.880 ;
        RECT  8.910 2.800 9.190 3.880 ;
        RECT  7.750 3.320 8.910 3.880 ;
        RECT  7.470 2.850 7.750 3.880 ;
        RECT  6.140 3.320 7.470 3.880 ;
        RECT  5.060 3.260 6.140 3.880 ;
        RECT  3.520 3.320 5.060 3.880 ;
        RECT  2.250 3.260 3.520 3.880 ;
        RECT  0.960 3.320 2.250 3.880 ;
        RECT  0.680 2.800 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.270 1.580 9.390 1.860 ;
        RECT  9.110 1.580 9.270 2.640 ;
        RECT  8.630 2.480 9.110 2.640 ;
        RECT  8.670 1.030 8.950 2.190 ;
        RECT  8.470 1.430 8.670 1.710 ;
        RECT  8.470 2.480 8.630 2.810 ;
        RECT  8.350 2.500 8.470 2.810 ;
        RECT  8.310 2.040 8.430 2.320 ;
        RECT  7.990 2.500 8.350 2.660 ;
        RECT  8.150 0.560 8.310 2.320 ;
        RECT  6.510 0.560 8.150 0.720 ;
        RECT  7.830 0.880 7.990 2.660 ;
        RECT  6.430 0.880 7.830 1.100 ;
        RECT  6.950 2.440 7.830 2.660 ;
        RECT  7.510 1.260 7.670 2.280 ;
        RECT  6.260 1.260 7.510 1.420 ;
        RECT  6.750 2.120 7.510 2.280 ;
        RECT  6.620 2.820 6.950 3.100 ;
        RECT  6.470 2.120 6.750 2.400 ;
        RECT  4.830 2.820 6.620 2.980 ;
        RECT  6.230 0.500 6.510 0.720 ;
        RECT  5.740 2.240 6.470 2.400 ;
        RECT  6.100 0.920 6.260 1.420 ;
        RECT  5.070 0.560 6.230 0.720 ;
        RECT  5.950 0.920 6.100 1.200 ;
        RECT  5.790 1.360 5.940 1.640 ;
        RECT  5.630 1.020 5.790 1.640 ;
        RECT  5.460 2.120 5.740 2.400 ;
        RECT  4.950 1.020 5.630 1.180 ;
        RECT  5.100 2.120 5.460 2.280 ;
        RECT  4.940 1.780 5.100 2.280 ;
        RECT  4.910 0.560 5.070 0.860 ;
        RECT  4.790 1.020 4.950 1.440 ;
        RECT  4.820 1.780 4.940 2.060 ;
        RECT  4.750 0.700 4.910 0.860 ;
        RECT  4.070 2.820 4.830 3.100 ;
        RECT  4.450 1.220 4.790 1.440 ;
        RECT  4.630 0.580 4.750 0.860 ;
        RECT  4.470 0.580 4.630 1.060 ;
        RECT  3.950 0.900 4.470 1.060 ;
        RECT  4.230 1.220 4.450 2.630 ;
        RECT  3.970 0.520 4.250 0.740 ;
        RECT  3.910 1.580 4.070 3.100 ;
        RECT  3.630 0.580 3.970 0.740 ;
        RECT  3.790 0.900 3.950 1.420 ;
        RECT  3.570 1.580 3.910 1.860 ;
        RECT  1.400 2.940 3.910 3.100 ;
        RECT  3.120 1.140 3.790 1.420 ;
        RECT  3.590 2.020 3.750 2.300 ;
        RECT  3.470 0.580 3.630 0.980 ;
        RECT  3.120 2.020 3.590 2.180 ;
        RECT  2.680 0.820 3.470 0.980 ;
        RECT  3.030 0.440 3.310 0.660 ;
        RECT  2.840 1.140 3.120 2.780 ;
        RECT  1.080 0.500 3.030 0.660 ;
        RECT  1.560 2.620 2.840 2.780 ;
        RECT  2.530 0.820 2.680 2.210 ;
        RECT  2.520 0.820 2.530 2.330 ;
        RECT  2.360 0.820 2.520 1.040 ;
        RECT  2.250 2.050 2.520 2.330 ;
        RECT  1.600 1.910 1.880 2.190 ;
        RECT  1.440 0.820 1.600 2.190 ;
        RECT  1.320 0.820 1.440 1.100 ;
        RECT  1.400 2.030 1.440 2.190 ;
        RECT  1.240 2.030 1.400 3.100 ;
        RECT  0.920 0.500 1.080 2.070 ;
        RECT  0.200 0.800 0.920 1.080 ;
        RECT  0.480 1.910 0.920 2.070 ;
        RECT  0.200 1.910 0.480 2.190 ;
    END
END DFFRHQX1TR

MACRO DFFRXLTR
    CLASS CORE ;
    FOREIGN DFFRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.470 6.050 1.520 ;
        RECT  4.810 0.470 5.890 0.630 ;
        RECT  4.650 0.470 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
        ANTENNAGATEAREA 0.1416 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.640 8.320 2.390 ;
        RECT  8.150 1.150 8.270 2.390 ;
        RECT  8.110 1.030 8.150 2.390 ;
        RECT  7.830 1.030 8.110 1.310 ;
        RECT  8.080 1.640 8.110 2.390 ;
        RECT  7.850 2.110 8.080 2.390 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.830 0.840 9.120 2.330 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.610 -0.280 9.200 0.280 ;
        RECT  8.330 -0.280 8.610 0.400 ;
        RECT  6.490 -0.280 8.330 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.580 3.320 9.200 3.880 ;
        RECT  7.290 3.200 8.580 3.880 ;
        RECT  6.080 3.320 7.290 3.880 ;
        RECT  5.800 3.200 6.080 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.640 2.600 8.920 2.880 ;
        RECT  7.010 2.680 8.640 2.880 ;
        RECT  7.670 1.670 7.730 1.950 ;
        RECT  7.670 0.450 7.710 0.670 ;
        RECT  7.650 0.450 7.670 1.950 ;
        RECT  7.510 0.450 7.650 2.520 ;
        RECT  7.430 0.450 7.510 0.670 ;
        RECT  7.490 1.410 7.510 2.520 ;
        RECT  7.370 2.240 7.490 2.520 ;
        RECT  7.010 1.030 7.350 1.310 ;
        RECT  6.850 1.030 7.010 3.160 ;
        RECT  6.290 1.900 6.850 2.060 ;
        RECT  6.260 2.940 6.850 3.160 ;
        RECT  6.470 2.500 6.690 2.780 ;
        RECT  5.730 2.500 6.470 2.660 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 0.790 5.730 2.880 ;
        RECT  5.450 0.790 5.570 1.070 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.970 0.790 5.190 1.830 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.970 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.660 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END DFFRXLTR

MACRO DFFRX4TR
    CLASS CORE ;
    FOREIGN DFFRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.110 1.360 6.430 1.520 ;
        RECT  5.950 0.440 6.110 1.520 ;
        RECT  4.810 0.440 5.950 0.600 ;
        RECT  4.650 0.440 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
        ANTENNAGATEAREA 0.2712 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.880 1.040 9.120 2.390 ;
        RECT  8.870 1.040 8.880 1.310 ;
        RECT  8.590 2.110 8.880 2.390 ;
        RECT  8.590 0.580 8.870 1.310 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.610 0.500 9.920 3.140 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
        ANTENNAGATEAREA 0.108 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.310 -0.280 10.400 0.280 ;
        RECT  10.090 -0.280 10.310 1.280 ;
        RECT  9.350 -0.280 10.090 0.280 ;
        RECT  9.070 -0.280 9.350 0.850 ;
        RECT  8.390 -0.280 9.070 0.280 ;
        RECT  8.110 -0.280 8.390 1.280 ;
        RECT  6.550 -0.280 8.110 0.280 ;
        RECT  6.270 -0.280 6.550 0.380 ;
        RECT  4.490 -0.280 6.270 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.310 3.320 10.400 3.880 ;
        RECT  10.090 2.060 10.310 3.880 ;
        RECT  9.350 3.320 10.090 3.880 ;
        RECT  9.070 2.990 9.350 3.880 ;
        RECT  8.390 3.320 9.070 3.880 ;
        RECT  8.110 2.990 8.390 3.880 ;
        RECT  7.380 3.320 8.110 3.880 ;
        RECT  7.100 3.260 7.380 3.880 ;
        RECT  6.250 3.320 7.100 3.880 ;
        RECT  5.890 2.750 6.250 3.880 ;
        RECT  3.670 3.320 5.890 3.880 ;
        RECT  3.390 2.470 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.290 1.590 9.450 2.710 ;
        RECT  7.820 2.550 9.290 2.710 ;
        RECT  7.950 1.670 8.050 1.950 ;
        RECT  7.790 0.450 7.950 2.350 ;
        RECT  7.660 2.550 7.820 2.940 ;
        RECT  7.610 0.450 7.790 0.780 ;
        RECT  7.650 1.670 7.790 2.350 ;
        RECT  7.450 2.780 7.660 2.940 ;
        RECT  7.290 0.530 7.450 2.940 ;
        RECT  7.130 0.530 7.290 1.310 ;
        RECT  6.110 1.900 7.290 2.060 ;
        RECT  6.770 2.780 7.290 2.940 ;
        RECT  5.730 2.320 6.950 2.480 ;
        RECT  6.490 2.660 6.770 2.940 ;
        RECT  5.890 1.780 6.110 2.060 ;
        RECT  5.570 0.980 5.730 2.880 ;
        RECT  5.470 0.980 5.570 1.260 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.970 0.930 5.190 1.830 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.970 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.660 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END DFFRX4TR

MACRO DFFRX2TR
    CLASS CORE ;
    FOREIGN DFFRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.610 6.050 1.520 ;
        RECT  4.810 0.610 5.890 0.770 ;
        RECT  4.650 0.610 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
        ANTENNAGATEAREA 0.1896 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.150 1.640 8.320 2.390 ;
        RECT  7.980 1.030 8.150 2.390 ;
        RECT  7.870 1.030 7.980 1.310 ;
        RECT  7.870 2.110 7.980 2.390 ;
        END
        ANTENNADIFFAREA 3.232 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.880 0.470 9.120 3.140 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.630 -0.280 9.200 0.280 ;
        RECT  8.350 -0.280 8.630 1.220 ;
        RECT  6.490 -0.280 8.350 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.630 3.320 9.200 3.880 ;
        RECT  8.350 2.990 8.630 3.880 ;
        RECT  7.380 3.320 8.350 3.880 ;
        RECT  7.100 3.260 7.380 3.880 ;
        RECT  6.250 3.320 7.100 3.880 ;
        RECT  5.800 3.200 6.250 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.560 1.590 8.720 2.710 ;
        RECT  7.230 2.550 8.560 2.710 ;
        RECT  7.670 0.450 7.810 0.670 ;
        RECT  7.690 1.670 7.760 1.950 ;
        RECT  7.670 1.670 7.690 2.350 ;
        RECT  7.510 0.450 7.670 2.350 ;
        RECT  7.410 2.070 7.510 2.350 ;
        RECT  7.230 1.030 7.350 1.250 ;
        RECT  7.070 1.030 7.230 2.710 ;
        RECT  6.290 1.900 7.070 2.060 ;
        RECT  6.490 2.430 7.070 2.710 ;
        RECT  6.660 2.870 6.940 3.140 ;
        RECT  5.730 2.870 6.660 3.030 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 1.020 5.730 3.030 ;
        RECT  5.450 1.020 5.570 1.310 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.890 1.170 5.170 1.830 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.890 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.590 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END DFFRX2TR

MACRO DFFRX1TR
    CLASS CORE ;
    FOREIGN DFFRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.470 6.050 1.520 ;
        RECT  4.810 0.470 5.890 0.630 ;
        RECT  4.650 0.470 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
        ANTENNAGATEAREA 0.1536 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.640 8.320 2.390 ;
        RECT  8.150 1.150 8.270 2.390 ;
        RECT  8.110 1.030 8.150 2.390 ;
        RECT  7.870 1.030 8.110 1.310 ;
        RECT  8.080 1.640 8.110 2.390 ;
        RECT  7.850 2.110 8.080 2.390 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.830 0.840 9.120 2.190 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.670 -0.280 9.200 0.280 ;
        RECT  8.390 -0.280 8.670 0.400 ;
        RECT  6.490 -0.280 8.390 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.580 3.320 9.200 3.880 ;
        RECT  7.290 3.200 8.580 3.880 ;
        RECT  6.080 3.320 7.290 3.880 ;
        RECT  5.800 3.200 6.080 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.640 2.600 8.920 2.880 ;
        RECT  7.010 2.680 8.640 2.880 ;
        RECT  7.670 1.670 7.730 1.950 ;
        RECT  7.670 0.450 7.710 0.670 ;
        RECT  7.650 0.450 7.670 1.950 ;
        RECT  7.510 0.450 7.650 2.520 ;
        RECT  7.430 0.450 7.510 0.670 ;
        RECT  7.490 1.410 7.510 2.520 ;
        RECT  7.370 2.240 7.490 2.520 ;
        RECT  7.010 1.030 7.350 1.250 ;
        RECT  6.850 1.030 7.010 3.160 ;
        RECT  6.290 1.900 6.850 2.060 ;
        RECT  6.260 2.940 6.850 3.160 ;
        RECT  6.470 2.500 6.690 2.780 ;
        RECT  5.730 2.500 6.470 2.660 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 0.790 5.730 2.880 ;
        RECT  5.450 0.790 5.570 1.070 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.970 0.790 5.190 1.830 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.970 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.660 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END DFFRX1TR

MACRO DFFQXLTR
    CLASS CORE ;
    FOREIGN DFFQXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.560 0.610 6.720 3.100 ;
        RECT  5.510 0.610 6.560 0.770 ;
        RECT  6.480 2.440 6.560 3.100 ;
        RECT  6.080 2.440 6.480 2.760 ;
        RECT  5.350 0.450 5.510 0.770 ;
        RECT  5.150 0.450 5.350 0.610 ;
        END
        ANTENNADIFFAREA 1.032 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 2.040 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.990 -0.280 6.800 0.280 ;
        RECT  5.710 -0.280 5.990 0.400 ;
        RECT  4.060 -0.280 5.710 0.280 ;
        RECT  3.900 -0.280 4.060 0.700 ;
        RECT  2.580 -0.280 3.900 0.280 ;
        RECT  1.860 -0.280 2.580 0.640 ;
        RECT  0.400 -0.280 1.860 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.220 3.320 6.800 3.880 ;
        RECT  5.940 2.920 6.220 3.880 ;
        RECT  4.140 3.320 5.940 3.880 ;
        RECT  3.850 3.260 4.140 3.880 ;
        RECT  2.920 3.320 3.850 3.880 ;
        RECT  2.640 3.260 2.920 3.880 ;
        RECT  1.940 3.320 2.640 3.880 ;
        RECT  1.660 3.260 1.940 3.880 ;
        RECT  0.400 3.320 1.660 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 1.030 6.400 2.230 ;
        RECT  6.120 1.800 6.240 2.230 ;
        RECT  5.670 1.800 6.120 1.960 ;
        RECT  5.890 1.350 6.050 1.640 ;
        RECT  5.180 1.350 5.890 1.510 ;
        RECT  5.390 1.680 5.670 1.960 ;
        RECT  5.020 1.030 5.180 3.160 ;
        RECT  4.850 1.030 5.020 1.310 ;
        RECT  4.830 0.570 4.990 0.870 ;
        RECT  4.700 1.660 4.860 2.990 ;
        RECT  4.690 0.710 4.830 0.870 ;
        RECT  4.690 1.660 4.700 1.940 ;
        RECT  2.340 2.830 4.700 2.990 ;
        RECT  4.530 0.710 4.690 1.940 ;
        RECT  4.380 2.110 4.540 2.670 ;
        RECT  4.110 1.660 4.530 1.940 ;
        RECT  3.950 2.110 4.380 2.270 ;
        RECT  3.240 2.510 4.380 2.670 ;
        RECT  4.190 1.000 4.350 1.310 ;
        RECT  3.950 1.150 4.190 1.310 ;
        RECT  3.790 1.150 3.950 2.270 ;
        RECT  3.470 0.690 3.630 2.270 ;
        RECT  3.410 0.690 3.470 0.850 ;
        RECT  3.250 0.440 3.410 0.850 ;
        RECT  3.240 1.110 3.310 1.880 ;
        RECT  2.910 0.440 3.250 0.600 ;
        RECT  3.150 1.110 3.240 2.670 ;
        RECT  3.080 1.720 3.150 2.670 ;
        RECT  1.770 1.720 3.080 1.880 ;
        RECT  1.160 1.400 2.990 1.560 ;
        RECT  1.660 1.020 2.470 1.180 ;
        RECT  2.180 2.520 2.340 2.990 ;
        RECT  1.360 2.830 2.180 2.990 ;
        RECT  1.610 1.720 1.770 2.000 ;
        RECT  1.500 0.590 1.660 1.180 ;
        RECT  0.800 0.590 1.500 0.750 ;
        RECT  1.200 2.830 1.360 3.110 ;
        RECT  0.800 2.830 1.200 2.990 ;
        RECT  1.130 1.400 1.160 2.670 ;
        RECT  1.000 0.930 1.130 2.670 ;
        RECT  0.970 0.930 1.000 1.560 ;
        RECT  0.640 0.590 0.800 2.990 ;
    END
END DFFQXLTR

MACRO DFFQX4TR
    CLASS CORE ;
    FOREIGN DFFQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.560 7.030 3.010 ;
        RECT  5.380 0.560 6.790 0.720 ;
        RECT  6.750 1.840 6.790 3.010 ;
        RECT  6.480 1.840 6.750 2.560 ;
        RECT  5.220 0.450 5.380 0.720 ;
        RECT  5.100 0.450 5.220 0.610 ;
        END
        ANTENNADIFFAREA 4.168 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 2.040 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.510 -0.280 7.600 0.280 ;
        RECT  7.230 -0.280 7.510 1.200 ;
        RECT  5.900 -0.280 7.230 0.280 ;
        RECT  5.620 -0.280 5.900 0.400 ;
        RECT  4.020 -0.280 5.620 0.280 ;
        RECT  3.860 -0.280 4.020 0.700 ;
        RECT  2.520 -0.280 3.860 0.280 ;
        RECT  1.860 -0.280 2.520 0.640 ;
        RECT  0.400 -0.280 1.860 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.510 3.320 7.600 3.880 ;
        RECT  7.230 2.020 7.510 3.880 ;
        RECT  6.290 3.320 7.230 3.880 ;
        RECT  5.600 2.920 6.290 3.880 ;
        RECT  4.030 3.320 5.600 3.880 ;
        RECT  3.740 3.260 4.030 3.880 ;
        RECT  2.820 3.320 3.740 3.880 ;
        RECT  2.540 3.260 2.820 3.880 ;
        RECT  1.840 3.320 2.540 3.880 ;
        RECT  1.560 3.260 1.840 3.880 ;
        RECT  0.400 3.320 1.560 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 1.420 6.630 1.580 ;
        RECT  6.080 1.030 6.240 2.230 ;
        RECT  5.960 1.910 6.080 2.230 ;
        RECT  5.580 1.910 5.960 2.070 ;
        RECT  5.760 1.360 5.920 1.640 ;
        RECT  5.070 1.360 5.760 1.520 ;
        RECT  5.300 1.680 5.580 2.070 ;
        RECT  4.910 1.030 5.070 3.160 ;
        RECT  4.780 0.590 4.940 0.870 ;
        RECT  4.770 1.030 4.910 1.310 ;
        RECT  4.610 0.710 4.780 0.870 ;
        RECT  4.610 1.660 4.750 2.990 ;
        RECT  4.590 0.710 4.610 2.990 ;
        RECT  4.450 0.710 4.590 1.940 ;
        RECT  2.240 2.830 4.590 2.990 ;
        RECT  4.110 1.660 4.450 1.940 ;
        RECT  4.270 2.110 4.430 2.670 ;
        RECT  4.130 1.000 4.290 1.310 ;
        RECT  3.950 2.110 4.270 2.270 ;
        RECT  3.100 2.510 4.270 2.670 ;
        RECT  3.950 1.150 4.130 1.310 ;
        RECT  3.790 1.150 3.950 2.270 ;
        RECT  3.470 0.690 3.630 2.210 ;
        RECT  3.370 0.690 3.470 0.850 ;
        RECT  3.350 2.050 3.470 2.210 ;
        RECT  3.210 0.440 3.370 0.850 ;
        RECT  3.120 1.110 3.280 1.880 ;
        RECT  2.870 0.440 3.210 0.600 ;
        RECT  3.100 1.720 3.120 1.880 ;
        RECT  2.940 1.720 3.100 2.670 ;
        RECT  1.770 1.720 2.940 1.880 ;
        RECT  1.100 1.400 2.890 1.560 ;
        RECT  1.630 1.020 2.440 1.180 ;
        RECT  2.080 2.520 2.240 2.990 ;
        RECT  1.260 2.830 2.080 2.990 ;
        RECT  1.580 1.720 1.770 2.000 ;
        RECT  1.470 0.590 1.630 1.180 ;
        RECT  0.730 0.590 1.470 0.750 ;
        RECT  1.100 2.830 1.260 3.110 ;
        RECT  1.060 0.930 1.100 1.560 ;
        RECT  0.730 2.830 1.100 2.990 ;
        RECT  0.900 0.930 1.060 2.670 ;
        RECT  0.570 0.590 0.730 2.990 ;
    END
END DFFQX4TR

MACRO DFFQX2TR
    CLASS CORE ;
    FOREIGN DFFQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.780 0.770 6.940 2.760 ;
        RECT  6.620 0.770 6.780 0.930 ;
        RECT  6.560 2.440 6.780 2.760 ;
        RECT  6.340 0.490 6.620 0.930 ;
        RECT  6.400 2.440 6.560 3.010 ;
        RECT  6.080 2.440 6.400 2.760 ;
        RECT  5.610 0.770 6.340 0.930 ;
        RECT  5.450 0.450 5.610 0.930 ;
        RECT  5.100 0.450 5.450 0.610 ;
        END
        ANTENNADIFFAREA 2.176 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 2.040 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.100 -0.280 7.200 0.280 ;
        RECT  6.820 -0.280 7.100 0.610 ;
        RECT  6.110 -0.280 6.820 0.280 ;
        RECT  5.830 -0.280 6.110 0.610 ;
        RECT  4.020 -0.280 5.830 0.280 ;
        RECT  3.860 -0.280 4.020 0.700 ;
        RECT  2.580 -0.280 3.860 0.280 ;
        RECT  1.860 -0.280 2.580 0.640 ;
        RECT  0.400 -0.280 1.860 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.100 3.320 7.200 3.880 ;
        RECT  6.820 2.920 7.100 3.880 ;
        RECT  6.140 3.320 6.820 3.880 ;
        RECT  5.860 2.920 6.140 3.880 ;
        RECT  4.140 3.320 5.860 3.880 ;
        RECT  3.850 3.260 4.140 3.880 ;
        RECT  2.920 3.320 3.850 3.880 ;
        RECT  2.640 3.260 2.920 3.880 ;
        RECT  1.940 3.320 2.640 3.880 ;
        RECT  1.660 3.260 1.940 3.880 ;
        RECT  0.400 3.320 1.660 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.450 1.090 6.610 2.170 ;
        RECT  6.120 1.090 6.450 1.250 ;
        RECT  5.640 2.010 6.450 2.170 ;
        RECT  5.820 1.360 5.980 1.640 ;
        RECT  5.180 1.360 5.820 1.520 ;
        RECT  5.360 1.680 5.640 2.170 ;
        RECT  5.020 1.030 5.180 3.160 ;
        RECT  4.770 1.030 5.020 1.310 ;
        RECT  4.780 0.570 4.940 0.870 ;
        RECT  4.700 1.660 4.860 2.990 ;
        RECT  4.610 0.710 4.780 0.870 ;
        RECT  4.610 1.660 4.700 1.940 ;
        RECT  2.340 2.830 4.700 2.990 ;
        RECT  4.450 0.710 4.610 1.940 ;
        RECT  4.380 2.110 4.540 2.670 ;
        RECT  4.110 1.660 4.450 1.940 ;
        RECT  3.950 2.110 4.380 2.270 ;
        RECT  3.240 2.510 4.380 2.670 ;
        RECT  4.130 1.000 4.290 1.310 ;
        RECT  3.950 1.150 4.130 1.310 ;
        RECT  3.790 1.150 3.950 2.270 ;
        RECT  3.470 0.690 3.630 2.270 ;
        RECT  3.370 0.690 3.470 0.850 ;
        RECT  3.210 0.440 3.370 0.850 ;
        RECT  3.240 1.110 3.310 1.880 ;
        RECT  3.150 1.110 3.240 2.670 ;
        RECT  2.870 0.440 3.210 0.600 ;
        RECT  3.080 1.720 3.150 2.670 ;
        RECT  1.770 1.720 3.080 1.880 ;
        RECT  1.160 1.400 2.990 1.560 ;
        RECT  1.660 1.020 2.470 1.180 ;
        RECT  2.180 2.520 2.340 2.990 ;
        RECT  1.360 2.830 2.180 2.990 ;
        RECT  1.610 1.720 1.770 2.000 ;
        RECT  1.500 0.590 1.660 1.180 ;
        RECT  0.800 0.590 1.500 0.750 ;
        RECT  1.200 2.830 1.360 3.110 ;
        RECT  0.800 2.830 1.200 2.990 ;
        RECT  1.130 1.400 1.160 2.670 ;
        RECT  1.000 0.930 1.130 2.670 ;
        RECT  0.970 0.930 1.000 1.560 ;
        RECT  0.640 0.590 0.800 2.990 ;
    END
END DFFQX2TR

MACRO DFFQX1TR
    CLASS CORE ;
    FOREIGN DFFQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.770 6.720 3.010 ;
        RECT  6.560 0.440 6.650 3.010 ;
        RECT  6.490 0.440 6.560 0.930 ;
        RECT  6.480 2.440 6.560 3.010 ;
        RECT  5.610 0.770 6.490 0.930 ;
        RECT  6.080 2.440 6.480 2.760 ;
        RECT  5.450 0.450 5.610 0.930 ;
        RECT  5.150 0.450 5.450 0.610 ;
        END
        ANTENNADIFFAREA 2.014 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.040 2.040 2.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.110 -0.280 6.800 0.280 ;
        RECT  5.830 -0.280 6.110 0.610 ;
        RECT  4.060 -0.280 5.830 0.280 ;
        RECT  3.900 -0.280 4.060 0.700 ;
        RECT  2.580 -0.280 3.900 0.280 ;
        RECT  1.860 -0.280 2.580 0.640 ;
        RECT  0.400 -0.280 1.860 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.220 3.320 6.800 3.880 ;
        RECT  5.940 2.920 6.220 3.880 ;
        RECT  4.140 3.320 5.940 3.880 ;
        RECT  3.850 3.260 4.140 3.880 ;
        RECT  2.920 3.320 3.850 3.880 ;
        RECT  2.640 3.260 2.920 3.880 ;
        RECT  1.940 3.320 2.640 3.880 ;
        RECT  1.660 3.260 1.940 3.880 ;
        RECT  0.400 3.320 1.660 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 1.090 6.400 2.230 ;
        RECT  6.120 1.090 6.240 1.250 ;
        RECT  6.120 1.800 6.240 2.230 ;
        RECT  5.640 1.800 6.120 1.960 ;
        RECT  5.820 1.350 5.980 1.640 ;
        RECT  5.180 1.350 5.820 1.510 ;
        RECT  5.380 1.680 5.640 1.960 ;
        RECT  5.020 1.030 5.180 3.160 ;
        RECT  4.850 1.030 5.020 1.310 ;
        RECT  4.830 0.570 4.990 0.870 ;
        RECT  4.700 1.660 4.860 2.990 ;
        RECT  4.690 0.710 4.830 0.870 ;
        RECT  4.690 1.660 4.700 1.940 ;
        RECT  2.340 2.830 4.700 2.990 ;
        RECT  4.530 0.710 4.690 1.940 ;
        RECT  4.380 2.110 4.540 2.670 ;
        RECT  4.110 1.660 4.530 1.940 ;
        RECT  3.950 2.110 4.380 2.270 ;
        RECT  3.240 2.510 4.380 2.670 ;
        RECT  4.190 1.000 4.350 1.310 ;
        RECT  3.950 1.150 4.190 1.310 ;
        RECT  3.790 1.150 3.950 2.270 ;
        RECT  3.470 0.690 3.630 2.270 ;
        RECT  3.410 0.690 3.470 0.850 ;
        RECT  3.250 0.440 3.410 0.850 ;
        RECT  3.240 1.110 3.310 1.880 ;
        RECT  2.910 0.440 3.250 0.600 ;
        RECT  3.150 1.110 3.240 2.670 ;
        RECT  3.080 1.720 3.150 2.670 ;
        RECT  1.770 1.720 3.080 1.880 ;
        RECT  1.160 1.400 2.990 1.560 ;
        RECT  1.660 1.020 2.470 1.180 ;
        RECT  2.180 2.520 2.340 2.990 ;
        RECT  1.360 2.830 2.180 2.990 ;
        RECT  1.610 1.720 1.770 2.000 ;
        RECT  1.500 0.590 1.660 1.180 ;
        RECT  0.800 0.590 1.500 0.750 ;
        RECT  1.200 2.830 1.360 3.110 ;
        RECT  0.800 2.830 1.200 2.990 ;
        RECT  1.130 1.400 1.160 2.670 ;
        RECT  1.000 0.930 1.130 2.670 ;
        RECT  0.970 0.930 1.000 1.560 ;
        RECT  0.640 0.590 0.800 2.990 ;
    END
END DFFQX1TR

MACRO DFFNSRXLTR
    CLASS CORE ;
    FOREIGN DFFNSRXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 2.440 7.520 2.800 ;
        RECT  6.970 2.520 7.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.470 3.230 1.750 ;
        RECT  2.880 1.240 3.120 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.030 9.520 2.360 ;
        END
        ANTENNADIFFAREA 1.1 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.440 2.040 8.720 2.360 ;
        RECT  8.280 1.030 8.440 2.360 ;
        END
        ANTENNADIFFAREA 1.1 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.470 2.720 1.960 ;
        RECT  2.440 1.470 2.480 1.640 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.070 -0.280 9.600 0.280 ;
        RECT  8.790 -0.280 9.070 0.340 ;
        RECT  7.660 -0.280 8.790 0.280 ;
        RECT  7.340 -0.280 7.660 0.400 ;
        RECT  3.530 -0.280 7.340 0.280 ;
        RECT  2.850 -0.280 3.530 0.290 ;
        RECT  1.890 -0.280 2.850 0.280 ;
        RECT  1.610 -0.280 1.890 0.290 ;
        RECT  0.000 -0.280 1.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.070 3.320 9.600 3.880 ;
        RECT  8.790 3.260 9.070 3.880 ;
        RECT  7.580 3.320 8.790 3.880 ;
        RECT  7.300 3.200 7.580 3.880 ;
        RECT  5.530 3.320 7.300 3.880 ;
        RECT  5.250 2.930 5.530 3.880 ;
        RECT  4.010 3.320 5.250 3.880 ;
        RECT  2.980 2.890 4.010 3.880 ;
        RECT  1.890 3.320 2.980 3.880 ;
        RECT  1.610 3.150 1.890 3.880 ;
        RECT  0.410 3.320 1.610 3.880 ;
        RECT  0.130 3.200 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.920 0.500 9.080 2.910 ;
        RECT  8.510 0.500 8.920 0.660 ;
        RECT  8.230 2.750 8.920 2.910 ;
        RECT  8.220 0.450 8.510 0.660 ;
        RECT  8.040 0.940 8.120 1.920 ;
        RECT  7.960 0.940 8.040 2.190 ;
        RECT  7.790 0.940 7.960 1.220 ;
        RECT  7.760 1.760 7.960 2.190 ;
        RECT  6.670 1.760 7.760 1.920 ;
        RECT  7.410 1.320 7.630 1.600 ;
        RECT  6.670 1.320 7.410 1.480 ;
        RECT  6.830 0.450 6.990 0.750 ;
        RECT  6.690 2.080 6.970 2.360 ;
        RECT  4.510 0.450 6.830 0.610 ;
        RECT  6.670 2.200 6.690 2.360 ;
        RECT  6.510 1.210 6.670 1.480 ;
        RECT  6.510 1.640 6.670 1.920 ;
        RECT  6.510 2.200 6.670 2.770 ;
        RECT  6.030 1.210 6.510 1.370 ;
        RECT  4.250 2.610 6.510 2.770 ;
        RECT  6.190 0.770 6.350 1.050 ;
        RECT  6.190 1.530 6.350 2.450 ;
        RECT  5.590 0.770 6.190 0.930 ;
        RECT  6.070 1.530 6.190 1.810 ;
        RECT  3.870 2.290 6.190 2.450 ;
        RECT  5.910 1.090 6.030 1.370 ;
        RECT  5.910 1.970 6.030 2.130 ;
        RECT  5.750 1.090 5.910 2.130 ;
        RECT  5.430 0.770 5.590 2.130 ;
        RECT  4.830 0.770 5.430 0.930 ;
        RECT  5.310 1.850 5.430 2.130 ;
        RECT  5.150 1.090 5.270 1.310 ;
        RECT  4.990 1.090 5.150 2.130 ;
        RECT  4.770 1.620 4.990 2.130 ;
        RECT  4.670 0.770 4.830 1.460 ;
        RECT  3.870 1.620 4.770 1.780 ;
        RECT  4.190 1.300 4.670 1.460 ;
        RECT  4.350 0.450 4.510 1.140 ;
        RECT  3.550 1.940 4.340 2.100 ;
        RECT  4.030 0.450 4.190 1.460 ;
        RECT  0.640 0.450 4.030 0.610 ;
        RECT  3.710 0.770 3.870 1.780 ;
        RECT  3.710 2.290 3.870 2.540 ;
        RECT  1.710 0.770 3.710 0.930 ;
        RECT  3.200 2.380 3.710 2.540 ;
        RECT  3.390 1.090 3.550 2.220 ;
        RECT  3.330 1.090 3.390 1.310 ;
        RECT  3.040 2.120 3.200 2.540 ;
        RECT  2.030 2.120 3.040 2.280 ;
        RECT  2.580 2.450 2.820 3.160 ;
        RECT  1.070 2.450 2.580 2.610 ;
        RECT  2.030 1.090 2.450 1.310 ;
        RECT  2.130 2.770 2.410 3.050 ;
        RECT  1.370 2.770 2.130 2.930 ;
        RECT  1.870 1.090 2.030 2.280 ;
        RECT  1.310 1.800 1.870 1.960 ;
        RECT  1.550 0.770 1.710 1.560 ;
        RECT  1.090 2.770 1.370 3.050 ;
        RECT  1.150 1.550 1.310 1.960 ;
        RECT  0.640 2.770 1.090 2.930 ;
        RECT  0.960 1.030 1.070 1.310 ;
        RECT  0.960 2.220 1.070 2.610 ;
        RECT  0.800 1.030 0.960 2.610 ;
        RECT  0.480 0.450 0.640 2.930 ;
    END
END DFFNSRXLTR

MACRO DFFNSRX4TR
    CLASS CORE ;
    FOREIGN DFFNSRX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.840 2.440 7.120 2.760 ;
        RECT  6.560 2.440 6.840 3.160 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.530 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.840 1.440 9.920 2.160 ;
        RECT  9.610 1.030 9.840 3.120 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.870 1.440 9.120 2.160 ;
        RECT  8.820 1.090 8.870 2.160 ;
        RECT  8.650 1.090 8.820 2.360 ;
        RECT  8.590 1.090 8.650 1.600 ;
        END
        ANTENNADIFFAREA 3.816 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.040 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 1.700 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.310 -0.280 10.400 0.280 ;
        RECT  10.030 -0.280 10.310 1.150 ;
        RECT  9.350 -0.280 10.030 0.280 ;
        RECT  9.070 -0.280 9.350 0.610 ;
        RECT  8.390 -0.280 9.070 0.280 ;
        RECT  8.110 -0.280 8.390 0.610 ;
        RECT  7.450 -0.280 8.110 0.280 ;
        RECT  7.170 -0.280 7.450 0.400 ;
        RECT  3.420 -0.280 7.170 0.280 ;
        RECT  2.740 -0.280 3.420 0.290 ;
        RECT  1.780 -0.280 2.740 0.280 ;
        RECT  1.500 -0.280 1.780 0.290 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.310 3.320 10.400 3.880 ;
        RECT  10.030 2.510 10.310 3.880 ;
        RECT  9.350 3.320 10.030 3.880 ;
        RECT  9.070 2.850 9.350 3.880 ;
        RECT  8.390 3.320 9.070 3.880 ;
        RECT  8.110 2.850 8.390 3.880 ;
        RECT  7.280 3.320 8.110 3.880 ;
        RECT  7.000 3.200 7.280 3.880 ;
        RECT  5.420 3.320 7.000 3.880 ;
        RECT  5.140 2.990 5.420 3.880 ;
        RECT  3.900 3.320 5.140 3.880 ;
        RECT  2.930 2.890 3.900 3.880 ;
        RECT  1.780 3.320 2.930 3.880 ;
        RECT  1.500 3.150 1.780 3.880 ;
        RECT  0.370 3.320 1.500 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.280 0.770 9.440 2.680 ;
        RECT  7.910 0.770 9.280 0.930 ;
        RECT  7.910 2.520 9.280 2.680 ;
        RECT  8.270 1.090 8.430 2.170 ;
        RECT  7.570 1.090 8.270 1.310 ;
        RECT  7.690 2.010 8.270 2.170 ;
        RECT  7.630 0.450 7.910 0.930 ;
        RECT  7.750 2.520 7.910 3.150 ;
        RECT  7.630 2.940 7.750 3.150 ;
        RECT  7.410 2.010 7.690 2.330 ;
        RECT  6.930 1.550 7.580 1.830 ;
        RECT  6.560 2.010 7.410 2.170 ;
        RECT  6.760 1.320 6.930 1.830 ;
        RECT  6.630 0.450 6.910 0.750 ;
        RECT  6.560 1.320 6.760 1.480 ;
        RECT  4.400 0.450 6.630 0.610 ;
        RECT  6.400 1.210 6.560 1.480 ;
        RECT  6.400 1.640 6.560 2.170 ;
        RECT  5.860 1.210 6.400 1.370 ;
        RECT  4.420 2.670 6.400 2.830 ;
        RECT  6.080 1.530 6.240 2.510 ;
        RECT  6.050 0.770 6.210 1.050 ;
        RECT  5.960 1.530 6.080 1.810 ;
        RECT  4.740 2.350 6.080 2.510 ;
        RECT  5.480 0.770 6.050 0.930 ;
        RECT  5.800 1.970 5.920 2.190 ;
        RECT  5.800 1.090 5.860 1.370 ;
        RECT  5.640 1.090 5.800 2.190 ;
        RECT  5.320 0.770 5.480 2.050 ;
        RECT  4.720 0.770 5.320 0.930 ;
        RECT  5.200 1.770 5.320 2.050 ;
        RECT  5.040 1.090 5.160 1.310 ;
        RECT  4.940 1.090 5.040 1.780 ;
        RECT  4.880 1.090 4.940 2.130 ;
        RECT  4.660 1.620 4.880 2.130 ;
        RECT  4.580 2.290 4.740 2.510 ;
        RECT  4.560 0.770 4.720 1.460 ;
        RECT  3.760 1.620 4.660 1.780 ;
        RECT  3.820 2.290 4.580 2.450 ;
        RECT  4.080 1.300 4.560 1.460 ;
        RECT  4.140 2.610 4.420 2.830 ;
        RECT  4.240 0.450 4.400 1.140 ;
        RECT  3.500 1.940 4.230 2.100 ;
        RECT  3.920 0.450 4.080 1.460 ;
        RECT  0.720 0.450 3.920 0.610 ;
        RECT  3.660 2.290 3.820 2.570 ;
        RECT  3.600 0.770 3.760 1.780 ;
        RECT  3.090 2.410 3.660 2.570 ;
        RECT  1.680 0.770 3.600 0.930 ;
        RECT  3.440 1.940 3.500 2.250 ;
        RECT  3.280 1.090 3.440 2.250 ;
        RECT  2.930 2.120 3.090 2.570 ;
        RECT  2.320 2.120 2.930 2.280 ;
        RECT  2.530 2.450 2.770 3.160 ;
        RECT  1.040 2.450 2.530 2.610 ;
        RECT  2.090 2.770 2.370 3.050 ;
        RECT  2.100 1.140 2.320 2.280 ;
        RECT  1.360 2.120 2.100 2.280 ;
        RECT  1.330 2.770 2.090 2.930 ;
        RECT  1.520 0.770 1.680 1.960 ;
        RECT  1.200 1.280 1.360 2.280 ;
        RECT  1.050 2.770 1.330 3.050 ;
        RECT  1.040 0.780 1.180 1.060 ;
        RECT  0.720 2.770 1.050 2.930 ;
        RECT  0.880 0.780 1.040 2.610 ;
        RECT  0.560 0.450 0.720 2.930 ;
    END
END DFFNSRX4TR

MACRO DFFNSRX2TR
    CLASS CORE ;
    FOREIGN DFFNSRX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 2.440 7.520 2.800 ;
        RECT  6.860 2.520 7.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.530 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 0.610 9.520 2.730 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.420 2.040 8.720 2.720 ;
        RECT  8.420 1.090 8.550 1.310 ;
        RECT  8.250 1.090 8.420 2.720 ;
        END
        ANTENNADIFFAREA 3.386 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.040 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 1.700 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.030 -0.280 9.600 0.280 ;
        RECT  8.750 -0.280 9.030 0.610 ;
        RECT  7.540 -0.280 8.750 0.280 ;
        RECT  7.260 -0.280 7.540 0.400 ;
        RECT  3.420 -0.280 7.260 0.280 ;
        RECT  2.740 -0.280 3.420 0.290 ;
        RECT  1.780 -0.280 2.740 0.280 ;
        RECT  1.500 -0.280 1.780 0.290 ;
        RECT  0.000 -0.280 1.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.990 3.320 9.600 3.880 ;
        RECT  8.710 3.260 8.990 3.880 ;
        RECT  7.460 3.320 8.710 3.880 ;
        RECT  7.180 3.200 7.460 3.880 ;
        RECT  5.420 3.320 7.180 3.880 ;
        RECT  5.140 2.990 5.420 3.880 ;
        RECT  3.900 3.320 5.140 3.880 ;
        RECT  2.930 2.890 3.900 3.880 ;
        RECT  1.780 3.320 2.930 3.880 ;
        RECT  1.500 3.150 1.780 3.880 ;
        RECT  0.370 3.320 1.500 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.960 0.770 9.120 3.100 ;
        RECT  8.210 0.770 8.960 0.930 ;
        RECT  8.900 1.350 8.960 1.640 ;
        RECT  7.980 2.940 8.960 3.100 ;
        RECT  7.930 0.450 8.210 0.930 ;
        RECT  7.930 1.090 8.090 1.950 ;
        RECT  7.700 2.940 7.980 3.150 ;
        RECT  7.640 1.090 7.930 1.310 ;
        RECT  7.920 1.790 7.930 1.950 ;
        RECT  7.760 1.790 7.920 2.190 ;
        RECT  6.560 1.790 7.760 1.950 ;
        RECT  6.930 1.470 7.580 1.630 ;
        RECT  6.760 1.210 6.930 1.630 ;
        RECT  6.630 0.450 6.910 0.750 ;
        RECT  6.580 2.110 6.860 2.360 ;
        RECT  5.860 1.210 6.760 1.370 ;
        RECT  4.400 0.450 6.630 0.610 ;
        RECT  6.560 2.200 6.580 2.360 ;
        RECT  6.400 1.640 6.560 1.950 ;
        RECT  6.400 2.200 6.560 2.830 ;
        RECT  4.420 2.670 6.400 2.830 ;
        RECT  6.080 1.530 6.240 2.510 ;
        RECT  6.050 0.770 6.210 1.050 ;
        RECT  5.960 1.530 6.080 1.810 ;
        RECT  4.740 2.350 6.080 2.510 ;
        RECT  5.480 0.770 6.050 0.930 ;
        RECT  5.800 1.970 5.920 2.190 ;
        RECT  5.800 1.090 5.860 1.370 ;
        RECT  5.640 1.090 5.800 2.190 ;
        RECT  5.320 0.770 5.480 2.190 ;
        RECT  4.720 0.770 5.320 0.930 ;
        RECT  5.200 1.910 5.320 2.190 ;
        RECT  5.040 1.090 5.160 1.310 ;
        RECT  4.880 1.090 5.040 2.130 ;
        RECT  4.660 1.620 4.880 2.130 ;
        RECT  4.580 2.290 4.740 2.510 ;
        RECT  4.560 0.770 4.720 1.460 ;
        RECT  3.760 1.620 4.660 1.780 ;
        RECT  3.820 2.290 4.580 2.450 ;
        RECT  4.080 1.300 4.560 1.460 ;
        RECT  4.140 2.610 4.420 2.830 ;
        RECT  4.240 0.450 4.400 1.140 ;
        RECT  3.500 1.940 4.230 2.100 ;
        RECT  3.920 0.450 4.080 1.460 ;
        RECT  0.720 0.450 3.920 0.610 ;
        RECT  3.660 2.290 3.820 2.570 ;
        RECT  3.600 0.770 3.760 1.780 ;
        RECT  3.090 2.410 3.660 2.570 ;
        RECT  1.680 0.770 3.600 0.930 ;
        RECT  3.440 1.940 3.500 2.250 ;
        RECT  3.280 1.090 3.440 2.250 ;
        RECT  2.930 2.120 3.090 2.570 ;
        RECT  2.320 2.120 2.930 2.280 ;
        RECT  2.530 2.450 2.770 3.160 ;
        RECT  1.040 2.450 2.530 2.610 ;
        RECT  2.090 2.770 2.370 3.050 ;
        RECT  2.100 1.140 2.320 2.280 ;
        RECT  1.360 2.120 2.100 2.280 ;
        RECT  1.330 2.770 2.090 2.930 ;
        RECT  1.520 0.770 1.680 1.960 ;
        RECT  1.200 1.280 1.360 2.280 ;
        RECT  1.050 2.770 1.330 3.050 ;
        RECT  1.040 0.780 1.180 1.060 ;
        RECT  0.720 2.770 1.050 2.930 ;
        RECT  0.880 0.780 1.040 2.610 ;
        RECT  0.560 0.450 0.720 2.930 ;
    END
END DFFNSRX2TR

MACRO DFFNSRX1TR
    CLASS CORE ;
    FOREIGN DFFNSRX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 2.440 7.520 2.800 ;
        RECT  6.970 2.520 7.280 2.800 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.470 3.230 1.750 ;
        RECT  2.880 1.240 3.120 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.030 9.520 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.520 2.040 8.720 2.360 ;
        RECT  8.360 1.030 8.520 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.470 2.720 1.960 ;
        RECT  2.440 1.470 2.480 1.640 ;
        END
        ANTENNAGATEAREA 0.0864 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 -0.280 9.600 0.280 ;
        RECT  8.830 -0.280 9.110 0.340 ;
        RECT  7.580 -0.280 8.830 0.280 ;
        RECT  7.300 -0.280 7.580 0.800 ;
        RECT  3.530 -0.280 7.300 0.280 ;
        RECT  2.850 -0.280 3.530 0.290 ;
        RECT  1.890 -0.280 2.850 0.280 ;
        RECT  1.610 -0.280 1.890 0.290 ;
        RECT  0.000 -0.280 1.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.110 3.320 9.600 3.880 ;
        RECT  8.830 3.260 9.110 3.880 ;
        RECT  7.570 3.320 8.830 3.880 ;
        RECT  7.290 3.200 7.570 3.880 ;
        RECT  5.530 3.320 7.290 3.880 ;
        RECT  5.250 2.930 5.530 3.880 ;
        RECT  4.010 3.320 5.250 3.880 ;
        RECT  2.980 2.890 4.010 3.880 ;
        RECT  1.890 3.320 2.980 3.880 ;
        RECT  1.610 3.150 1.890 3.880 ;
        RECT  0.410 3.320 1.610 3.880 ;
        RECT  0.130 3.200 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.120 2.910 9.130 3.070 ;
        RECT  8.960 0.500 9.120 3.070 ;
        RECT  8.440 0.500 8.960 0.660 ;
        RECT  7.810 2.910 8.960 3.070 ;
        RECT  8.160 0.450 8.440 0.660 ;
        RECT  8.030 1.000 8.140 1.920 ;
        RECT  7.980 1.000 8.030 2.190 ;
        RECT  7.840 1.000 7.980 1.160 ;
        RECT  7.870 1.760 7.980 2.190 ;
        RECT  6.670 1.760 7.870 1.920 ;
        RECT  7.520 1.320 7.740 1.600 ;
        RECT  6.670 1.320 7.520 1.480 ;
        RECT  6.930 0.470 6.990 0.750 ;
        RECT  6.690 2.080 6.970 2.360 ;
        RECT  6.830 0.450 6.930 0.750 ;
        RECT  4.510 0.450 6.830 0.610 ;
        RECT  6.670 2.200 6.690 2.360 ;
        RECT  6.510 1.210 6.670 1.480 ;
        RECT  6.510 1.640 6.670 1.920 ;
        RECT  6.510 2.200 6.670 2.770 ;
        RECT  6.030 1.210 6.510 1.370 ;
        RECT  4.250 2.610 6.510 2.770 ;
        RECT  6.190 0.770 6.350 1.050 ;
        RECT  6.190 1.530 6.350 2.450 ;
        RECT  5.590 0.770 6.190 0.930 ;
        RECT  6.070 1.530 6.190 1.810 ;
        RECT  3.870 2.290 6.190 2.450 ;
        RECT  5.910 1.090 6.030 1.370 ;
        RECT  5.910 1.970 6.030 2.130 ;
        RECT  5.750 1.090 5.910 2.130 ;
        RECT  5.430 0.770 5.590 2.130 ;
        RECT  4.830 0.770 5.430 0.930 ;
        RECT  5.310 1.850 5.430 2.130 ;
        RECT  5.150 1.090 5.270 1.310 ;
        RECT  4.990 1.090 5.150 2.130 ;
        RECT  4.770 1.620 4.990 2.130 ;
        RECT  4.670 0.770 4.830 1.460 ;
        RECT  3.870 1.620 4.770 1.780 ;
        RECT  4.190 1.300 4.670 1.460 ;
        RECT  4.350 0.450 4.510 1.140 ;
        RECT  3.550 1.940 4.340 2.100 ;
        RECT  4.030 0.450 4.190 1.460 ;
        RECT  0.640 0.450 4.030 0.610 ;
        RECT  3.710 0.770 3.870 1.780 ;
        RECT  3.710 2.290 3.870 2.540 ;
        RECT  1.710 0.770 3.710 0.930 ;
        RECT  3.200 2.380 3.710 2.540 ;
        RECT  3.390 1.090 3.550 2.220 ;
        RECT  3.280 1.090 3.390 1.310 ;
        RECT  3.040 2.120 3.200 2.540 ;
        RECT  2.030 2.120 3.040 2.280 ;
        RECT  2.580 2.450 2.820 3.160 ;
        RECT  1.070 2.450 2.580 2.610 ;
        RECT  2.030 1.090 2.450 1.310 ;
        RECT  2.130 2.770 2.410 3.050 ;
        RECT  1.370 2.770 2.130 2.930 ;
        RECT  1.870 1.090 2.030 2.280 ;
        RECT  1.310 1.800 1.870 1.960 ;
        RECT  1.550 0.770 1.710 1.560 ;
        RECT  1.090 2.770 1.370 3.050 ;
        RECT  1.150 1.550 1.310 1.960 ;
        RECT  0.640 2.770 1.090 2.930 ;
        RECT  0.960 1.030 1.070 1.310 ;
        RECT  0.960 2.220 1.070 2.610 ;
        RECT  0.800 1.030 0.960 2.610 ;
        RECT  0.480 0.450 0.640 2.930 ;
    END
END DFFNSRX1TR

MACRO DFFHQX8TR
    CLASS CORE ;
    FOREIGN DFFHQX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.750 0.620 13.030 3.030 ;
        RECT  12.070 1.470 12.750 1.940 ;
        RECT  11.800 0.630 12.070 2.990 ;
        RECT  11.790 1.440 11.800 2.990 ;
        RECT  11.330 1.440 11.790 1.930 ;
        RECT  11.130 1.440 11.330 2.160 ;
        RECT  11.120 1.440 11.130 2.990 ;
        RECT  10.820 0.630 11.120 2.990 ;
        RECT  10.810 1.430 10.820 2.990 ;
        RECT  10.680 1.430 10.810 2.160 ;
        END
        ANTENNADIFFAREA 9.984 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.580 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.160 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.3432 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.560 -0.280 13.200 0.280 ;
        RECT  12.270 -0.280 12.560 1.190 ;
        RECT  11.610 -0.280 12.270 0.280 ;
        RECT  11.310 -0.280 11.610 1.200 ;
        RECT  10.600 -0.280 11.310 0.280 ;
        RECT  10.300 -0.280 10.600 0.800 ;
        RECT  6.340 -0.280 10.300 0.280 ;
        RECT  6.060 -0.280 6.340 0.340 ;
        RECT  5.300 -0.280 6.060 0.280 ;
        RECT  5.020 -0.280 5.300 0.340 ;
        RECT  3.700 -0.280 5.020 0.280 ;
        RECT  3.540 -0.280 3.700 1.050 ;
        RECT  2.340 -0.280 3.540 0.280 ;
        RECT  3.220 0.770 3.540 1.050 ;
        RECT  2.180 -0.280 2.340 0.870 ;
        RECT  0.780 -0.280 2.180 0.280 ;
        RECT  0.500 -0.280 0.780 0.340 ;
        RECT  0.000 -0.280 0.500 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.550 3.320 13.200 3.880 ;
        RECT  12.270 2.130 12.550 3.880 ;
        RECT  11.590 3.320 12.270 3.880 ;
        RECT  11.310 2.470 11.590 3.880 ;
        RECT  10.630 3.320 11.310 3.880 ;
        RECT  9.970 2.700 10.630 3.880 ;
        RECT  7.380 3.320 9.970 3.880 ;
        RECT  7.100 3.260 7.380 3.880 ;
        RECT  6.340 3.320 7.100 3.880 ;
        RECT  6.060 3.260 6.340 3.880 ;
        RECT  4.660 3.320 6.060 3.880 ;
        RECT  4.380 3.260 4.660 3.880 ;
        RECT  3.400 3.320 4.380 3.880 ;
        RECT  3.120 3.260 3.400 3.880 ;
        RECT  2.360 3.320 3.120 3.880 ;
        RECT  2.080 3.260 2.360 3.880 ;
        RECT  0.780 3.320 2.080 3.880 ;
        RECT  0.500 3.260 0.780 3.880 ;
        RECT  0.000 3.320 0.500 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.290 1.480 10.450 2.530 ;
        RECT  9.810 2.370 10.290 2.530 ;
        RECT  9.970 1.030 10.130 2.190 ;
        RECT  9.710 1.490 9.970 1.650 ;
        RECT  9.650 2.370 9.810 2.840 ;
        RECT  9.110 2.680 9.650 2.840 ;
        RECT  9.490 0.440 9.550 1.790 ;
        RECT  9.390 0.440 9.490 2.510 ;
        RECT  7.540 0.440 9.390 0.600 ;
        RECT  9.330 1.610 9.390 2.510 ;
        RECT  9.070 0.760 9.230 1.240 ;
        RECT  8.950 1.900 9.110 2.840 ;
        RECT  8.230 1.080 9.070 1.240 ;
        RECT  8.350 1.900 8.950 2.060 ;
        RECT  7.910 0.760 8.830 0.920 ;
        RECT  8.550 2.220 8.790 2.960 ;
        RECT  7.910 2.800 8.550 2.960 ;
        RECT  8.230 1.900 8.350 2.640 ;
        RECT  8.070 1.080 8.230 2.640 ;
        RECT  7.750 0.760 7.910 2.960 ;
        RECT  7.650 1.020 7.750 1.300 ;
        RECT  7.590 1.930 7.750 2.580 ;
        RECT  6.800 1.140 7.650 1.300 ;
        RECT  6.800 1.930 7.590 2.090 ;
        RECT  7.430 2.760 7.590 3.040 ;
        RECT  7.380 0.440 7.540 0.720 ;
        RECT  3.440 2.880 7.430 3.040 ;
        RECT  5.800 0.560 7.380 0.720 ;
        RECT  6.440 1.460 7.060 1.620 ;
        RECT  6.640 1.020 6.800 1.300 ;
        RECT  6.640 1.930 6.800 2.610 ;
        RECT  6.120 1.930 6.640 2.090 ;
        RECT  6.280 0.880 6.440 1.620 ;
        RECT  5.080 0.880 6.280 1.040 ;
        RECT  5.960 1.600 6.120 2.090 ;
        RECT  5.640 0.440 5.800 0.720 ;
        RECT  4.020 0.560 5.640 0.720 ;
        RECT  5.080 2.260 5.500 2.420 ;
        RECT  4.920 0.880 5.080 2.420 ;
        RECT  4.180 0.880 4.920 1.040 ;
        RECT  3.760 2.260 4.920 2.420 ;
        RECT  4.200 1.810 4.760 2.090 ;
        RECT  4.020 1.810 4.200 1.970 ;
        RECT  3.860 0.560 4.020 1.970 ;
        RECT  2.980 1.210 3.860 1.370 ;
        RECT  3.600 2.140 3.760 2.420 ;
        RECT  3.440 1.530 3.700 1.690 ;
        RECT  3.280 1.530 3.440 3.040 ;
        RECT  2.660 0.440 3.380 0.600 ;
        RECT  1.560 2.880 3.280 3.040 ;
        RECT  2.820 1.030 2.980 2.720 ;
        RECT  2.660 2.440 2.820 2.720 ;
        RECT  2.500 0.440 2.660 1.190 ;
        RECT  1.360 2.560 2.660 2.720 ;
        RECT  1.820 1.030 2.500 1.190 ;
        RECT  1.820 2.120 1.900 2.400 ;
        RECT  1.660 1.030 1.820 2.400 ;
        RECT  1.540 0.440 1.700 0.720 ;
        RECT  1.400 2.880 1.560 3.160 ;
        RECT  0.320 0.560 1.540 0.720 ;
        RECT  1.040 2.880 1.400 3.040 ;
        RECT  1.200 1.580 1.360 2.720 ;
        RECT  1.040 1.090 1.300 1.250 ;
        RECT  0.880 1.090 1.040 3.040 ;
        RECT  0.160 0.560 0.320 2.190 ;
    END
END DFFHQX8TR

MACRO DFFHQX4TR
    CLASS CORE ;
    FOREIGN DFFHQX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.040 1.430 11.160 2.180 ;
        RECT  10.720 0.630 11.040 2.990 ;
        END
        ANTENNADIFFAREA 3.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 1.580 2.330 1.960 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.160 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.3432 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.500 -0.280 11.600 0.280 ;
        RECT  11.220 -0.280 11.500 1.200 ;
        RECT  10.510 -0.280 11.220 0.280 ;
        RECT  10.210 -0.280 10.510 0.800 ;
        RECT  6.250 -0.280 10.210 0.280 ;
        RECT  5.970 -0.280 6.250 0.340 ;
        RECT  5.210 -0.280 5.970 0.280 ;
        RECT  4.930 -0.280 5.210 0.340 ;
        RECT  3.610 -0.280 4.930 0.280 ;
        RECT  3.450 -0.280 3.610 1.050 ;
        RECT  2.250 -0.280 3.450 0.280 ;
        RECT  3.130 0.770 3.450 1.050 ;
        RECT  2.090 -0.280 2.250 0.870 ;
        RECT  0.770 -0.280 2.090 0.280 ;
        RECT  0.490 -0.280 0.770 0.340 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.510 3.320 11.600 3.880 ;
        RECT  11.220 2.470 11.510 3.880 ;
        RECT  10.540 3.320 11.220 3.880 ;
        RECT  9.880 2.700 10.540 3.880 ;
        RECT  7.290 3.320 9.880 3.880 ;
        RECT  7.010 3.260 7.290 3.880 ;
        RECT  6.250 3.320 7.010 3.880 ;
        RECT  5.970 3.260 6.250 3.880 ;
        RECT  4.570 3.320 5.970 3.880 ;
        RECT  4.290 3.260 4.570 3.880 ;
        RECT  3.390 3.320 4.290 3.880 ;
        RECT  3.110 3.260 3.390 3.880 ;
        RECT  2.350 3.320 3.110 3.880 ;
        RECT  2.070 3.260 2.350 3.880 ;
        RECT  0.770 3.320 2.070 3.880 ;
        RECT  0.490 3.260 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.200 1.480 10.360 2.530 ;
        RECT  9.720 2.370 10.200 2.530 ;
        RECT  9.880 1.030 10.040 2.190 ;
        RECT  9.620 1.490 9.880 1.650 ;
        RECT  9.560 2.370 9.720 2.840 ;
        RECT  9.020 2.680 9.560 2.840 ;
        RECT  9.400 0.440 9.460 1.790 ;
        RECT  9.300 0.440 9.400 2.510 ;
        RECT  7.450 0.440 9.300 0.600 ;
        RECT  9.240 1.610 9.300 2.510 ;
        RECT  8.980 0.760 9.140 1.240 ;
        RECT  8.860 1.900 9.020 2.840 ;
        RECT  8.140 1.080 8.980 1.240 ;
        RECT  8.260 1.900 8.860 2.060 ;
        RECT  7.820 0.760 8.740 0.920 ;
        RECT  8.460 2.220 8.700 2.960 ;
        RECT  7.820 2.800 8.460 2.960 ;
        RECT  8.140 1.900 8.260 2.640 ;
        RECT  7.980 1.080 8.140 2.640 ;
        RECT  7.660 0.760 7.820 2.960 ;
        RECT  7.560 1.020 7.660 1.300 ;
        RECT  7.500 1.930 7.660 2.580 ;
        RECT  6.710 1.140 7.560 1.300 ;
        RECT  6.710 1.930 7.500 2.090 ;
        RECT  7.340 2.760 7.500 3.040 ;
        RECT  7.290 0.440 7.450 0.720 ;
        RECT  3.350 2.880 7.340 3.040 ;
        RECT  5.710 0.560 7.290 0.720 ;
        RECT  6.350 1.460 6.970 1.620 ;
        RECT  6.550 1.020 6.710 1.300 ;
        RECT  6.550 1.930 6.710 2.610 ;
        RECT  6.030 1.930 6.550 2.090 ;
        RECT  6.190 0.880 6.350 1.620 ;
        RECT  4.990 0.880 6.190 1.040 ;
        RECT  5.870 1.600 6.030 2.090 ;
        RECT  5.550 0.440 5.710 0.720 ;
        RECT  3.930 0.560 5.550 0.720 ;
        RECT  4.990 2.260 5.410 2.420 ;
        RECT  4.830 0.880 4.990 2.420 ;
        RECT  4.090 0.880 4.830 1.040 ;
        RECT  3.670 2.260 4.830 2.420 ;
        RECT  4.110 1.810 4.670 2.090 ;
        RECT  3.930 1.810 4.110 1.970 ;
        RECT  3.770 0.560 3.930 1.970 ;
        RECT  2.890 1.210 3.770 1.370 ;
        RECT  3.510 2.140 3.670 2.420 ;
        RECT  3.350 1.530 3.610 1.690 ;
        RECT  3.190 1.530 3.350 3.040 ;
        RECT  2.570 0.440 3.290 0.600 ;
        RECT  1.550 2.880 3.190 3.040 ;
        RECT  2.730 1.030 2.890 2.720 ;
        RECT  2.650 2.440 2.730 2.720 ;
        RECT  1.450 2.560 2.650 2.720 ;
        RECT  2.410 0.440 2.570 1.190 ;
        RECT  1.770 1.030 2.410 1.190 ;
        RECT  1.770 2.120 1.890 2.400 ;
        RECT  1.610 1.030 1.770 2.400 ;
        RECT  1.440 0.440 1.670 0.720 ;
        RECT  1.510 1.030 1.610 1.320 ;
        RECT  1.390 2.880 1.550 3.160 ;
        RECT  1.290 1.580 1.450 2.720 ;
        RECT  0.310 0.560 1.440 0.720 ;
        RECT  1.130 2.880 1.390 3.040 ;
        RECT  1.130 1.090 1.310 1.250 ;
        RECT  0.970 1.090 1.130 3.040 ;
        RECT  0.140 0.560 0.310 2.190 ;
    END
END DFFHQX4TR

MACRO DFFHQX2TR
    CLASS CORE ;
    FOREIGN DFFHQX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.710 0.440 8.720 2.070 ;
        RECT  8.430 0.440 8.710 3.140 ;
        END
        ANTENNADIFFAREA 3.488 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 0.840 0.760 1.480 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.840 1.960 1.320 ;
        END
        ANTENNAGATEAREA 0.216 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.230 -0.280 8.800 0.280 ;
        RECT  7.420 -0.280 8.230 0.780 ;
        RECT  3.380 -0.280 7.420 0.340 ;
        RECT  3.100 -0.280 3.380 0.670 ;
        RECT  0.910 -0.280 3.100 0.340 ;
        RECT  0.620 -0.280 0.910 0.430 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.190 3.320 8.800 3.880 ;
        RECT  7.910 2.500 8.190 3.880 ;
        RECT  5.400 3.260 7.910 3.880 ;
        RECT  4.320 3.200 5.400 3.880 ;
        RECT  2.880 3.320 4.320 3.880 ;
        RECT  2.600 3.200 2.880 3.880 ;
        RECT  1.000 3.320 2.600 3.880 ;
        RECT  0.660 3.200 1.000 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.110 1.110 8.270 2.070 ;
        RECT  7.790 1.110 8.110 1.270 ;
        RECT  7.790 1.910 8.110 2.070 ;
        RECT  7.670 1.430 7.950 1.710 ;
        RECT  7.510 0.990 7.790 1.270 ;
        RECT  7.670 1.910 7.790 2.190 ;
        RECT  7.350 1.430 7.670 1.590 ;
        RECT  7.510 1.910 7.670 3.040 ;
        RECT  7.180 2.870 7.510 3.040 ;
        RECT  7.190 1.110 7.350 2.630 ;
        RECT  6.780 1.110 7.190 1.270 ;
        RECT  6.820 2.470 7.190 2.630 ;
        RECT  6.750 1.440 7.030 2.310 ;
        RECT  6.540 2.470 6.820 2.750 ;
        RECT  6.500 0.500 6.780 1.270 ;
        RECT  6.340 1.440 6.750 1.600 ;
        RECT  5.860 2.470 6.540 2.630 ;
        RECT  6.180 0.500 6.340 1.600 ;
        RECT  6.060 1.990 6.340 2.270 ;
        RECT  3.700 0.500 6.180 0.660 ;
        RECT  6.030 1.320 6.180 1.600 ;
        RECT  5.860 2.820 6.140 3.100 ;
        RECT  5.870 1.990 6.060 2.150 ;
        RECT  5.870 0.880 6.020 1.160 ;
        RECT  5.710 0.880 5.870 2.150 ;
        RECT  5.580 2.350 5.860 2.630 ;
        RECT  4.250 2.820 5.860 2.980 ;
        RECT  5.000 1.990 5.710 2.150 ;
        RECT  5.020 1.120 5.300 1.620 ;
        RECT  4.220 1.120 5.020 1.280 ;
        RECT  4.860 1.990 5.000 2.550 ;
        RECT  4.700 1.440 4.860 2.550 ;
        RECT  4.580 1.440 4.700 1.740 ;
        RECT  4.090 2.500 4.250 2.980 ;
        RECT  4.100 0.880 4.220 1.280 ;
        RECT  3.940 0.880 4.100 1.720 ;
        RECT  3.280 2.500 4.090 2.720 ;
        RECT  3.720 1.560 3.940 1.720 ;
        RECT  3.650 2.880 3.930 3.160 ;
        RECT  3.440 1.560 3.720 2.170 ;
        RECT  3.540 0.500 3.700 0.990 ;
        RECT  0.420 2.880 3.650 3.040 ;
        RECT  3.280 1.180 3.580 1.400 ;
        RECT  2.860 0.830 3.540 0.990 ;
        RECT  3.120 1.180 3.280 2.720 ;
        RECT  1.080 2.550 3.120 2.720 ;
        RECT  2.860 1.560 2.960 1.840 ;
        RECT  2.840 0.790 2.860 1.840 ;
        RECT  2.680 0.790 2.840 2.110 ;
        RECT  2.580 0.790 2.680 1.070 ;
        RECT  1.960 1.950 2.680 2.110 ;
        RECT  2.400 1.360 2.520 1.640 ;
        RECT  2.240 0.690 2.400 1.640 ;
        RECT  2.120 0.690 2.240 0.970 ;
        RECT  1.520 1.480 2.240 1.640 ;
        RECT  1.680 1.950 1.960 2.280 ;
        RECT  1.240 1.480 1.520 2.030 ;
        RECT  1.080 0.680 1.380 0.960 ;
        RECT  0.920 0.680 1.080 2.720 ;
        RECT  0.310 1.910 0.420 3.040 ;
        RECT  0.260 0.870 0.310 3.040 ;
        RECT  0.090 0.870 0.260 2.190 ;
    END
END DFFHQX2TR

MACRO DFFHQX1TR
    CLASS CORE ;
    FOREIGN DFFHQX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.660 0.840 7.920 3.020 ;
        END
        ANTENNADIFFAREA 1.957 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.220 0.760 1.660 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.620 0.840 1.960 1.410 ;
        END
        ANTENNAGATEAREA 0.1752 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 -0.280 8.000 0.280 ;
        RECT  7.020 -0.280 7.320 0.690 ;
        RECT  3.290 -0.280 7.020 0.290 ;
        RECT  2.960 -0.280 3.290 0.370 ;
        RECT  1.930 -0.280 2.960 0.290 ;
        RECT  1.700 -0.280 1.930 0.390 ;
        RECT  0.880 -0.280 1.700 0.290 ;
        RECT  0.600 -0.280 0.880 0.740 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.360 3.320 8.000 3.880 ;
        RECT  7.080 2.860 7.360 3.880 ;
        RECT  6.570 3.320 7.080 3.880 ;
        RECT  6.330 2.800 6.570 3.880 ;
        RECT  4.510 3.320 6.330 3.880 ;
        RECT  4.290 2.700 4.510 3.880 ;
        RECT  2.970 3.320 4.290 3.880 ;
        RECT  2.690 3.200 2.970 3.880 ;
        RECT  0.440 3.320 2.690 3.880 ;
        RECT  0.160 2.720 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.210 1.100 7.380 2.060 ;
        RECT  6.890 1.100 7.210 1.260 ;
        RECT  6.940 1.900 7.210 2.060 ;
        RECT  6.890 1.420 7.050 1.700 ;
        RECT  6.780 1.900 6.940 2.560 ;
        RECT  6.610 0.980 6.890 1.260 ;
        RECT  6.200 1.420 6.890 1.580 ;
        RECT  6.430 1.900 6.780 2.180 ;
        RECT  6.190 1.420 6.200 2.560 ;
        RECT  6.000 0.910 6.190 2.560 ;
        RECT  4.830 3.000 6.030 3.160 ;
        RECT  5.790 0.910 6.000 1.230 ;
        RECT  5.630 2.400 6.000 2.560 ;
        RECT  5.630 1.960 5.840 2.180 ;
        RECT  5.470 0.450 5.630 2.180 ;
        RECT  5.470 2.400 5.630 2.620 ;
        RECT  5.290 0.450 5.470 0.690 ;
        RECT  5.150 0.850 5.310 2.140 ;
        RECT  3.020 0.530 5.290 0.690 ;
        RECT  4.990 1.980 5.150 2.790 ;
        RECT  4.830 1.110 4.990 1.630 ;
        RECT  4.400 1.980 4.990 2.140 ;
        RECT  4.010 1.110 4.830 1.270 ;
        RECT  4.670 2.340 4.830 3.160 ;
        RECT  3.990 2.340 4.670 2.500 ;
        RECT  4.240 1.460 4.400 2.140 ;
        RECT  3.860 0.850 4.010 1.270 ;
        RECT  3.830 2.340 3.990 2.930 ;
        RECT  3.700 0.850 3.860 2.130 ;
        RECT  3.360 2.340 3.830 2.500 ;
        RECT  3.530 1.880 3.700 2.130 ;
        RECT  2.600 2.730 3.610 2.890 ;
        RECT  3.190 1.120 3.360 2.500 ;
        RECT  2.280 2.340 3.190 2.500 ;
        RECT  2.860 0.530 3.020 2.130 ;
        RECT  2.440 0.530 2.860 0.740 ;
        RECT  1.900 1.970 2.860 2.130 ;
        RECT  2.340 1.450 2.610 1.730 ;
        RECT  2.440 2.730 2.600 3.050 ;
        RECT  0.760 2.890 2.440 3.050 ;
        RECT  2.180 0.960 2.340 1.730 ;
        RECT  2.120 2.340 2.280 2.720 ;
        RECT  1.520 1.570 2.180 1.730 ;
        RECT  1.080 2.560 2.120 2.720 ;
        RECT  1.740 1.970 1.900 2.340 ;
        RECT  1.240 1.570 1.520 2.190 ;
        RECT  1.080 0.780 1.360 1.060 ;
        RECT  0.920 0.900 1.080 2.720 ;
        RECT  0.600 1.980 0.760 3.050 ;
        RECT  0.320 1.980 0.600 2.140 ;
        RECT  0.100 0.980 0.320 2.190 ;
    END
END DFFHQX1TR

MACRO DFFXLTR
    CLASS CORE ;
    FOREIGN DFFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.840 1.030 7.120 2.360 ;
        END
        ANTENNADIFFAREA 1.158 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.520 0.560 6.680 2.200 ;
        RECT  5.940 0.560 6.520 0.720 ;
        RECT  6.360 2.040 6.520 2.200 ;
        RECT  6.240 2.040 6.360 2.360 ;
        RECT  6.080 2.040 6.240 3.070 ;
        RECT  5.700 2.790 6.080 3.070 ;
        RECT  5.660 0.440 5.940 0.720 ;
        END
        ANTENNADIFFAREA 0.996 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 2.440 0.720 2.760 ;
        RECT  0.270 1.960 0.430 2.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.590 3.120 1.960 ;
        RECT  2.770 1.680 2.840 1.960 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.500 -0.280 7.200 0.280 ;
        RECT  6.220 -0.280 6.500 0.400 ;
        RECT  5.480 -0.280 6.220 0.280 ;
        RECT  5.200 -0.280 5.480 0.400 ;
        RECT  3.480 -0.280 5.200 0.340 ;
        RECT  2.210 -0.280 3.480 0.280 ;
        RECT  1.930 -0.280 2.210 0.670 ;
        RECT  0.400 -0.280 1.930 0.340 ;
        RECT  0.120 -0.280 0.400 0.400 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.680 3.320 7.200 3.880 ;
        RECT  6.400 2.640 6.680 3.880 ;
        RECT  5.360 3.320 6.400 3.880 ;
        RECT  5.080 2.710 5.360 3.880 ;
        RECT  3.360 3.260 5.080 3.880 ;
        RECT  2.490 3.320 3.360 3.880 ;
        RECT  1.810 3.260 2.490 3.880 ;
        RECT  0.400 3.320 1.810 3.880 ;
        RECT  0.120 3.200 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 1.580 6.360 1.880 ;
        RECT  6.080 0.900 6.240 1.880 ;
        RECT  5.660 0.900 6.080 1.120 ;
        RECT  5.800 1.720 6.080 1.880 ;
        RECT  5.640 1.280 5.920 1.560 ;
        RECT  5.800 2.270 5.920 2.550 ;
        RECT  5.640 1.720 5.800 2.550 ;
        RECT  5.040 1.280 5.640 1.440 ;
        RECT  5.480 1.720 5.640 1.880 ;
        RECT  5.200 1.600 5.480 1.880 ;
        RECT  4.880 0.590 5.040 2.390 ;
        RECT  4.240 0.590 4.880 0.870 ;
        RECT  4.580 2.230 4.880 2.390 ;
        RECT  4.440 1.030 4.720 1.950 ;
        RECT  4.360 2.230 4.580 2.510 ;
        RECT  3.760 1.030 4.440 1.190 ;
        RECT  4.320 1.790 4.440 1.950 ;
        RECT  4.200 1.790 4.320 2.070 ;
        RECT  4.000 1.350 4.280 1.630 ;
        RECT  4.040 1.790 4.200 3.100 ;
        RECT  1.530 2.880 4.040 3.100 ;
        RECT  3.440 1.350 4.000 1.510 ;
        RECT  3.600 1.790 3.880 2.720 ;
        RECT  3.600 0.500 3.760 1.190 ;
        RECT  2.840 0.500 3.600 0.780 ;
        RECT  2.530 2.560 3.600 2.720 ;
        RECT  3.280 1.060 3.440 2.400 ;
        RECT  3.190 1.060 3.280 1.220 ;
        RECT  2.910 2.120 3.280 2.400 ;
        RECT  2.910 0.940 3.190 1.220 ;
        RECT  1.770 0.940 2.910 1.100 ;
        RECT  2.680 0.450 2.840 0.780 ;
        RECT  2.560 0.450 2.680 0.670 ;
        RECT  2.530 1.260 2.610 2.240 ;
        RECT  2.450 1.260 2.530 2.720 ;
        RECT  2.330 1.260 2.450 1.480 ;
        RECT  2.250 2.080 2.450 2.720 ;
        RECT  2.170 1.640 2.290 1.920 ;
        RECT  1.850 2.080 2.250 2.240 ;
        RECT  2.010 1.260 2.170 1.920 ;
        RECT  1.450 1.260 2.010 1.420 ;
        RECT  1.570 1.960 1.850 2.240 ;
        RECT  1.610 0.500 1.770 1.100 ;
        RECT  1.120 0.500 1.610 0.720 ;
        RECT  1.390 2.400 1.530 3.100 ;
        RECT  1.290 0.880 1.450 1.420 ;
        RECT  1.370 1.580 1.390 3.100 ;
        RECT  1.230 1.580 1.370 2.560 ;
        RECT  0.450 0.880 1.290 1.100 ;
        RECT  1.130 1.580 1.230 1.740 ;
        RECT  1.050 2.880 1.210 3.160 ;
        RECT  0.970 1.260 1.130 1.740 ;
        RECT  0.890 1.900 1.050 3.160 ;
        RECT  0.640 1.260 0.970 1.480 ;
        RECT  0.810 1.900 0.890 2.060 ;
        RECT  0.650 1.640 0.810 2.060 ;
        RECT  0.450 1.640 0.650 1.800 ;
        RECT  0.290 0.880 0.450 1.800 ;
    END
END DFFXLTR

MACRO DFFX4TR
    CLASS CORE ;
    FOREIGN DFFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.230 1.440 10.320 2.160 ;
        RECT  10.030 0.500 10.230 3.160 ;
        RECT  9.950 0.500 10.030 1.320 ;
        RECT  9.950 2.020 10.030 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.990 0.500 9.270 2.300 ;
        RECT  8.880 1.440 8.990 2.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.640 0.530 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.820 2.760 2.360 ;
        END
        ANTENNAGATEAREA 0.228 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 -0.280 10.800 0.280 ;
        RECT  10.430 -0.280 10.710 1.180 ;
        RECT  9.750 -0.280 10.430 0.280 ;
        RECT  9.470 -0.280 9.750 1.310 ;
        RECT  8.790 -0.280 9.470 0.280 ;
        RECT  8.510 -0.280 8.790 1.080 ;
        RECT  7.850 -0.280 8.510 0.280 ;
        RECT  7.630 -0.280 7.850 1.310 ;
        RECT  6.120 -0.280 7.630 0.340 ;
        RECT  5.840 -0.280 6.120 0.610 ;
        RECT  4.400 -0.280 5.840 0.280 ;
        RECT  4.120 -0.280 4.400 0.990 ;
        RECT  2.910 -0.280 4.120 0.280 ;
        RECT  2.630 -0.280 2.910 0.890 ;
        RECT  2.090 -0.280 2.630 0.280 ;
        RECT  1.810 -0.280 2.090 0.990 ;
        RECT  0.370 -0.280 1.810 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.710 3.320 10.800 3.880 ;
        RECT  10.430 2.480 10.710 3.880 ;
        RECT  9.750 3.320 10.430 3.880 ;
        RECT  9.470 2.930 9.750 3.880 ;
        RECT  8.790 3.320 9.470 3.880 ;
        RECT  8.510 2.930 8.790 3.880 ;
        RECT  7.850 3.320 8.510 3.880 ;
        RECT  7.570 2.340 7.850 3.880 ;
        RECT  6.080 3.320 7.570 3.880 ;
        RECT  5.800 2.900 6.080 3.880 ;
        RECT  4.360 3.320 5.800 3.880 ;
        RECT  4.080 3.240 4.360 3.880 ;
        RECT  2.750 3.260 4.080 3.880 ;
        RECT  2.050 3.320 2.750 3.880 ;
        RECT  1.770 3.260 2.050 3.880 ;
        RECT  0.410 3.320 1.770 3.880 ;
        RECT  0.130 2.740 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.750 1.580 9.870 1.860 ;
        RECT  9.590 1.580 9.750 2.620 ;
        RECT  8.330 2.460 9.590 2.620 ;
        RECT  8.420 1.260 8.580 2.180 ;
        RECT  8.330 1.260 8.420 1.420 ;
        RECT  8.330 2.020 8.420 2.180 ;
        RECT  8.050 0.600 8.330 1.420 ;
        RECT  8.050 2.020 8.330 3.160 ;
        RECT  7.460 1.580 8.260 1.860 ;
        RECT  7.410 2.020 8.050 2.180 ;
        RECT  7.300 0.770 7.460 1.860 ;
        RECT  7.250 2.020 7.410 3.160 ;
        RECT  5.000 0.770 7.300 0.990 ;
        RECT  7.000 1.700 7.300 1.860 ;
        RECT  7.130 2.880 7.250 3.160 ;
        RECT  6.920 1.150 7.140 1.430 ;
        RECT  6.880 1.700 7.000 2.600 ;
        RECT  6.560 1.150 6.920 1.310 ;
        RECT  6.840 1.700 6.880 3.160 ;
        RECT  6.600 2.440 6.840 3.160 ;
        RECT  6.560 1.870 6.680 2.280 ;
        RECT  5.280 2.440 6.600 2.600 ;
        RECT  6.400 1.150 6.560 2.280 ;
        RECT  4.240 1.150 6.400 1.310 ;
        RECT  5.120 2.120 6.400 2.280 ;
        RECT  5.600 1.530 6.240 1.810 ;
        RECT  4.680 1.530 5.600 1.690 ;
        RECT  5.000 2.440 5.280 3.160 ;
        RECT  4.840 1.850 5.120 2.280 ;
        RECT  4.600 2.120 4.840 2.280 ;
        RECT  4.400 1.530 4.680 1.960 ;
        RECT  4.440 2.120 4.600 3.080 ;
        RECT  1.540 2.920 4.440 3.080 ;
        RECT  4.280 1.800 4.400 1.960 ;
        RECT  4.120 1.800 4.280 2.760 ;
        RECT  4.080 1.150 4.240 1.640 ;
        RECT  3.430 2.600 4.120 2.760 ;
        RECT  3.910 1.360 4.080 1.640 ;
        RECT  3.750 2.030 3.960 2.310 ;
        RECT  3.750 0.920 3.920 1.200 ;
        RECT  3.590 0.440 3.750 2.310 ;
        RECT  3.430 0.440 3.590 0.720 ;
        RECT  3.270 0.910 3.430 2.760 ;
        RECT  3.150 0.910 3.270 1.190 ;
        RECT  1.930 2.600 3.270 2.760 ;
        RECT  1.330 1.500 3.100 1.660 ;
        RECT  2.290 1.070 2.570 1.340 ;
        RECT  1.650 1.180 2.290 1.340 ;
        RECT  1.770 1.870 1.930 2.760 ;
        RECT  1.650 1.870 1.770 2.150 ;
        RECT  1.490 0.560 1.650 1.340 ;
        RECT  1.530 2.860 1.540 3.080 ;
        RECT  1.250 2.860 1.530 3.140 ;
        RECT  0.770 0.560 1.490 0.720 ;
        RECT  1.170 0.880 1.330 2.700 ;
        RECT  0.850 2.860 1.250 3.020 ;
        RECT  0.930 0.880 1.170 1.160 ;
        RECT  1.010 2.020 1.170 2.700 ;
        RECT  0.850 1.320 1.010 1.630 ;
        RECT  0.770 1.320 0.850 3.020 ;
        RECT  0.690 0.560 0.770 3.020 ;
        RECT  0.610 0.560 0.690 1.480 ;
    END
END DFFX4TR

MACRO DFFX2TR
    CLASS CORE ;
    FOREIGN DFFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.430 1.240 9.520 2.360 ;
        RECT  9.230 0.500 9.430 3.160 ;
        RECT  9.150 0.500 9.230 1.320 ;
        RECT  9.150 2.020 9.230 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.190 0.500 8.470 2.300 ;
        RECT  8.080 1.640 8.190 1.960 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.740 0.400 2.030 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0792 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.820 2.380 2.360 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.950 -0.280 9.600 0.280 ;
        RECT  8.670 -0.280 8.950 1.310 ;
        RECT  7.450 -0.280 8.670 0.280 ;
        RECT  7.230 -0.280 7.450 1.110 ;
        RECT  5.720 -0.280 7.230 0.340 ;
        RECT  5.440 -0.280 5.720 0.610 ;
        RECT  4.200 -0.280 5.440 0.280 ;
        RECT  3.920 -0.280 4.200 0.990 ;
        RECT  2.740 -0.280 3.920 0.280 ;
        RECT  2.460 -0.280 2.740 0.840 ;
        RECT  1.880 -0.280 2.460 0.280 ;
        RECT  1.600 -0.280 1.880 0.810 ;
        RECT  0.400 -0.280 1.600 0.280 ;
        RECT  0.120 -0.280 0.400 0.680 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.950 3.320 9.600 3.880 ;
        RECT  8.670 2.930 8.950 3.880 ;
        RECT  7.450 3.320 8.670 3.880 ;
        RECT  7.170 2.340 7.450 3.880 ;
        RECT  5.680 3.320 7.170 3.880 ;
        RECT  5.400 2.680 5.680 3.880 ;
        RECT  4.320 3.320 5.400 3.880 ;
        RECT  4.040 3.240 4.320 3.880 ;
        RECT  2.580 3.260 4.040 3.880 ;
        RECT  1.880 3.320 2.580 3.880 ;
        RECT  1.600 3.260 1.880 3.880 ;
        RECT  0.400 3.320 1.600 3.880 ;
        RECT  0.120 3.150 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.950 1.580 9.070 1.860 ;
        RECT  8.790 1.580 8.950 2.620 ;
        RECT  7.930 2.460 8.790 2.620 ;
        RECT  7.920 2.460 7.930 2.780 ;
        RECT  7.760 0.900 7.920 2.780 ;
        RECT  7.650 0.900 7.760 1.420 ;
        RECT  7.650 2.020 7.760 2.780 ;
        RECT  7.010 2.020 7.650 2.180 ;
        RECT  7.060 1.580 7.600 1.860 ;
        RECT  6.900 0.770 7.060 1.860 ;
        RECT  6.850 2.020 7.010 3.160 ;
        RECT  4.600 0.770 6.900 0.990 ;
        RECT  6.600 1.700 6.900 1.860 ;
        RECT  6.730 2.880 6.850 3.160 ;
        RECT  6.520 1.150 6.740 1.430 ;
        RECT  6.440 1.700 6.600 2.600 ;
        RECT  6.160 1.150 6.520 1.310 ;
        RECT  6.200 2.360 6.440 2.600 ;
        RECT  6.160 1.870 6.280 2.200 ;
        RECT  4.880 2.360 6.200 2.520 ;
        RECT  6.000 1.150 6.160 2.200 ;
        RECT  4.060 1.150 6.000 1.310 ;
        RECT  5.080 2.040 6.000 2.200 ;
        RECT  5.340 1.530 5.720 1.810 ;
        RECT  4.420 1.530 5.340 1.690 ;
        RECT  4.800 1.850 5.080 2.200 ;
        RECT  4.600 2.360 4.880 2.690 ;
        RECT  4.440 2.040 4.800 2.200 ;
        RECT  4.280 2.040 4.440 3.080 ;
        RECT  4.220 1.530 4.420 1.880 ;
        RECT  1.370 2.920 4.280 3.080 ;
        RECT  4.120 1.720 4.220 1.880 ;
        RECT  3.960 1.720 4.120 2.760 ;
        RECT  3.900 1.150 4.060 1.560 ;
        RECT  3.200 2.600 3.960 2.760 ;
        RECT  3.710 1.340 3.900 1.560 ;
        RECT  3.550 2.030 3.790 2.310 ;
        RECT  3.550 0.820 3.720 1.100 ;
        RECT  3.390 0.440 3.550 2.310 ;
        RECT  3.230 0.440 3.390 0.720 ;
        RECT  3.040 0.910 3.200 2.760 ;
        RECT  2.980 0.910 3.040 1.190 ;
        RECT  1.890 2.600 3.040 2.760 ;
        RECT  2.710 1.440 2.870 1.720 ;
        RECT  1.060 1.500 2.710 1.660 ;
        RECT  2.120 1.020 2.400 1.340 ;
        RECT  1.380 1.180 2.120 1.340 ;
        RECT  1.730 1.870 1.890 2.760 ;
        RECT  1.610 1.870 1.730 2.150 ;
        RECT  1.220 0.700 1.380 1.340 ;
        RECT  1.360 2.860 1.370 3.080 ;
        RECT  1.080 2.860 1.360 3.140 ;
        RECT  0.720 0.700 1.220 0.860 ;
        RECT  0.720 2.860 1.080 3.020 ;
        RECT  0.900 1.020 1.060 2.700 ;
        RECT  0.880 2.020 0.900 2.700 ;
        RECT  0.560 0.700 0.720 3.020 ;
    END
END DFFX2TR

MACRO DFFX1TR
    CLASS CORE ;
    FOREIGN DFFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 0.620 7.520 3.010 ;
        RECT  6.960 2.730 7.280 3.010 ;
        END
        ANTENNADIFFAREA 2.496 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 0.690 7.120 2.330 ;
        RECT  6.080 0.690 6.960 0.850 ;
        RECT  6.320 2.170 6.960 2.330 ;
        RECT  6.240 2.170 6.320 2.760 ;
        RECT  6.160 2.170 6.240 3.030 ;
        RECT  6.080 2.440 6.160 3.030 ;
        RECT  5.920 0.570 6.080 0.850 ;
        RECT  5.940 2.870 6.080 3.030 ;
        END
        ANTENNADIFFAREA 1.544 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.980 0.560 2.140 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.590 3.120 1.960 ;
        RECT  2.770 1.800 2.880 1.960 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.660 -0.280 7.600 0.280 ;
        RECT  6.380 -0.280 6.660 0.340 ;
        RECT  5.540 -0.280 6.380 0.280 ;
        RECT  5.260 -0.280 5.540 0.800 ;
        RECT  3.790 -0.280 5.260 0.280 ;
        RECT  3.510 -0.280 3.790 0.340 ;
        RECT  2.160 -0.280 3.510 0.280 ;
        RECT  2.000 -0.280 2.160 0.670 ;
        RECT  0.410 -0.280 2.000 0.280 ;
        RECT  0.130 -0.280 0.410 0.350 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.640 3.320 7.600 3.880 ;
        RECT  6.480 2.490 6.640 3.880 ;
        RECT  5.360 3.320 6.480 3.880 ;
        RECT  5.080 2.860 5.360 3.880 ;
        RECT  3.660 3.320 5.080 3.880 ;
        RECT  3.380 3.260 3.660 3.880 ;
        RECT  2.550 3.320 3.380 3.880 ;
        RECT  1.870 3.260 2.550 3.880 ;
        RECT  0.410 3.320 1.870 3.880 ;
        RECT  0.130 3.260 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.570 1.090 6.800 2.010 ;
        RECT  5.820 1.090 6.570 1.250 ;
        RECT  5.820 1.850 6.570 2.010 ;
        RECT  5.670 1.410 6.240 1.690 ;
        RECT  5.660 1.850 5.820 2.630 ;
        RECT  4.980 1.410 5.670 1.570 ;
        RECT  5.420 1.850 5.660 2.010 ;
        RECT  5.140 1.740 5.420 2.010 ;
        RECT  4.820 0.840 4.980 2.420 ;
        RECT  4.270 0.840 4.820 1.000 ;
        RECT  4.440 2.260 4.820 2.420 ;
        RECT  4.500 1.160 4.660 2.100 ;
        RECT  3.760 1.160 4.500 1.320 ;
        RECT  4.120 1.940 4.500 2.100 ;
        RECT  4.280 2.260 4.440 3.010 ;
        RECT  3.440 1.540 4.310 1.700 ;
        RECT  3.960 1.940 4.120 3.070 ;
        RECT  1.530 2.910 3.960 3.070 ;
        RECT  3.640 1.880 3.800 2.750 ;
        RECT  3.600 0.640 3.760 1.320 ;
        RECT  2.490 2.590 3.640 2.750 ;
        RECT  2.870 0.640 3.600 0.800 ;
        RECT  3.280 1.150 3.440 2.430 ;
        RECT  3.160 1.150 3.280 1.310 ;
        RECT  2.940 2.270 3.280 2.430 ;
        RECT  3.000 0.960 3.160 1.310 ;
        RECT  1.840 0.960 3.000 1.120 ;
        RECT  2.710 0.510 2.870 0.800 ;
        RECT  2.590 0.510 2.710 0.670 ;
        RECT  2.490 1.280 2.610 2.260 ;
        RECT  2.450 1.280 2.490 2.750 ;
        RECT  2.330 1.280 2.450 1.440 ;
        RECT  2.330 2.100 2.450 2.750 ;
        RECT  1.850 2.100 2.330 2.260 ;
        RECT  2.130 1.600 2.290 1.940 ;
        RECT  1.520 1.600 2.130 1.760 ;
        RECT  1.690 1.920 1.850 2.260 ;
        RECT  1.680 0.450 1.840 1.120 ;
        RECT  1.220 0.450 1.680 0.610 ;
        RECT  1.370 1.980 1.530 3.070 ;
        RECT  1.360 0.850 1.520 1.760 ;
        RECT  1.200 1.980 1.370 2.140 ;
        RECT  0.650 0.850 1.360 1.010 ;
        RECT  1.050 2.300 1.210 2.580 ;
        RECT  1.040 1.200 1.200 2.140 ;
        RECT  0.880 2.300 1.050 2.460 ;
        RECT  0.820 1.200 1.040 1.480 ;
        RECT  0.720 1.660 0.880 2.460 ;
        RECT  0.650 1.660 0.720 1.820 ;
        RECT  0.490 0.850 0.650 1.820 ;
    END
END DFFX1TR

MACRO CLKXOR2X8TR
    CLASS CORE ;
    FOREIGN CLKXOR2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.110 0.980 8.390 3.160 ;
        RECT  7.430 1.230 8.110 2.170 ;
        RECT  7.170 0.980 7.430 3.160 ;
        RECT  7.150 0.980 7.170 1.390 ;
        RECT  7.150 1.990 7.170 3.160 ;
        END
        ANTENNADIFFAREA 6.3 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.580 1.050 1.860 ;
        RECT  0.440 1.580 0.760 1.960 ;
        RECT  0.370 1.580 0.440 1.860 ;
        END
        ANTENNAGATEAREA 0.6552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.690 2.670 1.970 ;
        RECT  1.640 1.240 1.960 1.970 ;
        END
        ANTENNAGATEAREA 0.7032 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.870 -0.280 9.200 0.280 ;
        RECT  8.590 -0.280 8.870 1.070 ;
        RECT  7.910 -0.280 8.590 0.280 ;
        RECT  7.630 -0.280 7.910 1.070 ;
        RECT  6.910 -0.280 7.630 0.280 ;
        RECT  6.630 -0.280 6.910 0.400 ;
        RECT  5.870 -0.280 6.630 0.280 ;
        RECT  5.590 -0.280 5.870 0.400 ;
        RECT  1.850 -0.280 5.590 0.280 ;
        RECT  1.570 -0.280 1.850 0.320 ;
        RECT  0.850 -0.280 1.570 0.280 ;
        RECT  0.570 -0.280 0.850 1.000 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.870 3.320 9.200 3.880 ;
        RECT  8.590 1.910 8.870 3.880 ;
        RECT  7.910 3.320 8.590 3.880 ;
        RECT  7.630 2.400 7.910 3.880 ;
        RECT  6.950 3.320 7.630 3.880 ;
        RECT  6.670 2.670 6.950 3.880 ;
        RECT  5.990 3.260 6.670 3.880 ;
        RECT  5.710 2.670 5.990 3.880 ;
        RECT  1.810 3.320 5.710 3.880 ;
        RECT  1.530 2.930 1.810 3.880 ;
        RECT  0.850 3.320 1.530 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.790 1.550 7.010 1.830 ;
        RECT  6.630 0.590 6.790 2.510 ;
        RECT  4.750 0.590 6.630 0.750 ;
        RECT  5.550 2.350 6.630 2.510 ;
        RECT  6.390 1.030 6.470 2.190 ;
        RECT  6.310 0.910 6.390 2.190 ;
        RECT  6.110 0.910 6.310 1.190 ;
        RECT  6.190 1.910 6.310 2.190 ;
        RECT  5.510 1.910 6.190 2.070 ;
        RECT  5.510 1.470 6.150 1.750 ;
        RECT  4.270 1.030 6.110 1.190 ;
        RECT  5.390 2.350 5.550 2.990 ;
        RECT  4.670 1.590 5.510 1.750 ;
        RECT  5.230 1.910 5.510 2.190 ;
        RECT  5.030 2.830 5.390 2.990 ;
        RECT  5.070 1.910 5.230 2.500 ;
        RECT  4.550 2.340 5.070 2.500 ;
        RECT  4.750 2.710 5.030 2.990 ;
        RECT  4.470 0.590 4.750 0.870 ;
        RECT  4.070 2.830 4.750 2.990 ;
        RECT  4.510 1.590 4.670 2.180 ;
        RECT  4.270 2.340 4.550 2.620 ;
        RECT  3.590 2.020 4.510 2.180 ;
        RECT  3.790 0.590 4.470 0.750 ;
        RECT  3.510 1.580 4.350 1.860 ;
        RECT  3.990 0.910 4.270 1.190 ;
        RECT  3.790 2.340 4.070 2.990 ;
        RECT  3.670 0.590 3.790 0.870 ;
        RECT  3.110 2.820 3.790 2.990 ;
        RECT  3.510 0.590 3.670 1.190 ;
        RECT  3.310 2.020 3.590 2.660 ;
        RECT  2.830 1.030 3.510 1.190 ;
        RECT  3.350 1.350 3.510 1.860 ;
        RECT  2.990 1.350 3.350 1.630 ;
        RECT  3.030 0.480 3.310 0.870 ;
        RECT  2.630 2.500 3.310 2.660 ;
        RECT  2.830 2.820 3.110 3.100 ;
        RECT  1.370 0.480 3.030 0.640 ;
        RECT  2.830 1.350 2.990 2.330 ;
        RECT  2.550 0.910 2.830 1.190 ;
        RECT  2.370 1.350 2.830 1.510 ;
        RECT  2.290 2.170 2.830 2.330 ;
        RECT  2.470 2.500 2.630 3.100 ;
        RECT  2.350 2.610 2.470 3.100 ;
        RECT  2.210 0.800 2.370 1.510 ;
        RECT  1.370 2.610 2.350 2.770 ;
        RECT  2.010 2.170 2.290 2.450 ;
        RECT  2.090 0.800 2.210 1.080 ;
        RECT  1.330 0.480 1.370 2.770 ;
        RECT  1.210 0.480 1.330 3.160 ;
        RECT  1.050 0.970 1.210 1.320 ;
        RECT  1.050 2.120 1.210 3.160 ;
        RECT  0.370 1.160 1.050 1.320 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 0.970 0.370 1.320 ;
        RECT  0.090 2.120 0.370 3.160 ;
    END
END CLKXOR2X8TR

MACRO CLKXOR2X4TR
    CLASS CORE ;
    FOREIGN CLKXOR2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.030 1.020 5.120 1.760 ;
        RECT  4.970 0.560 5.030 1.760 ;
        RECT  4.750 0.560 4.970 3.100 ;
        RECT  4.690 1.020 4.750 3.100 ;
        END
        ANTENNADIFFAREA 3.132 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.570 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.240 1.590 1.880 ;
        END
        ANTENNAGATEAREA 0.3552 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 -0.280 5.600 0.280 ;
        RECT  5.230 -0.280 5.510 0.720 ;
        RECT  4.550 -0.280 5.230 0.280 ;
        RECT  4.270 -0.280 4.550 0.720 ;
        RECT  1.330 -0.280 4.270 0.280 ;
        RECT  1.050 -0.280 1.330 1.080 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.470 3.320 5.600 3.880 ;
        RECT  5.190 1.940 5.470 3.880 ;
        RECT  4.490 3.320 5.190 3.880 ;
        RECT  4.270 1.940 4.490 3.880 ;
        RECT  1.370 3.260 4.270 3.880 ;
        RECT  1.090 2.800 1.370 3.880 ;
        RECT  0.370 3.320 1.090 3.880 ;
        RECT  0.090 2.590 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.310 0.880 4.490 1.370 ;
        RECT  4.110 0.880 4.310 1.040 ;
        RECT  3.950 0.440 4.110 1.040 ;
        RECT  3.950 1.260 4.110 3.100 ;
        RECT  3.350 0.440 3.950 0.600 ;
        RECT  3.830 1.260 3.950 1.540 ;
        RECT  2.870 2.940 3.950 3.100 ;
        RECT  3.670 0.760 3.790 1.040 ;
        RECT  3.670 1.700 3.790 2.780 ;
        RECT  3.510 0.760 3.670 2.780 ;
        RECT  3.190 0.440 3.350 2.780 ;
        RECT  3.030 0.440 3.190 1.020 ;
        RECT  3.070 2.020 3.190 2.780 ;
        RECT  2.390 0.440 3.030 0.600 ;
        RECT  2.710 2.020 2.870 3.100 ;
        RECT  2.710 0.760 2.830 1.040 ;
        RECT  2.550 0.760 2.710 3.100 ;
        RECT  1.690 2.940 2.550 3.100 ;
        RECT  2.230 0.440 2.390 2.780 ;
        RECT  2.070 0.740 2.230 1.020 ;
        RECT  2.110 2.020 2.230 2.780 ;
        RECT  1.910 1.350 2.070 1.630 ;
        RECT  1.750 0.800 1.910 2.320 ;
        RECT  1.610 0.800 1.750 1.080 ;
        RECT  1.610 2.040 1.750 2.320 ;
        RECT  1.530 2.480 1.690 3.100 ;
        RECT  0.890 2.480 1.530 2.640 ;
        RECT  0.850 0.800 0.890 2.640 ;
        RECT  0.730 0.800 0.850 3.100 ;
        RECT  0.570 0.800 0.730 1.080 ;
        RECT  0.570 2.020 0.730 3.100 ;
    END
END CLKXOR2X4TR

MACRO CLKXOR2X2TR
    CLASS CORE ;
    FOREIGN CLKXOR2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 0.840 3.520 2.540 ;
        RECT  3.280 0.840 3.410 3.100 ;
        RECT  3.140 0.840 3.280 1.120 ;
        RECT  3.140 2.280 3.280 3.100 ;
        END
        ANTENNADIFFAREA 2.848 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.240 1.120 2.030 ;
        RECT  0.880 1.030 1.040 2.030 ;
        RECT  0.820 1.030 0.880 1.360 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.530 0.720 1.970 ;
        END
        ANTENNAGATEAREA 0.2208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 -0.280 3.600 0.280 ;
        RECT  2.620 -0.280 2.900 0.600 ;
        RECT  0.720 -0.280 2.620 0.280 ;
        RECT  0.440 -0.280 0.720 0.400 ;
        RECT  0.000 -0.280 0.440 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 3.320 3.600 3.880 ;
        RECT  2.620 3.200 2.900 3.880 ;
        RECT  0.980 3.320 2.620 3.880 ;
        RECT  0.700 2.890 0.980 3.880 ;
        RECT  0.000 3.320 0.700 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.900 1.580 3.060 2.060 ;
        RECT  2.740 1.900 2.900 2.060 ;
        RECT  2.580 0.760 2.740 1.740 ;
        RECT  2.580 1.900 2.740 2.710 ;
        RECT  1.500 0.760 2.580 0.920 ;
        RECT  2.420 1.460 2.580 1.740 ;
        RECT  1.940 2.550 2.580 2.710 ;
        RECT  2.260 1.080 2.420 1.240 ;
        RECT  2.260 2.020 2.420 2.300 ;
        RECT  2.100 1.080 2.260 2.300 ;
        RECT  1.300 2.930 2.220 3.090 ;
        RECT  1.820 1.090 1.940 1.250 ;
        RECT  1.820 2.020 1.940 2.710 ;
        RECT  1.660 1.090 1.820 2.710 ;
        RECT  1.040 0.440 1.700 0.600 ;
        RECT  1.340 0.760 1.500 2.350 ;
        RECT  1.200 0.760 1.340 1.040 ;
        RECT  1.180 2.190 1.340 2.350 ;
        RECT  1.140 2.570 1.300 3.090 ;
        RECT  0.320 2.570 1.140 2.730 ;
        RECT  0.880 0.440 1.040 0.720 ;
        RECT  0.320 0.560 0.880 0.720 ;
        RECT  0.160 0.560 0.320 2.730 ;
        RECT  0.150 0.560 0.160 0.980 ;
    END
END CLKXOR2X2TR

MACRO CLKXOR2X1TR
    CLASS CORE ;
    FOREIGN CLKXOR2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.840 3.520 2.660 ;
        RECT  3.240 2.280 3.280 2.660 ;
        END
        ANTENNADIFFAREA 1.554 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.240 1.120 2.030 ;
        RECT  0.880 1.030 0.990 2.030 ;
        RECT  0.820 1.030 0.880 1.460 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.640 0.720 2.110 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.940 -0.280 3.600 0.280 ;
        RECT  2.660 -0.280 2.940 0.600 ;
        RECT  0.000 -0.280 2.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.940 3.320 3.600 3.880 ;
        RECT  2.660 2.870 2.940 3.880 ;
        RECT  0.940 3.320 2.660 3.880 ;
        RECT  0.650 2.890 0.940 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 1.690 3.080 2.710 ;
        RECT  1.940 2.550 2.920 2.710 ;
        RECT  2.600 0.760 2.760 1.740 ;
        RECT  1.500 0.760 2.600 0.920 ;
        RECT  2.420 1.520 2.600 1.740 ;
        RECT  2.260 1.080 2.440 1.310 ;
        RECT  2.260 2.130 2.420 2.390 ;
        RECT  2.100 1.080 2.260 2.390 ;
        RECT  1.300 2.930 2.220 3.090 ;
        RECT  1.820 1.090 1.940 1.310 ;
        RECT  1.820 2.270 1.940 2.710 ;
        RECT  1.660 1.090 1.820 2.710 ;
        RECT  0.990 0.440 1.700 0.600 ;
        RECT  1.340 0.760 1.500 2.350 ;
        RECT  1.150 0.760 1.340 1.040 ;
        RECT  1.180 2.190 1.340 2.350 ;
        RECT  1.140 2.570 1.300 3.090 ;
        RECT  0.320 2.570 1.140 2.730 ;
        RECT  0.830 0.440 0.990 0.720 ;
        RECT  0.320 0.560 0.830 0.720 ;
        RECT  0.160 0.560 0.320 2.730 ;
        RECT  0.150 0.560 0.160 0.980 ;
    END
END CLKXOR2X1TR

MACRO CLKMX2X8TR
    CLASS CORE ;
    FOREIGN CLKMX2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 1.040 6.230 3.160 ;
        RECT  5.510 1.040 5.950 2.400 ;
        RECT  5.270 0.450 5.510 2.400 ;
        RECT  5.230 0.450 5.270 3.160 ;
        RECT  4.990 1.910 5.230 3.160 ;
        END
        ANTENNADIFFAREA 6.632 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.730 1.560 3.160 ;
        END
        ANTENNAGATEAREA 0.1056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.120 1.620 ;
        END
        ANTENNAGATEAREA 0.1056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.030 -0.280 6.800 0.280 ;
        RECT  5.750 -0.280 6.030 0.800 ;
        RECT  4.950 -0.280 5.750 0.280 ;
        RECT  4.670 -0.280 4.950 1.310 ;
        RECT  3.480 -0.280 4.670 0.340 ;
        RECT  3.200 -0.280 3.480 1.080 ;
        RECT  1.040 -0.280 3.200 0.340 ;
        RECT  0.760 -0.280 1.040 0.760 ;
        RECT  0.000 -0.280 0.760 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.710 3.320 6.800 3.880 ;
        RECT  6.430 1.910 6.710 3.880 ;
        RECT  5.750 3.320 6.430 3.880 ;
        RECT  5.470 2.560 5.750 3.880 ;
        RECT  4.790 3.320 5.470 3.880 ;
        RECT  4.510 2.230 4.790 3.880 ;
        RECT  3.830 3.320 4.510 3.880 ;
        RECT  3.610 1.910 3.830 3.880 ;
        RECT  2.730 3.320 3.610 3.880 ;
        RECT  2.450 3.200 2.730 3.880 ;
        RECT  0.920 3.320 2.450 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.790 1.470 5.070 1.750 ;
        RECT  4.470 1.470 4.790 1.630 ;
        RECT  4.310 0.590 4.470 2.070 ;
        RECT  4.190 0.590 4.310 1.310 ;
        RECT  4.030 1.910 4.310 2.920 ;
        RECT  3.960 1.470 4.110 1.750 ;
        RECT  3.800 0.810 3.960 1.750 ;
        RECT  3.680 0.810 3.800 1.090 ;
        RECT  3.440 1.590 3.800 1.750 ;
        RECT  3.280 1.590 3.440 2.680 ;
        RECT  3.090 2.000 3.280 2.680 ;
        RECT  2.890 2.880 3.170 3.160 ;
        RECT  2.680 0.800 2.920 1.080 ;
        RECT  2.000 2.880 2.890 3.040 ;
        RECT  2.640 0.800 2.680 2.720 ;
        RECT  2.520 0.920 2.640 2.720 ;
        RECT  2.160 2.440 2.520 2.720 ;
        RECT  1.360 0.500 2.480 0.720 ;
        RECT  2.080 1.030 2.360 2.280 ;
        RECT  2.000 2.120 2.080 2.280 ;
        RECT  1.840 2.120 2.000 3.040 ;
        RECT  1.800 1.040 1.920 1.960 ;
        RECT  1.680 2.120 1.840 2.400 ;
        RECT  1.760 0.920 1.800 1.960 ;
        RECT  1.520 0.920 1.760 1.200 ;
        RECT  1.480 1.800 1.760 1.960 ;
        RECT  1.360 1.360 1.600 1.640 ;
        RECT  1.200 1.800 1.480 2.570 ;
        RECT  1.320 0.500 1.360 1.640 ;
        RECT  1.200 0.500 1.320 1.520 ;
        RECT  1.040 1.320 1.200 1.520 ;
        RECT  0.880 1.320 1.040 2.280 ;
        RECT  0.480 1.320 0.880 1.480 ;
        RECT  0.380 2.120 0.880 2.280 ;
        RECT  0.200 1.030 0.480 1.480 ;
        RECT  0.100 2.120 0.380 2.400 ;
    END
END CLKMX2X8TR

MACRO CLKMX2X6TR
    CLASS CORE ;
    FOREIGN CLKMX2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.490 1.840 7.770 3.160 ;
        RECT  7.060 1.840 7.490 2.650 ;
        RECT  6.810 0.440 7.060 2.650 ;
        RECT  6.700 0.440 6.810 3.160 ;
        RECT  6.530 2.040 6.700 3.160 ;
        END
        ANTENNADIFFAREA 5.772 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.240 0.730 1.630 ;
        END
        ANTENNAGATEAREA 0.6672 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.960 ;
        RECT  1.050 1.670 1.280 1.960 ;
        END
        ANTENNAGATEAREA 0.5016 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 1.240 5.960 1.560 ;
        END
        ANTENNAGATEAREA 0.4896 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.500 -0.280 8.000 0.280 ;
        RECT  7.220 -0.280 7.500 1.140 ;
        RECT  6.460 -0.280 7.220 0.280 ;
        RECT  6.180 -0.280 6.460 1.140 ;
        RECT  5.420 -0.280 6.180 0.280 ;
        RECT  5.140 -0.280 5.420 0.340 ;
        RECT  1.550 -0.280 5.140 0.280 ;
        RECT  0.610 -0.280 1.550 0.760 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.290 3.320 8.000 3.880 ;
        RECT  7.010 2.930 7.290 3.880 ;
        RECT  6.330 3.320 7.010 3.880 ;
        RECT  6.050 2.930 6.330 3.880 ;
        RECT  5.370 3.320 6.050 3.880 ;
        RECT  5.090 2.930 5.370 3.880 ;
        RECT  1.810 3.260 5.090 3.880 ;
        RECT  1.530 2.440 1.810 3.880 ;
        RECT  0.850 3.320 1.530 3.880 ;
        RECT  0.570 2.530 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.260 1.600 6.540 1.880 ;
        RECT  6.170 1.720 6.260 1.880 ;
        RECT  6.010 1.720 6.170 2.500 ;
        RECT  4.720 2.340 6.010 2.500 ;
        RECT  5.480 0.570 5.940 0.850 ;
        RECT  5.480 1.900 5.850 2.180 ;
        RECT  5.320 0.500 5.480 2.180 ;
        RECT  4.480 0.500 5.320 0.660 ;
        RECT  4.240 2.020 5.320 2.180 ;
        RECT  5.000 0.820 5.160 1.860 ;
        RECT  4.680 0.820 5.000 1.100 ;
        RECT  3.780 1.700 5.000 1.860 ;
        RECT  4.100 1.260 4.840 1.540 ;
        RECT  4.440 2.340 4.720 3.100 ;
        RECT  4.260 0.500 4.480 0.900 ;
        RECT  3.760 2.940 4.440 3.100 ;
        RECT  3.960 2.020 4.240 2.780 ;
        RECT  3.940 0.440 4.100 1.540 ;
        RECT  1.870 0.440 3.940 0.600 ;
        RECT  3.760 0.860 3.780 1.860 ;
        RECT  3.560 0.860 3.760 3.100 ;
        RECT  3.480 1.910 3.560 3.100 ;
        RECT  2.840 2.940 3.480 3.100 ;
        RECT  3.160 0.760 3.360 1.040 ;
        RECT  3.160 1.910 3.280 2.780 ;
        RECT  3.000 0.760 3.160 2.780 ;
        RECT  2.260 0.760 3.000 0.920 ;
        RECT  2.680 1.080 2.840 3.100 ;
        RECT  2.560 1.080 2.680 1.300 ;
        RECT  2.520 1.910 2.680 3.100 ;
        RECT  2.260 2.120 2.320 2.930 ;
        RECT  2.100 0.760 2.260 2.930 ;
        RECT  2.030 1.000 2.100 1.280 ;
        RECT  2.040 2.120 2.100 2.930 ;
        RECT  1.330 2.120 2.040 2.280 ;
        RECT  1.870 1.450 1.940 1.730 ;
        RECT  1.710 0.440 1.870 1.730 ;
        RECT  0.370 0.920 1.710 1.080 ;
        RECT  1.050 2.120 1.330 3.150 ;
        RECT  0.250 0.760 0.370 1.080 ;
        RECT  0.250 1.800 0.370 3.150 ;
        RECT  0.090 0.760 0.250 3.150 ;
    END
END CLKMX2X6TR

MACRO CLKMX2X4TR
    CLASS CORE ;
    FOREIGN CLKMX2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 0.580 3.890 2.360 ;
        RECT  3.410 0.580 3.570 1.340 ;
        RECT  3.520 2.120 3.570 2.360 ;
        RECT  3.140 2.120 3.520 3.160 ;
        END
        ANTENNADIFFAREA 3.564 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.440 0.720 2.920 ;
        END
        ANTENNAGATEAREA 0.2928 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.170 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.840 3.160 1.160 ;
        RECT  2.970 0.840 3.040 1.480 ;
        RECT  2.880 0.840 2.970 1.640 ;
        RECT  2.690 1.320 2.880 1.640 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.210 -0.280 4.000 0.280 ;
        RECT  2.930 -0.280 3.210 0.680 ;
        RECT  0.870 -0.280 2.930 0.280 ;
        RECT  0.650 -0.280 0.870 0.760 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.900 3.320 4.000 3.880 ;
        RECT  3.680 2.520 3.900 3.880 ;
        RECT  2.940 3.320 3.680 3.880 ;
        RECT  2.660 2.930 2.940 3.880 ;
        RECT  0.890 3.320 2.660 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 1.680 3.410 1.960 ;
        RECT  2.850 1.800 3.130 1.960 ;
        RECT  2.690 1.800 2.850 2.740 ;
        RECT  2.530 0.880 2.690 1.160 ;
        RECT  1.930 2.580 2.690 2.740 ;
        RECT  2.370 0.880 2.530 2.420 ;
        RECT  1.830 0.440 2.490 0.660 ;
        RECT  2.180 2.200 2.370 2.420 ;
        RECT  1.990 1.120 2.210 2.040 ;
        RECT  1.930 1.880 1.990 2.040 ;
        RECT  1.890 1.880 1.930 2.740 ;
        RECT  1.770 1.880 1.890 3.160 ;
        RECT  1.670 0.440 1.830 1.720 ;
        RECT  1.610 2.030 1.770 3.160 ;
        RECT  1.190 0.440 1.670 0.600 ;
        RECT  1.610 1.560 1.670 1.720 ;
        RECT  1.330 1.560 1.610 1.870 ;
        RECT  1.350 1.120 1.510 1.400 ;
        RECT  1.130 2.120 1.410 3.160 ;
        RECT  0.720 1.240 1.350 1.400 ;
        RECT  1.030 0.440 1.190 1.080 ;
        RECT  0.720 2.120 1.130 2.280 ;
        RECT  0.250 0.920 1.030 1.080 ;
        RECT  0.560 1.240 0.720 2.280 ;
        RECT  0.250 2.030 0.400 2.250 ;
        RECT  0.090 0.920 0.250 2.250 ;
    END
END CLKMX2X4TR

MACRO CLKMX2X3TR
    CLASS CORE ;
    FOREIGN CLKMX2X3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 0.760 3.660 1.310 ;
        RECT  3.200 0.760 3.480 2.720 ;
        END
        ANTENNADIFFAREA 2.712 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 2.440 0.730 2.760 ;
        END
        ANTENNAGATEAREA 0.3 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.640 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.2136 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.640 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2136 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.280 4.000 0.280 ;
        RECT  2.860 -0.280 3.140 0.460 ;
        RECT  0.840 -0.280 2.860 0.340 ;
        RECT  0.560 -0.280 0.840 0.750 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.880 3.320 4.000 3.880 ;
        RECT  2.800 3.200 3.880 3.880 ;
        RECT  0.840 3.320 2.800 3.880 ;
        RECT  0.560 2.930 0.840 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.800 1.640 3.920 1.920 ;
        RECT  3.640 1.640 3.800 3.040 ;
        RECT  2.080 2.880 3.640 3.040 ;
        RECT  2.880 1.150 3.040 2.280 ;
        RECT  2.600 1.150 2.880 1.310 ;
        RECT  2.560 2.120 2.880 2.280 ;
        RECT  2.320 1.030 2.600 1.310 ;
        RECT  2.280 2.120 2.560 2.630 ;
        RECT  1.200 0.500 2.370 0.660 ;
        RECT  1.920 0.920 2.080 3.040 ;
        RECT  1.860 2.560 1.920 3.040 ;
        RECT  1.500 2.560 1.860 3.120 ;
        RECT  1.600 0.880 1.760 2.280 ;
        RECT  1.360 0.880 1.600 1.160 ;
        RECT  1.340 2.120 1.600 2.280 ;
        RECT  1.280 1.320 1.440 1.920 ;
        RECT  1.070 2.120 1.340 3.160 ;
        RECT  1.200 1.320 1.280 1.480 ;
        RECT  1.040 0.500 1.200 1.480 ;
        RECT  0.400 1.320 1.040 1.480 ;
        RECT  0.280 2.070 0.440 2.240 ;
        RECT  0.280 1.030 0.400 1.480 ;
        RECT  0.120 1.030 0.280 2.240 ;
    END
END CLKMX2X3TR

MACRO CLKMX2X2TR
    CLASS CORE ;
    FOREIGN CLKMX2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 1.030 3.520 3.160 ;
        RECT  3.200 1.030 3.360 1.310 ;
        RECT  3.200 1.930 3.360 3.160 ;
        END
        ANTENNADIFFAREA 2.816 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.360 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.140 1.140 1.560 ;
        END
        ANTENNAGATEAREA 0.1656 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.210 2.720 1.670 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 -0.280 3.600 0.280 ;
        RECT  2.760 -0.280 3.040 0.350 ;
        RECT  0.930 -0.280 2.760 0.340 ;
        RECT  0.650 -0.280 0.930 0.940 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 3.320 3.600 3.880 ;
        RECT  2.720 2.670 3.000 3.880 ;
        RECT  0.970 3.260 2.720 3.880 ;
        RECT  0.690 2.500 0.970 3.880 ;
        RECT  0.000 3.320 0.690 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.040 1.470 3.200 1.750 ;
        RECT  2.880 0.510 3.040 2.470 ;
        RECT  1.960 0.510 2.880 0.670 ;
        RECT  2.280 2.310 2.880 2.470 ;
        RECT  2.280 0.830 2.440 1.050 ;
        RECT  2.280 1.930 2.410 2.150 ;
        RECT  2.120 0.830 2.280 2.150 ;
        RECT  2.120 2.310 2.280 2.520 ;
        RECT  1.930 2.360 2.120 2.520 ;
        RECT  1.760 0.510 1.960 0.950 ;
        RECT  1.800 1.110 1.960 2.200 ;
        RECT  1.650 2.360 1.930 2.640 ;
        RECT  1.520 1.110 1.800 1.270 ;
        RECT  1.450 2.040 1.800 2.200 ;
        RECT  1.680 0.670 1.760 0.950 ;
        RECT  1.360 1.430 1.640 1.880 ;
        RECT  1.360 0.670 1.520 1.270 ;
        RECT  1.290 2.040 1.450 2.720 ;
        RECT  1.170 0.670 1.360 0.950 ;
        RECT  1.080 1.720 1.360 1.880 ;
        RECT  1.170 2.440 1.290 2.720 ;
        RECT  0.920 1.720 1.080 2.280 ;
        RECT  0.320 2.120 0.920 2.280 ;
        RECT  0.160 0.720 0.320 2.280 ;
        RECT  0.090 0.720 0.160 1.070 ;
        RECT  0.100 2.000 0.160 2.280 ;
    END
END CLKMX2X2TR

MACRO CLKMX2X12TR
    CLASS CORE ;
    FOREIGN CLKMX2X12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.460 1.030 7.740 3.160 ;
        RECT  6.780 1.030 7.460 1.760 ;
        RECT  6.500 0.500 6.780 3.160 ;
        RECT  6.070 0.770 6.500 2.400 ;
        RECT  5.820 0.770 6.070 1.370 ;
        RECT  5.820 1.910 6.070 2.400 ;
        RECT  5.540 0.440 5.820 1.370 ;
        RECT  5.540 1.910 5.820 3.160 ;
        END
        ANTENNADIFFAREA 9.986 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 2.440 0.720 2.780 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.440 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.240 3.160 1.620 ;
        END
        ANTENNAGATEAREA 0.168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.300 -0.280 8.400 0.280 ;
        RECT  6.020 -0.280 6.300 0.610 ;
        RECT  5.340 -0.280 6.020 0.280 ;
        RECT  5.060 -0.280 5.340 1.310 ;
        RECT  4.340 -0.280 5.060 0.280 ;
        RECT  4.060 -0.280 4.340 1.020 ;
        RECT  3.400 -0.280 4.060 0.340 ;
        RECT  3.120 -0.280 3.400 1.080 ;
        RECT  1.040 -0.280 3.120 0.280 ;
        RECT  0.760 -0.280 1.040 0.960 ;
        RECT  0.000 -0.280 0.760 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.220 3.320 8.400 3.880 ;
        RECT  7.940 1.910 8.220 3.880 ;
        RECT  7.260 3.320 7.940 3.880 ;
        RECT  6.980 1.920 7.260 3.880 ;
        RECT  6.300 3.320 6.980 3.880 ;
        RECT  6.020 2.560 6.300 3.880 ;
        RECT  5.340 3.320 6.020 3.880 ;
        RECT  5.060 1.910 5.340 3.880 ;
        RECT  4.340 3.320 5.060 3.880 ;
        RECT  4.060 3.200 4.340 3.880 ;
        RECT  2.960 3.320 4.060 3.880 ;
        RECT  2.680 3.200 2.960 3.880 ;
        RECT  1.040 3.260 2.680 3.880 ;
        RECT  0.760 3.200 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 1.530 5.890 1.750 ;
        RECT  4.700 1.030 4.860 3.160 ;
        RECT  4.540 1.030 4.700 1.310 ;
        RECT  4.580 1.910 4.700 3.160 ;
        RECT  3.940 1.910 4.580 2.070 ;
        RECT  4.100 1.470 4.370 1.750 ;
        RECT  3.880 1.470 4.100 1.630 ;
        RECT  3.660 1.910 3.940 2.470 ;
        RECT  3.720 0.900 3.880 1.630 ;
        RECT  3.600 0.900 3.720 1.180 ;
        RECT  3.480 1.470 3.720 1.630 ;
        RECT  3.120 2.880 3.690 3.160 ;
        RECT  3.320 1.470 3.480 2.590 ;
        RECT  3.200 1.910 3.320 2.590 ;
        RECT  2.120 2.880 3.120 3.040 ;
        RECT  2.680 0.800 2.840 1.080 ;
        RECT  2.560 0.800 2.680 2.720 ;
        RECT  1.440 0.480 2.560 0.640 ;
        RECT  2.520 0.920 2.560 2.720 ;
        RECT  2.280 2.440 2.520 2.720 ;
        RECT  2.140 0.900 2.360 2.280 ;
        RECT  2.120 2.120 2.140 2.280 ;
        RECT  1.760 2.120 2.120 3.040 ;
        RECT  1.880 1.020 1.980 1.960 ;
        RECT  1.820 0.900 1.880 1.960 ;
        RECT  1.600 0.900 1.820 1.180 ;
        RECT  1.560 1.800 1.820 1.960 ;
        RECT  1.440 1.340 1.660 1.640 ;
        RECT  1.280 1.800 1.560 2.930 ;
        RECT  1.280 0.480 1.440 1.500 ;
        RECT  0.480 1.120 1.280 1.280 ;
        RECT  0.360 1.910 0.520 2.190 ;
        RECT  0.360 0.900 0.480 1.280 ;
        RECT  0.200 0.900 0.360 2.190 ;
    END
END CLKMX2X12TR

MACRO CLKINVX8TR
    CLASS CORE ;
    FOREIGN CLKINVX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.920 1.920 1.210 ;
        RECT  1.650 0.920 1.850 3.080 ;
        RECT  1.570 1.040 1.650 3.080 ;
        RECT  0.890 1.040 1.570 1.760 ;
        RECT  0.610 0.800 0.890 3.160 ;
        END
        ANTENNADIFFAREA 6.334 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.360 0.450 1.680 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.8352 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 -0.280 2.800 0.280 ;
        RECT  2.170 -0.280 2.450 1.230 ;
        RECT  1.410 -0.280 2.170 0.280 ;
        RECT  1.130 -0.280 1.410 0.760 ;
        RECT  0.370 -0.280 1.130 0.280 ;
        RECT  0.090 -0.280 0.370 0.680 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 3.320 2.800 3.880 ;
        RECT  2.050 1.910 2.330 3.880 ;
        RECT  1.370 3.320 2.050 3.880 ;
        RECT  1.090 2.040 1.370 3.880 ;
        RECT  0.410 3.320 1.090 3.880 ;
        RECT  0.130 2.190 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
END CLKINVX8TR

MACRO CLKINVX6TR
    CLASS CORE ;
    FOREIGN CLKINVX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.210 1.900 3.080 ;
        RECT  1.610 0.710 1.890 3.080 ;
        RECT  1.050 0.710 1.610 2.160 ;
        RECT  0.570 0.710 1.050 1.080 ;
        RECT  0.850 1.800 1.050 2.160 ;
        RECT  0.570 1.800 0.850 3.160 ;
        END
        ANTENNADIFFAREA 5.96 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.240 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.6312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.370 -0.280 2.000 0.280 ;
        RECT  0.090 -0.280 0.370 1.070 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.380 3.320 2.000 3.880 ;
        RECT  1.070 2.350 1.380 3.880 ;
        RECT  0.370 3.320 1.070 3.880 ;
        RECT  0.090 1.910 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END CLKINVX6TR

MACRO CLKINVX4TR
    CLASS CORE ;
    FOREIGN CLKINVX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.940 0.800 1.120 2.160 ;
        RECT  0.880 0.800 0.940 3.020 ;
        RECT  0.660 0.800 0.880 1.080 ;
        RECT  0.660 1.910 0.880 3.020 ;
        END
        ANTENNADIFFAREA 3.132 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.720 1.630 ;
        END
        ANTENNAGATEAREA 0.4176 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.450 -0.280 1.600 0.280 ;
        RECT  1.280 -0.280 1.450 1.060 ;
        RECT  0.420 -0.280 1.280 0.340 ;
        RECT  0.140 -0.280 0.420 1.080 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 3.320 1.600 3.880 ;
        RECT  1.180 2.400 1.460 3.880 ;
        RECT  0.460 3.320 1.180 3.880 ;
        RECT  0.180 1.910 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
END CLKINVX4TR

MACRO CLKINVX3TR
    CLASS CORE ;
    FOREIGN CLKINVX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.600 1.120 2.160 ;
        RECT  0.940 0.800 1.060 2.160 ;
        RECT  0.880 0.800 0.940 2.660 ;
        RECT  0.660 0.800 0.880 1.080 ;
        RECT  0.660 1.910 0.880 2.660 ;
        END
        ANTENNADIFFAREA 2.394 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.720 1.630 ;
        END
        ANTENNAGATEAREA 0.3192 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.510 -0.280 1.600 0.280 ;
        RECT  1.220 -0.280 1.510 1.100 ;
        RECT  0.420 -0.280 1.220 0.340 ;
        RECT  0.140 -0.280 0.420 1.080 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 3.320 1.600 3.880 ;
        RECT  1.180 2.400 1.460 3.880 ;
        RECT  0.460 3.320 1.180 3.880 ;
        RECT  0.180 1.910 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
END CLKINVX3TR

MACRO CLKINVX2TR
    CLASS CORE ;
    FOREIGN CLKINVX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 0.440 1.120 1.560 ;
        RECT  0.950 0.440 1.110 3.100 ;
        RECT  0.880 0.440 0.950 1.560 ;
        RECT  0.790 2.400 0.950 3.100 ;
        RECT  0.800 0.840 0.880 1.160 ;
        END
        ANTENNADIFFAREA 2.848 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2136 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 -0.280 1.200 0.280 ;
        RECT  0.270 -0.280 0.550 1.250 ;
        RECT  0.000 -0.280 0.270 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 3.320 1.200 3.880 ;
        RECT  0.250 2.350 0.550 3.880 ;
        RECT  0.000 3.320 0.250 3.880 ;
        END
    END VDD
END CLKINVX2TR

MACRO CLKINVX20TR
    CLASS CORE ;
    FOREIGN CLKINVX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 0.650 4.720 2.830 ;
        RECT  3.740 1.000 4.420 2.370 ;
        RECT  3.460 0.540 3.740 3.160 ;
        RECT  2.780 1.000 3.460 2.200 ;
        RECT  2.500 0.540 2.780 3.160 ;
        RECT  1.820 1.000 2.500 2.200 ;
        RECT  1.540 0.570 1.820 3.160 ;
        RECT  0.870 1.000 1.540 2.200 ;
        RECT  0.860 0.630 0.870 2.200 ;
        RECT  0.580 0.630 0.860 2.890 ;
        END
        ANTENNADIFFAREA 16.1 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.420 1.640 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 2.0832 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.180 -0.280 5.600 0.280 ;
        RECT  4.900 -0.280 5.180 1.060 ;
        RECT  4.220 -0.280 4.900 0.280 ;
        RECT  3.940 -0.280 4.220 0.770 ;
        RECT  3.260 -0.280 3.940 0.280 ;
        RECT  2.980 -0.280 3.260 0.760 ;
        RECT  2.300 -0.280 2.980 0.280 ;
        RECT  2.020 -0.280 2.300 0.760 ;
        RECT  1.340 -0.280 2.020 0.280 ;
        RECT  1.060 -0.280 1.340 0.760 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 1.060 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.200 3.320 5.600 3.880 ;
        RECT  4.900 2.020 5.200 3.880 ;
        RECT  4.220 3.320 4.900 3.880 ;
        RECT  3.940 2.570 4.220 3.880 ;
        RECT  3.260 3.320 3.940 3.880 ;
        RECT  2.980 2.480 3.260 3.880 ;
        RECT  2.300 3.320 2.980 3.880 ;
        RECT  2.020 2.490 2.300 3.880 ;
        RECT  1.340 3.320 2.020 3.880 ;
        RECT  1.060 2.480 1.340 3.880 ;
        RECT  0.380 3.320 1.060 3.880 ;
        RECT  0.100 2.530 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
END CLKINVX20TR

MACRO CLKINVX1TR
    CLASS CORE ;
    FOREIGN CLKINVX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.840 1.120 2.470 ;
        RECT  0.770 1.070 0.880 1.310 ;
        RECT  0.730 2.170 0.880 2.470 ;
        END
        ANTENNADIFFAREA 1.526 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.520 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 -0.280 1.200 0.280 ;
        RECT  0.210 -0.280 0.490 1.310 ;
        RECT  0.000 -0.280 0.210 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 3.320 1.200 3.880 ;
        RECT  0.210 2.170 0.520 3.880 ;
        RECT  0.000 3.320 0.210 3.880 ;
        END
    END VDD
END CLKINVX1TR

MACRO CLKINVX16TR
    CLASS CORE ;
    FOREIGN CLKINVX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.440 4.580 2.820 ;
        RECT  1.020 0.500 3.280 1.370 ;
        RECT  1.060 1.850 3.280 2.820 ;
        END
        ANTENNADIFFAREA 12.762 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.530 3.120 1.690 ;
        RECT  0.480 1.530 0.720 1.960 ;
        END
        ANTENNAGATEAREA 1.7016 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 -0.280 4.800 0.280 ;
        RECT  2.580 -0.280 2.860 0.340 ;
        RECT  1.820 -0.280 2.580 0.280 ;
        RECT  1.540 -0.280 1.820 0.340 ;
        RECT  0.820 -0.280 1.540 0.280 ;
        RECT  0.540 -0.280 0.820 1.220 ;
        RECT  0.000 -0.280 0.540 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.420 2.990 4.700 3.880 ;
        RECT  3.740 3.320 4.420 3.880 ;
        RECT  3.460 2.990 3.740 3.880 ;
        RECT  2.780 3.320 3.460 3.880 ;
        RECT  2.500 2.990 2.780 3.880 ;
        RECT  1.820 3.320 2.500 3.880 ;
        RECT  1.540 2.990 1.820 3.880 ;
        RECT  0.860 3.320 1.540 3.880 ;
        RECT  0.580 2.280 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
END CLKINVX16TR

MACRO CLKINVX12TR
    CLASS CORE ;
    FOREIGN CLKINVX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 0.660 3.350 3.020 ;
        RECT  2.390 1.010 3.070 1.770 ;
        RECT  2.320 1.010 2.390 3.030 ;
        RECT  2.110 0.650 2.320 3.030 ;
        RECT  2.030 0.650 2.110 1.740 ;
        RECT  1.430 1.010 2.030 1.740 ;
        RECT  1.350 1.010 1.430 3.010 ;
        RECT  1.150 0.590 1.350 3.010 ;
        RECT  1.070 0.590 1.150 0.910 ;
        END
        ANTENNADIFFAREA 9.396 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.100 0.990 1.600 ;
        END
        ANTENNAGATEAREA 1.2528 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.280 4.000 0.280 ;
        RECT  3.590 -0.280 3.870 0.400 ;
        RECT  2.830 -0.280 3.590 0.280 ;
        RECT  2.550 -0.280 2.830 0.400 ;
        RECT  1.840 -0.280 2.550 0.280 ;
        RECT  1.550 -0.280 1.840 0.820 ;
        RECT  0.840 -0.280 1.550 0.280 ;
        RECT  0.550 -0.280 0.840 0.900 ;
        RECT  0.000 -0.280 0.550 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 3.320 4.000 3.880 ;
        RECT  3.550 2.040 3.830 3.880 ;
        RECT  2.870 3.320 3.550 3.880 ;
        RECT  2.590 2.140 2.870 3.880 ;
        RECT  1.910 3.320 2.590 3.880 ;
        RECT  1.630 2.110 1.910 3.880 ;
        RECT  0.950 3.320 1.630 3.880 ;
        RECT  0.670 2.050 0.950 3.880 ;
        RECT  0.000 3.320 0.670 3.880 ;
        END
    END VDD
END CLKINVX12TR

MACRO CLKBUFX8TR
    CLASS CORE ;
    FOREIGN CLKBUFX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 1.040 2.850 3.160 ;
        RECT  1.850 1.040 2.570 1.760 ;
        RECT  1.810 0.440 1.850 1.760 ;
        RECT  1.550 0.440 1.810 3.160 ;
        RECT  1.530 1.910 1.550 3.160 ;
        END
        ANTENNADIFFAREA 6.264 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.400 1.050 1.640 ;
        RECT  0.080 0.440 0.330 1.640 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.280 3.600 0.280 ;
        RECT  2.050 -0.280 2.330 0.670 ;
        RECT  1.370 -0.280 2.050 0.280 ;
        RECT  1.090 -0.280 1.370 0.760 ;
        RECT  0.000 -0.280 1.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 3.320 3.600 3.880 ;
        RECT  3.050 1.910 3.330 3.880 ;
        RECT  2.330 3.320 3.050 3.880 ;
        RECT  2.050 2.030 2.330 3.880 ;
        RECT  1.330 3.320 2.050 3.880 ;
        RECT  1.050 2.120 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 1.990 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.370 1.470 1.390 1.750 ;
        RECT  1.210 0.920 1.370 1.960 ;
        RECT  0.810 0.920 1.210 1.080 ;
        RECT  0.850 1.800 1.210 1.960 ;
        RECT  0.690 1.800 0.850 2.800 ;
        RECT  0.530 0.710 0.810 1.080 ;
        RECT  0.570 1.990 0.690 2.800 ;
    END
END CLKBUFX8TR

MACRO CLKBUFX6TR
    CLASS CORE ;
    FOREIGN CLKBUFX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.440 2.640 3.100 ;
        RECT  1.680 1.440 2.360 2.160 ;
        RECT  1.480 0.890 1.680 3.160 ;
        RECT  1.400 0.890 1.480 1.350 ;
        RECT  1.400 2.060 1.480 3.160 ;
        END
        ANTENNADIFFAREA 5.63 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.840 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 -0.280 2.800 0.280 ;
        RECT  1.920 -0.280 2.200 1.080 ;
        RECT  1.160 -0.280 1.920 0.280 ;
        RECT  0.880 -0.280 1.160 0.760 ;
        RECT  0.000 -0.280 0.880 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 3.320 2.800 3.880 ;
        RECT  1.880 2.480 2.160 3.880 ;
        RECT  1.200 3.320 1.880 3.880 ;
        RECT  0.920 2.340 1.200 3.880 ;
        RECT  0.000 3.320 0.920 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.160 1.560 1.270 1.840 ;
        RECT  1.000 0.920 1.160 2.070 ;
        RECT  0.640 0.920 1.000 1.080 ;
        RECT  0.720 1.910 1.000 2.070 ;
        RECT  0.440 1.910 0.720 3.040 ;
        RECT  0.360 0.800 0.640 1.080 ;
    END
END CLKBUFX6TR

MACRO CLKBUFX4TR
    CLASS CORE ;
    FOREIGN CLKBUFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.940 1.980 1.900 ;
        RECT  1.510 0.940 1.740 1.110 ;
        RECT  1.520 1.660 1.740 1.900 ;
        RECT  1.230 1.660 1.520 3.160 ;
        RECT  1.230 0.840 1.510 1.110 ;
        END
        ANTENNADIFFAREA 3.132 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.720 1.560 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 -0.280 2.400 0.280 ;
        RECT  1.750 -0.280 2.030 0.740 ;
        RECT  0.990 -0.280 1.750 0.340 ;
        RECT  0.710 -0.280 0.990 0.760 ;
        RECT  0.000 -0.280 0.710 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 3.320 2.400 3.880 ;
        RECT  1.750 2.060 2.030 3.880 ;
        RECT  0.990 3.320 1.750 3.880 ;
        RECT  0.710 2.040 0.990 3.880 ;
        RECT  0.000 3.320 0.710 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 1.270 1.540 1.500 ;
        RECT  0.880 0.920 1.040 1.880 ;
        RECT  0.470 0.920 0.880 1.080 ;
        RECT  0.470 1.720 0.880 1.880 ;
        RECT  0.190 0.800 0.470 1.080 ;
        RECT  0.190 1.720 0.470 2.710 ;
    END
END CLKBUFX4TR

MACRO CLKBUFX3TR
    CLASS CORE ;
    FOREIGN CLKBUFX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.000 1.920 2.160 ;
        RECT  1.570 1.000 1.760 1.160 ;
        RECT  1.430 2.000 1.760 2.160 ;
        RECT  1.240 0.840 1.570 1.160 ;
        RECT  1.150 2.000 1.430 2.880 ;
        END
        ANTENNADIFFAREA 2.898 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.790 ;
        END
        ANTENNAGATEAREA 0.0984 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.280 2.000 0.280 ;
        RECT  0.720 -0.280 1.000 0.400 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.630 2.470 1.910 3.880 ;
        RECT  0.950 3.320 1.630 3.880 ;
        RECT  0.670 2.160 0.950 3.880 ;
        RECT  0.000 3.320 0.670 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 1.560 1.570 1.840 ;
        RECT  0.920 0.920 1.080 1.840 ;
        RECT  0.440 0.920 0.920 1.080 ;
        RECT  0.320 0.800 0.440 1.080 ;
        RECT  0.160 0.800 0.320 2.560 ;
    END
END CLKBUFX3TR

MACRO CLKBUFX2TR
    CLASS CORE ;
    FOREIGN CLKBUFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.840 1.520 2.940 ;
        RECT  1.280 0.840 1.350 1.960 ;
        RECT  1.230 2.230 1.350 2.940 ;
        RECT  1.200 0.840 1.280 1.220 ;
        END
        ANTENNADIFFAREA 2.848 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.240 0.720 1.560 ;
        RECT  0.480 1.240 0.680 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.0888 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.280 1.600 0.280 ;
        RECT  0.720 -0.280 1.000 1.080 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 3.320 1.600 3.880 ;
        RECT  0.750 2.230 1.030 3.880 ;
        RECT  0.000 3.320 0.750 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 1.520 1.120 2.070 ;
        RECT  0.530 1.910 0.950 2.070 ;
        RECT  0.240 1.910 0.530 2.350 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.230 1.030 0.240 2.350 ;
        RECT  0.080 1.030 0.230 2.070 ;
    END
END CLKBUFX2TR

MACRO CLKBUFX20TR
    CLASS CORE ;
    FOREIGN CLKBUFX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.520 0.440 6.730 1.560 ;
        RECT  5.680 0.440 6.520 2.820 ;
        RECT  5.400 0.500 5.680 2.820 ;
        RECT  2.360 0.500 5.400 1.370 ;
        RECT  2.400 1.850 5.400 2.820 ;
        END
        ANTENNADIFFAREA 15.966 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.460 1.400 1.780 ;
        RECT  0.480 1.460 0.770 1.960 ;
        END
        ANTENNAGATEAREA 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 -0.280 7.200 0.280 ;
        RECT  4.960 -0.280 5.240 0.340 ;
        RECT  4.200 -0.280 4.960 0.280 ;
        RECT  3.920 -0.280 4.200 0.340 ;
        RECT  3.160 -0.280 3.920 0.280 ;
        RECT  2.880 -0.280 3.160 0.340 ;
        RECT  2.160 -0.280 2.880 0.280 ;
        RECT  1.880 -0.280 2.160 0.980 ;
        RECT  1.200 -0.280 1.880 0.280 ;
        RECT  0.920 -0.280 1.200 0.980 ;
        RECT  0.000 -0.280 0.920 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.000 3.320 7.200 3.880 ;
        RECT  6.720 1.910 7.000 3.880 ;
        RECT  6.040 3.320 6.720 3.880 ;
        RECT  5.760 2.990 6.040 3.880 ;
        RECT  5.080 3.320 5.760 3.880 ;
        RECT  4.800 2.990 5.080 3.880 ;
        RECT  4.120 3.320 4.800 3.880 ;
        RECT  3.840 2.990 4.120 3.880 ;
        RECT  3.160 3.320 3.840 3.880 ;
        RECT  2.880 2.990 3.160 3.880 ;
        RECT  2.200 3.320 2.880 3.880 ;
        RECT  1.920 1.910 2.200 3.880 ;
        RECT  1.240 3.320 1.920 3.880 ;
        RECT  0.960 2.650 1.240 3.880 ;
        RECT  0.000 3.320 0.960 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 1.530 5.240 1.690 ;
        RECT  1.680 1.140 1.720 2.890 ;
        RECT  1.560 0.700 1.680 2.890 ;
        RECT  1.400 0.700 1.560 1.300 ;
        RECT  1.440 2.210 1.560 2.890 ;
        RECT  0.760 2.210 1.440 2.370 ;
        RECT  0.720 1.140 1.400 1.300 ;
        RECT  0.480 2.210 0.760 2.860 ;
        RECT  0.440 0.700 0.720 1.300 ;
    END
END CLKBUFX20TR

MACRO CLKBUFX16TR
    CLASS CORE ;
    FOREIGN CLKBUFX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 0.440 5.580 2.820 ;
        RECT  2.020 0.500 4.480 1.370 ;
        RECT  2.060 1.850 4.480 2.820 ;
        END
        ANTENNADIFFAREA 12.762 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.510 1.060 1.780 ;
        RECT  0.390 1.510 0.780 1.960 ;
        END
        ANTENNAGATEAREA 0.5424 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.860 -0.280 6.000 0.280 ;
        RECT  3.580 -0.280 3.860 0.340 ;
        RECT  2.820 -0.280 3.580 0.280 ;
        RECT  2.540 -0.280 2.820 0.340 ;
        RECT  1.820 -0.280 2.540 0.280 ;
        RECT  1.540 -0.280 1.820 1.220 ;
        RECT  0.860 -0.280 1.540 0.280 ;
        RECT  0.580 -0.280 0.860 1.030 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.700 3.320 6.000 3.880 ;
        RECT  5.420 2.990 5.700 3.880 ;
        RECT  4.740 3.320 5.420 3.880 ;
        RECT  4.460 2.990 4.740 3.880 ;
        RECT  3.780 3.320 4.460 3.880 ;
        RECT  3.500 2.990 3.780 3.880 ;
        RECT  2.820 3.320 3.500 3.880 ;
        RECT  2.540 2.990 2.820 3.880 ;
        RECT  1.860 3.320 2.540 3.880 ;
        RECT  1.580 1.910 1.860 3.880 ;
        RECT  0.900 3.320 1.580 3.880 ;
        RECT  0.620 2.650 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.380 1.530 4.180 1.690 ;
        RECT  1.220 0.800 1.380 2.890 ;
        RECT  1.060 0.800 1.220 1.350 ;
        RECT  1.100 2.210 1.220 2.890 ;
        RECT  0.420 2.210 1.100 2.370 ;
        RECT  0.380 1.190 1.060 1.350 ;
        RECT  0.140 2.210 0.420 2.860 ;
        RECT  0.100 0.700 0.380 1.350 ;
    END
END CLKBUFX16TR

MACRO CLKBUFX12TR
    CLASS CORE ;
    FOREIGN CLKBUFX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.660 4.150 3.020 ;
        RECT  3.190 1.010 3.870 1.770 ;
        RECT  3.120 1.010 3.190 3.030 ;
        RECT  2.910 0.650 3.120 3.030 ;
        RECT  2.830 0.650 2.910 1.740 ;
        RECT  2.230 1.010 2.830 1.740 ;
        RECT  2.150 1.010 2.230 3.010 ;
        RECT  1.950 0.590 2.150 3.010 ;
        RECT  1.870 0.590 1.950 0.910 ;
        END
        ANTENNADIFFAREA 9.396 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.470 0.920 1.720 ;
        RECT  0.480 1.240 0.720 1.720 ;
        END
        ANTENNAGATEAREA 0.4008 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.670 -0.280 4.800 0.280 ;
        RECT  4.390 -0.280 4.670 0.400 ;
        RECT  3.630 -0.280 4.390 0.280 ;
        RECT  3.350 -0.280 3.630 0.400 ;
        RECT  2.640 -0.280 3.350 0.280 ;
        RECT  2.350 -0.280 2.640 0.820 ;
        RECT  1.640 -0.280 2.350 0.280 ;
        RECT  1.350 -0.280 1.640 0.900 ;
        RECT  0.000 -0.280 1.350 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.630 3.320 4.800 3.880 ;
        RECT  4.350 2.040 4.630 3.880 ;
        RECT  3.670 3.320 4.350 3.880 ;
        RECT  3.390 2.140 3.670 3.880 ;
        RECT  2.710 3.320 3.390 3.880 ;
        RECT  2.430 2.110 2.710 3.880 ;
        RECT  1.750 3.320 2.430 3.880 ;
        RECT  1.470 2.050 1.750 3.880 ;
        RECT  0.790 3.320 1.470 3.880 ;
        RECT  0.530 1.970 0.790 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.280 1.100 1.790 1.370 ;
        RECT  1.270 1.100 1.280 1.670 ;
        RECT  1.150 1.100 1.270 2.990 ;
        RECT  1.080 0.490 1.150 2.990 ;
        RECT  0.920 0.490 1.080 1.310 ;
        RECT  0.990 2.010 1.080 2.990 ;
    END
END CLKBUFX12TR

MACRO CLKAND2X8TR
    CLASS CORE ;
    FOREIGN CLKAND2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 1.040 3.840 3.160 ;
        RECT  3.280 1.040 3.480 1.760 ;
        RECT  3.000 0.670 3.280 1.760 ;
        RECT  2.800 0.750 3.000 1.760 ;
        RECT  2.520 0.750 2.800 3.160 ;
        RECT  2.320 0.750 2.520 1.060 ;
        RECT  2.040 0.670 2.320 1.060 ;
        END
        ANTENNADIFFAREA 7.04 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.640 2.020 1.900 ;
        RECT  0.760 1.740 1.720 1.900 ;
        RECT  0.480 1.240 0.760 1.900 ;
        RECT  0.380 1.240 0.480 1.600 ;
        END
        ANTENNAGATEAREA 0.336 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.240 1.560 1.580 ;
        END
        ANTENNAGATEAREA 0.336 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.760 -0.280 4.000 0.280 ;
        RECT  3.480 -0.280 3.760 0.650 ;
        RECT  2.800 -0.280 3.480 0.280 ;
        RECT  2.520 -0.280 2.800 0.590 ;
        RECT  0.880 -0.280 2.520 0.280 ;
        RECT  0.600 -0.280 0.880 1.080 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 3.320 4.000 3.880 ;
        RECT  3.000 2.080 3.280 3.880 ;
        RECT  2.300 3.320 3.000 3.880 ;
        RECT  2.020 2.660 2.300 3.880 ;
        RECT  1.340 3.320 2.020 3.880 ;
        RECT  1.060 2.660 1.340 3.880 ;
        RECT  0.320 3.320 1.060 3.880 ;
        RECT  0.100 2.200 0.320 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.180 1.220 2.340 2.220 ;
        RECT  1.880 1.220 2.180 1.380 ;
        RECT  1.820 2.060 2.180 2.220 ;
        RECT  1.720 0.630 1.880 1.380 ;
        RECT  1.540 2.060 1.820 2.940 ;
        RECT  1.680 0.630 1.720 0.790 ;
        RECT  1.400 0.510 1.680 0.790 ;
        RECT  0.860 2.060 1.540 2.220 ;
        RECT  0.580 2.060 0.860 2.940 ;
    END
END CLKAND2X8TR

MACRO CLKAND2X6TR
    CLASS CORE ;
    FOREIGN CLKAND2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.030 2.920 2.800 ;
        RECT  1.880 1.030 2.640 1.770 ;
        RECT  1.620 0.520 1.880 2.820 ;
        RECT  1.600 0.520 1.620 0.930 ;
        RECT  1.600 1.640 1.620 2.820 ;
        END
        ANTENNADIFFAREA 4.526 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.200 1.120 1.560 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.090 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2112 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.280 3.200 0.280 ;
        RECT  2.120 -0.280 2.400 0.720 ;
        RECT  0.000 -0.280 2.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 3.320 3.200 3.880 ;
        RECT  2.120 2.280 2.400 3.880 ;
        RECT  1.400 3.320 2.120 3.880 ;
        RECT  1.120 2.040 1.400 3.880 ;
        RECT  0.440 3.320 1.120 3.880 ;
        RECT  0.160 2.550 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.200 1.460 1.480 ;
        RECT  1.280 0.770 1.440 1.880 ;
        RECT  0.440 0.770 1.280 0.930 ;
        RECT  0.920 1.720 1.280 1.880 ;
        RECT  0.640 1.720 0.920 2.950 ;
        RECT  0.160 0.500 0.440 0.930 ;
    END
END CLKAND2X6TR

MACRO CLKAND2X4TR
    CLASS CORE ;
    FOREIGN CLKAND2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.590 2.320 1.360 ;
        RECT  1.760 0.500 2.040 3.160 ;
        END
        ANTENNADIFFAREA 3.758 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.160 1.750 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.680 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.560 -0.280 2.800 0.280 ;
        RECT  1.280 -0.280 1.560 0.760 ;
        RECT  0.000 -0.280 1.280 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 3.320 2.800 3.880 ;
        RECT  2.240 1.910 2.520 3.880 ;
        RECT  1.560 3.320 2.240 3.880 ;
        RECT  1.280 2.230 1.560 3.880 ;
        RECT  0.520 3.320 1.280 3.880 ;
        RECT  0.240 2.620 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.360 1.600 1.640 ;
        RECT  1.320 0.920 1.480 2.070 ;
        RECT  0.680 0.920 1.320 1.080 ;
        RECT  1.000 1.910 1.320 2.070 ;
        RECT  0.720 1.910 1.000 2.660 ;
        RECT  0.400 0.800 0.680 1.080 ;
    END
END CLKAND2X4TR

MACRO CLKAND2X3TR
    CLASS CORE ;
    FOREIGN CLKAND2X3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.900 0.840 1.930 2.070 ;
        RECT  1.810 0.590 1.900 2.070 ;
        RECT  1.770 0.590 1.810 2.820 ;
        RECT  1.600 0.590 1.770 1.310 ;
        RECT  1.650 1.910 1.770 2.820 ;
        RECT  1.530 2.260 1.650 2.820 ;
        END
        ANTENNADIFFAREA 3.222 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.240 1.120 1.560 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.450 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1272 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.280 2.400 0.280 ;
        RECT  1.010 -0.280 1.290 0.760 ;
        RECT  0.000 -0.280 1.010 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 3.320 2.400 3.880 ;
        RECT  2.010 2.260 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.040 2.410 1.330 3.880 ;
        RECT  0.380 3.320 1.040 3.880 ;
        RECT  0.090 2.520 0.380 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.470 1.610 1.750 ;
        RECT  1.280 0.920 1.440 2.070 ;
        RECT  0.450 0.920 1.280 1.080 ;
        RECT  0.850 1.910 1.280 2.070 ;
        RECT  0.570 1.910 0.850 2.690 ;
        RECT  0.170 0.800 0.450 1.080 ;
    END
END CLKAND2X3TR

MACRO CLKAND2X2TR
    CLASS CORE ;
    FOREIGN CLKAND2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.030 1.920 3.160 ;
        RECT  1.600 1.030 1.760 1.310 ;
        RECT  1.600 1.910 1.760 3.160 ;
        END
        ANTENNADIFFAREA 2.848 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.830 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.520 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0912 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.080 -0.280 1.360 0.400 ;
        RECT  0.000 -0.280 1.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 3.320 2.000 3.880 ;
        RECT  1.080 2.590 1.360 3.880 ;
        RECT  0.380 3.320 1.080 3.880 ;
        RECT  0.090 2.140 0.380 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.470 1.600 1.750 ;
        RECT  1.280 0.910 1.440 2.370 ;
        RECT  0.480 0.910 1.280 1.070 ;
        RECT  0.560 2.210 1.280 2.370 ;
        RECT  0.200 0.910 0.480 1.160 ;
    END
END CLKAND2X2TR

MACRO CLKAND2X12TR
    CLASS CORE ;
    FOREIGN CLKAND2X12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 0.490 4.720 3.160 ;
        RECT  4.280 0.490 4.440 1.370 ;
        RECT  3.760 0.560 4.280 1.370 ;
        RECT  3.520 0.560 3.760 3.160 ;
        RECT  3.480 0.440 3.520 3.160 ;
        RECT  3.240 0.440 3.480 0.720 ;
        RECT  2.480 0.560 3.240 0.720 ;
        RECT  2.200 0.440 2.480 0.720 ;
        END
        ANTENNADIFFAREA 9.024 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.700 3.000 1.860 ;
        RECT  0.320 1.240 0.590 1.860 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.4872 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.380 2.520 1.540 ;
        RECT  0.890 0.920 1.130 1.540 ;
        RECT  0.760 0.920 0.890 1.080 ;
        RECT  0.600 0.440 0.760 1.080 ;
        RECT  0.480 0.440 0.600 0.760 ;
        END
        ANTENNAGATEAREA 0.4872 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.040 -0.280 5.600 0.280 ;
        RECT  3.760 -0.280 4.040 0.400 ;
        RECT  3.000 -0.280 3.760 0.280 ;
        RECT  2.720 -0.280 3.000 0.400 ;
        RECT  2.000 -0.280 2.720 0.280 ;
        RECT  1.730 -0.280 2.000 0.670 ;
        RECT  0.320 -0.280 1.730 0.280 ;
        RECT  0.100 -0.280 0.320 0.670 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 3.320 5.600 3.880 ;
        RECT  4.960 1.950 5.240 3.880 ;
        RECT  4.240 3.320 4.960 3.880 ;
        RECT  3.960 1.710 4.240 3.880 ;
        RECT  3.280 3.320 3.960 3.880 ;
        RECT  3.000 2.400 3.280 3.880 ;
        RECT  2.320 3.320 3.000 3.880 ;
        RECT  2.040 2.400 2.320 3.880 ;
        RECT  1.350 3.320 2.040 3.880 ;
        RECT  1.070 2.400 1.350 3.880 ;
        RECT  0.390 3.320 1.070 3.880 ;
        RECT  0.110 2.250 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.160 0.880 3.320 2.240 ;
        RECT  3.040 0.880 3.160 1.160 ;
        RECT  2.800 2.080 3.160 2.240 ;
        RECT  1.570 0.880 3.040 1.040 ;
        RECT  2.520 2.080 2.800 2.950 ;
        RECT  1.840 2.080 2.520 2.240 ;
        RECT  1.560 2.080 1.840 2.950 ;
        RECT  1.410 0.600 1.570 1.040 ;
        RECT  0.870 2.080 1.560 2.240 ;
        RECT  1.200 0.600 1.410 0.760 ;
        RECT  0.920 0.440 1.200 0.760 ;
        RECT  0.590 2.080 0.870 2.950 ;
    END
END CLKAND2X12TR

MACRO BUFX8TR
    CLASS CORE ;
    FOREIGN BUFX8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.840 2.920 2.560 ;
        RECT  2.810 1.840 2.850 3.160 ;
        RECT  2.530 0.590 2.810 3.160 ;
        RECT  2.080 0.840 2.530 2.560 ;
        RECT  1.850 0.840 2.080 1.320 ;
        RECT  1.810 1.920 2.080 2.560 ;
        RECT  1.570 0.610 1.850 1.320 ;
        RECT  1.530 1.920 1.810 3.160 ;
        END
        ANTENNADIFFAREA 7.92 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 1.050 1.650 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.408 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 -0.280 3.600 0.280 ;
        RECT  3.010 -0.280 3.290 1.240 ;
        RECT  2.330 -0.280 3.010 0.280 ;
        RECT  2.050 -0.280 2.330 0.680 ;
        RECT  1.370 -0.280 2.050 0.280 ;
        RECT  1.090 -0.280 1.370 0.760 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 3.320 3.600 3.880 ;
        RECT  3.110 1.920 3.330 3.880 ;
        RECT  2.330 3.320 3.110 3.880 ;
        RECT  2.050 2.780 2.330 3.880 ;
        RECT  1.330 3.320 2.050 3.880 ;
        RECT  1.050 2.270 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.560 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.370 1.480 1.920 1.760 ;
        RECT  1.210 0.920 1.370 2.080 ;
        RECT  0.850 0.920 1.210 1.080 ;
        RECT  0.850 1.920 1.210 2.080 ;
        RECT  0.570 0.650 0.850 1.080 ;
        RECT  0.570 1.920 0.850 2.950 ;
    END
END BUFX8TR

MACRO BUFX6TR
    CLASS CORE ;
    FOREIGN BUFX6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.830 0.440 3.100 3.160 ;
        RECT  2.820 0.950 2.830 3.160 ;
        RECT  2.710 0.950 2.820 2.570 ;
        RECT  2.070 0.950 2.710 1.310 ;
        RECT  2.060 1.840 2.710 2.570 ;
        RECT  1.790 0.550 2.070 1.310 ;
        RECT  1.780 1.840 2.060 3.160 ;
        END
        ANTENNADIFFAREA 7.466 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 1.270 1.640 ;
        END
        ANTENNAGATEAREA 0.3168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.280 3.200 0.280 ;
        RECT  2.310 -0.280 2.590 0.730 ;
        RECT  1.590 -0.280 2.310 0.280 ;
        RECT  1.310 -0.280 1.590 0.760 ;
        RECT  0.590 -0.280 1.310 0.280 ;
        RECT  0.310 -0.280 0.590 1.040 ;
        RECT  0.000 -0.280 0.310 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 3.320 3.200 3.880 ;
        RECT  2.300 2.860 2.580 3.880 ;
        RECT  1.580 3.320 2.300 3.880 ;
        RECT  1.260 2.400 1.580 3.880 ;
        RECT  0.620 3.320 1.260 3.880 ;
        RECT  0.340 1.910 0.620 3.880 ;
        RECT  0.000 3.320 0.340 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.590 1.470 2.260 1.680 ;
        RECT  1.430 0.920 1.590 2.070 ;
        RECT  1.070 0.920 1.430 1.080 ;
        RECT  1.100 1.910 1.430 2.070 ;
        RECT  0.880 1.910 1.100 2.680 ;
        RECT  0.790 0.800 1.070 1.080 ;
    END
END BUFX6TR

MACRO BUFX4TR
    CLASS CORE ;
    FOREIGN BUFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.010 1.920 2.200 ;
        RECT  1.520 1.010 1.680 1.310 ;
        RECT  1.520 1.930 1.680 2.200 ;
        RECT  1.240 0.450 1.520 1.310 ;
        RECT  1.240 1.930 1.520 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.760 1.660 ;
        RECT  0.440 1.380 0.480 1.660 ;
        END
        ANTENNAGATEAREA 0.204 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.040 -0.280 2.400 0.280 ;
        RECT  1.760 -0.280 2.040 0.840 ;
        RECT  1.000 -0.280 1.760 0.280 ;
        RECT  0.720 -0.280 1.000 0.800 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.040 3.320 2.400 3.880 ;
        RECT  1.760 2.460 2.040 3.880 ;
        RECT  1.040 3.320 1.760 3.880 ;
        RECT  0.760 2.140 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 1.490 1.290 1.770 ;
        RECT  0.920 1.490 1.080 1.980 ;
        RECT  0.560 1.820 0.920 1.980 ;
        RECT  0.280 1.820 0.560 2.950 ;
        RECT  0.260 0.650 0.320 1.260 ;
        RECT  0.260 1.820 0.280 1.980 ;
        RECT  0.100 0.650 0.260 1.980 ;
    END
END BUFX4TR

MACRO BUFX3TR
    CLASS CORE ;
    FOREIGN BUFX3TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.240 1.920 2.360 ;
        RECT  1.640 1.040 1.800 2.360 ;
        RECT  1.440 1.040 1.640 1.200 ;
        RECT  1.430 2.160 1.640 2.360 ;
        RECT  1.160 0.920 1.440 1.200 ;
        RECT  1.130 2.160 1.430 2.870 ;
        END
        ANTENNADIFFAREA 2.97 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.1608 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.280 2.000 0.280 ;
        RECT  1.630 -0.280 1.910 0.870 ;
        RECT  0.930 -0.280 1.630 0.280 ;
        RECT  0.610 -0.280 0.930 1.030 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.600 2.580 1.910 3.880 ;
        RECT  0.910 3.320 1.600 3.880 ;
        RECT  0.610 2.350 0.910 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.270 1.360 1.390 1.680 ;
        RECT  1.100 1.360 1.270 1.960 ;
        RECT  0.380 1.800 1.100 1.960 ;
        RECT  0.260 0.800 0.410 1.080 ;
        RECT  0.260 1.800 0.380 2.690 ;
        RECT  0.100 0.800 0.260 2.690 ;
    END
END BUFX3TR

MACRO BUFX2TR
    CLASS CORE ;
    FOREIGN BUFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 0.840 1.620 1.160 ;
        RECT  1.300 0.840 1.460 2.420 ;
        RECT  1.040 0.840 1.300 1.250 ;
        RECT  1.120 2.120 1.300 2.420 ;
        END
        ANTENNADIFFAREA 2.1 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 0.840 0.820 1.160 ;
        RECT  0.480 0.840 0.680 1.640 ;
        RECT  0.460 1.420 0.480 1.640 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.280 2.000 0.280 ;
        RECT  1.550 -0.280 1.840 0.680 ;
        RECT  0.800 -0.280 1.550 0.280 ;
        RECT  0.520 -0.280 0.800 0.600 ;
        RECT  0.000 -0.280 0.520 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 3.320 2.000 3.880 ;
        RECT  1.630 2.060 1.870 3.880 ;
        RECT  0.890 3.320 1.630 3.880 ;
        RECT  0.600 2.160 0.890 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 1.510 1.120 1.790 ;
        RECT  0.840 1.510 1.000 1.960 ;
        RECT  0.400 1.800 0.840 1.960 ;
        RECT  0.300 1.800 0.400 2.280 ;
        RECT  0.300 1.000 0.320 1.290 ;
        RECT  0.140 1.000 0.300 2.280 ;
    END
END BUFX2TR

MACRO BUFX20TR
    CLASS CORE ;
    FOREIGN BUFX20TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.610 0.840 6.760 2.070 ;
        RECT  6.330 0.840 6.610 2.770 ;
        RECT  5.650 0.840 6.330 2.070 ;
        RECT  5.370 0.440 5.650 3.160 ;
        RECT  4.690 1.110 5.370 2.070 ;
        RECT  4.410 0.440 4.690 3.160 ;
        RECT  3.730 1.110 4.410 2.070 ;
        RECT  3.450 0.440 3.730 3.160 ;
        RECT  2.770 1.110 3.450 2.070 ;
        RECT  2.520 0.440 2.770 3.160 ;
        RECT  2.490 0.440 2.520 1.370 ;
        RECT  2.490 1.870 2.520 3.160 ;
        END
        ANTENNADIFFAREA 19.696 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 1.530 1.640 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 1.056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.210 -0.280 7.600 0.280 ;
        RECT  6.920 -0.280 7.210 1.310 ;
        RECT  6.130 -0.280 6.920 0.340 ;
        RECT  5.850 -0.280 6.130 0.670 ;
        RECT  5.170 -0.280 5.850 0.280 ;
        RECT  4.890 -0.280 5.170 0.760 ;
        RECT  4.210 -0.280 4.890 0.280 ;
        RECT  3.930 -0.280 4.210 0.800 ;
        RECT  3.250 -0.280 3.930 0.280 ;
        RECT  2.960 -0.280 3.250 0.810 ;
        RECT  2.290 -0.280 2.960 0.280 ;
        RECT  2.010 -0.280 2.290 1.190 ;
        RECT  1.330 -0.280 2.010 0.280 ;
        RECT  1.050 -0.280 1.330 0.760 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.090 3.320 7.600 3.880 ;
        RECT  6.810 2.270 7.090 3.880 ;
        RECT  6.130 3.260 6.810 3.880 ;
        RECT  5.850 2.480 6.130 3.880 ;
        RECT  5.170 3.320 5.850 3.880 ;
        RECT  4.890 2.400 5.170 3.880 ;
        RECT  4.210 3.320 4.890 3.880 ;
        RECT  3.930 2.390 4.210 3.880 ;
        RECT  3.250 3.320 3.930 3.880 ;
        RECT  2.970 2.390 3.250 3.880 ;
        RECT  2.290 3.320 2.970 3.880 ;
        RECT  2.010 1.910 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.120 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.270 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.850 1.470 2.350 1.750 ;
        RECT  1.810 0.920 1.850 3.120 ;
        RECT  1.690 0.440 1.810 3.120 ;
        RECT  1.530 0.440 1.690 1.080 ;
        RECT  1.530 1.800 1.690 3.120 ;
        RECT  0.850 0.920 1.530 1.080 ;
        RECT  0.850 1.800 1.530 1.960 ;
        RECT  0.570 0.440 0.850 1.080 ;
        RECT  0.570 1.800 0.850 3.130 ;
    END
END BUFX20TR

MACRO BUFX16TR
    CLASS CORE ;
    FOREIGN BUFX16TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.170 0.840 5.670 2.080 ;
        RECT  4.890 0.840 5.170 2.810 ;
        RECT  4.370 0.840 4.890 2.080 ;
        RECT  4.210 0.500 4.370 2.080 ;
        RECT  4.090 0.500 4.210 3.160 ;
        RECT  3.930 1.100 4.090 3.160 ;
        RECT  3.330 1.100 3.930 2.070 ;
        RECT  3.250 0.500 3.330 2.070 ;
        RECT  3.050 0.500 3.250 3.160 ;
        RECT  2.970 1.100 3.050 3.160 ;
        RECT  2.290 1.100 2.970 2.070 ;
        RECT  2.090 0.500 2.290 3.160 ;
        RECT  2.010 0.500 2.090 1.280 ;
        RECT  2.010 1.980 2.090 3.160 ;
        END
        ANTENNADIFFAREA 15.032 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.240 1.530 1.640 ;
        END
        ANTENNAGATEAREA 0.7992 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 -0.280 6.000 0.280 ;
        RECT  5.530 -0.280 5.810 0.610 ;
        RECT  4.610 -0.280 5.530 0.340 ;
        RECT  3.850 -0.280 4.610 0.280 ;
        RECT  3.570 -0.280 3.850 0.800 ;
        RECT  2.810 -0.280 3.570 0.280 ;
        RECT  2.530 -0.280 2.810 0.790 ;
        RECT  1.810 -0.280 2.530 0.280 ;
        RECT  1.530 -0.280 1.810 0.670 ;
        RECT  0.850 -0.280 1.530 0.280 ;
        RECT  0.570 -0.280 0.850 0.670 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 3.320 6.000 3.880 ;
        RECT  5.410 2.400 5.690 3.880 ;
        RECT  4.690 3.260 5.410 3.880 ;
        RECT  4.410 2.330 4.690 3.880 ;
        RECT  3.730 3.320 4.410 3.880 ;
        RECT  3.450 2.490 3.730 3.880 ;
        RECT  2.770 3.320 3.450 3.880 ;
        RECT  2.490 2.390 2.770 3.880 ;
        RECT  1.810 3.320 2.490 3.880 ;
        RECT  1.530 2.120 1.810 3.880 ;
        RECT  0.850 3.320 1.530 3.880 ;
        RECT  0.570 2.120 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.850 1.470 1.930 1.750 ;
        RECT  1.690 0.920 1.850 1.960 ;
        RECT  1.330 0.920 1.690 1.080 ;
        RECT  1.330 1.800 1.690 1.960 ;
        RECT  1.050 0.540 1.330 1.080 ;
        RECT  1.050 1.800 1.330 3.160 ;
        RECT  0.370 0.920 1.050 1.080 ;
        RECT  0.370 1.800 1.050 1.960 ;
        RECT  0.090 0.540 0.370 1.080 ;
        RECT  0.090 1.800 0.370 3.160 ;
    END
END BUFX16TR

MACRO BUFX12TR
    CLASS CORE ;
    FOREIGN BUFX12TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.720 1.260 3.850 2.760 ;
        RECT  3.450 1.040 3.720 2.760 ;
        RECT  3.080 1.040 3.450 1.980 ;
        RECT  2.770 1.260 3.080 1.980 ;
        RECT  2.490 0.440 2.770 3.160 ;
        RECT  1.810 1.260 2.490 1.980 ;
        RECT  1.550 0.440 1.810 3.160 ;
        RECT  1.530 0.440 1.550 0.730 ;
        RECT  1.530 2.180 1.550 3.160 ;
        END
        ANTENNADIFFAREA 10.872 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 1.050 1.610 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 -0.280 4.400 0.280 ;
        RECT  4.080 -0.280 4.240 1.110 ;
        RECT  3.250 -0.280 4.080 0.280 ;
        RECT  2.970 -0.280 3.250 0.620 ;
        RECT  2.290 -0.280 2.970 0.280 ;
        RECT  2.010 -0.280 2.290 1.100 ;
        RECT  1.330 -0.280 2.010 0.280 ;
        RECT  1.050 -0.280 1.330 0.760 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 3.320 4.400 3.880 ;
        RECT  4.010 1.930 4.170 3.880 ;
        RECT  3.250 3.320 4.010 3.880 ;
        RECT  2.970 2.250 3.250 3.880 ;
        RECT  2.290 3.320 2.970 3.880 ;
        RECT  2.010 2.380 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.090 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.230 0.920 1.390 1.930 ;
        RECT  0.850 0.920 1.230 1.080 ;
        RECT  0.850 1.770 1.230 1.930 ;
        RECT  0.570 0.440 0.850 1.080 ;
        RECT  0.570 1.770 0.850 3.160 ;
    END
END BUFX12TR

MACRO AOI33XLTR
    CLASS CORE ;
    FOREIGN AOI33XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 2.160 3.400 2.600 ;
        RECT  2.440 2.160 3.120 2.320 ;
        RECT  2.360 0.840 2.720 1.160 ;
        RECT  2.360 2.160 2.440 2.600 ;
        RECT  2.200 0.840 2.360 2.600 ;
        RECT  1.850 0.840 2.200 1.080 ;
        RECT  2.160 2.320 2.200 2.600 ;
        RECT  1.560 0.800 1.850 1.080 ;
        END
        ANTENNADIFFAREA 2.936 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.640 1.610 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.120 2.000 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.410 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.840 3.520 1.960 ;
        RECT  3.090 1.220 3.280 1.480 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.640 3.120 1.960 ;
        RECT  2.520 1.680 2.880 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 2.040 1.610 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.200 -0.280 3.600 0.280 ;
        RECT  2.920 -0.280 3.200 0.680 ;
        RECT  0.600 -0.280 2.920 0.280 ;
        RECT  0.320 -0.280 0.600 1.080 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 3.600 3.880 ;
        RECT  1.120 2.480 1.400 3.880 ;
        RECT  0.440 3.260 1.120 3.880 ;
        RECT  0.160 2.540 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.640 2.480 2.920 2.920 ;
        RECT  1.880 2.760 2.640 2.920 ;
        RECT  1.720 2.160 1.880 2.920 ;
        RECT  1.600 2.160 1.720 2.600 ;
        RECT  0.920 2.160 1.600 2.320 ;
        RECT  0.640 2.160 0.920 2.600 ;
    END
END AOI33XLTR

MACRO AOI33X4TR
    CLASS CORE ;
    FOREIGN AOI33X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.920 1.040 5.120 2.010 ;
        RECT  4.900 0.440 4.920 2.010 ;
        RECT  4.880 0.440 4.900 3.160 ;
        RECT  4.640 0.440 4.880 1.310 ;
        RECT  4.660 1.790 4.880 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.240 0.660 1.560 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.180 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.840 1.520 1.520 ;
        RECT  1.280 0.840 1.360 1.160 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.490 3.120 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.580 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.580 1.990 1.960 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.400 -0.280 5.600 0.280 ;
        RECT  5.110 -0.280 5.400 0.670 ;
        RECT  4.380 -0.280 5.110 0.280 ;
        RECT  4.220 -0.280 4.380 1.310 ;
        RECT  3.100 -0.280 4.220 0.280 ;
        RECT  2.820 -0.280 3.100 1.010 ;
        RECT  0.680 -0.280 2.820 0.280 ;
        RECT  0.360 -0.280 0.680 1.010 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.390 3.320 5.600 3.880 ;
        RECT  5.120 2.170 5.390 3.880 ;
        RECT  4.380 3.320 5.120 3.880 ;
        RECT  4.220 1.910 4.380 3.880 ;
        RECT  1.420 3.320 4.220 3.880 ;
        RECT  1.130 2.520 1.420 3.880 ;
        RECT  0.460 3.320 1.130 3.880 ;
        RECT  0.160 2.520 0.460 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.060 1.470 4.640 1.630 ;
        RECT  3.940 1.090 4.060 2.360 ;
        RECT  3.900 1.090 3.940 2.950 ;
        RECT  3.740 0.870 3.900 1.250 ;
        RECT  3.680 1.980 3.900 2.950 ;
        RECT  3.440 1.420 3.740 1.580 ;
        RECT  3.280 1.170 3.440 2.290 ;
        RECT  2.310 1.170 3.280 1.330 ;
        RECT  1.910 2.520 2.980 2.680 ;
        RECT  2.310 2.180 2.490 2.340 ;
        RECT  2.150 1.170 2.310 2.340 ;
        RECT  1.980 1.170 2.150 1.330 ;
        RECT  1.680 0.800 1.980 1.330 ;
        RECT  1.750 2.170 1.910 2.680 ;
        RECT  0.870 2.170 1.750 2.330 ;
        RECT  0.710 2.170 0.870 2.750 ;
    END
END AOI33X4TR

MACRO AOI33X2TR
    CLASS CORE ;
    FOREIGN AOI33X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.070 6.200 2.200 ;
        RECT  5.920 1.070 6.040 1.230 ;
        RECT  5.680 2.040 6.040 2.200 ;
        RECT  5.640 0.500 5.920 1.230 ;
        RECT  5.400 2.040 5.680 2.780 ;
        RECT  3.200 0.560 5.640 0.720 ;
        RECT  5.160 2.040 5.400 2.200 ;
        RECT  4.840 2.040 5.160 2.360 ;
        RECT  4.720 2.120 4.840 2.360 ;
        RECT  4.440 2.120 4.720 2.780 ;
        RECT  3.760 2.120 4.440 2.280 ;
        RECT  3.480 2.120 3.760 2.780 ;
        RECT  2.920 0.560 3.200 1.080 ;
        RECT  0.640 0.920 2.920 1.080 ;
        RECT  0.360 0.790 0.640 1.120 ;
        END
        ANTENNADIFFAREA 9 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 2.040 1.580 ;
        RECT  1.360 1.300 1.640 1.580 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.640 2.520 1.920 ;
        RECT  1.160 1.760 2.240 1.920 ;
        RECT  0.880 1.240 1.160 1.920 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.830 3.000 2.110 ;
        RECT  2.720 1.830 2.880 2.240 ;
        RECT  0.720 2.080 2.720 2.240 ;
        RECT  0.560 1.640 0.720 2.240 ;
        RECT  0.400 1.640 0.560 1.960 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.240 4.920 1.560 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.720 5.400 1.880 ;
        RECT  3.680 1.640 3.960 1.960 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.600 1.390 5.880 1.670 ;
        RECT  5.240 1.390 5.600 1.550 ;
        RECT  5.080 0.920 5.240 1.550 ;
        RECT  3.520 0.920 5.080 1.080 ;
        RECT  3.360 0.920 3.520 1.560 ;
        RECT  3.200 1.240 3.360 1.560 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 -0.280 6.400 0.280 ;
        RECT  4.400 -0.280 4.680 0.400 ;
        RECT  1.950 -0.280 4.400 0.280 ;
        RECT  1.660 -0.280 1.950 0.760 ;
        RECT  0.000 -0.280 1.660 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.800 3.320 6.400 3.880 ;
        RECT  2.520 2.720 2.800 3.880 ;
        RECT  1.840 3.320 2.520 3.880 ;
        RECT  1.560 2.720 1.840 3.880 ;
        RECT  0.880 3.320 1.560 3.880 ;
        RECT  0.600 2.720 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.040 2.550 6.160 2.830 ;
        RECT  5.880 2.550 6.040 3.100 ;
        RECT  5.200 2.940 5.880 3.100 ;
        RECT  4.920 2.550 5.200 3.100 ;
        RECT  4.240 2.940 4.920 3.100 ;
        RECT  3.960 2.550 4.240 3.100 ;
        RECT  3.280 2.940 3.960 3.100 ;
        RECT  3.120 2.400 3.280 3.100 ;
        RECT  3.000 2.400 3.120 2.680 ;
        RECT  2.320 2.400 3.000 2.560 ;
        RECT  2.040 2.400 2.320 3.000 ;
        RECT  1.360 2.400 2.040 2.560 ;
        RECT  1.080 2.400 1.360 3.000 ;
        RECT  0.400 2.400 1.080 2.560 ;
        RECT  0.120 2.400 0.400 3.000 ;
    END
END AOI33X2TR

MACRO AOI33X1TR
    CLASS CORE ;
    FOREIGN AOI33X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 2.160 3.480 2.890 ;
        RECT  2.440 2.160 3.200 2.320 ;
        RECT  2.440 1.240 2.720 1.560 ;
        RECT  2.280 1.080 2.440 2.440 ;
        RECT  1.960 1.080 2.280 1.240 ;
        RECT  2.160 2.120 2.280 2.440 ;
        RECT  1.680 0.650 1.960 1.240 ;
        END
        ANTENNADIFFAREA 5.352 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.400 0.640 1.680 ;
        RECT  0.320 1.400 0.360 2.360 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.480 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.200 1.520 1.680 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.440 3.520 1.560 ;
        RECT  3.010 1.200 3.280 1.480 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.640 3.120 2.000 ;
        RECT  2.600 1.720 2.880 2.000 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.500 2.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 -0.280 3.600 0.280 ;
        RECT  2.840 -0.280 3.120 0.800 ;
        RECT  0.600 -0.280 2.840 0.340 ;
        RECT  0.320 -0.280 0.600 0.970 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 3.600 3.880 ;
        RECT  1.120 2.610 1.400 3.880 ;
        RECT  0.440 3.320 1.120 3.880 ;
        RECT  0.160 2.610 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.720 2.610 3.000 2.890 ;
        RECT  1.880 2.730 2.720 2.890 ;
        RECT  1.600 2.160 1.880 2.890 ;
        RECT  0.920 2.160 1.600 2.320 ;
        RECT  0.640 2.160 0.920 2.890 ;
    END
END AOI33X1TR

MACRO AOI32XLTR
    CLASS CORE ;
    FOREIGN AOI32XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.840 2.320 1.160 ;
        RECT  2.110 0.840 2.270 2.540 ;
        RECT  2.080 0.840 2.110 1.160 ;
        RECT  1.950 2.380 2.110 2.540 ;
        RECT  1.350 1.000 2.080 1.160 ;
        END
        ANTENNADIFFAREA 1.72 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        RECT  2.430 1.720 2.480 2.360 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.600 1.950 1.980 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.410 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.720 0.970 2.360 ;
        RECT  0.480 2.040 0.810 2.360 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.400 1.430 1.680 ;
        RECT  1.150 1.240 1.190 1.680 ;
        RECT  0.880 1.240 1.150 1.560 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.280 2.800 0.280 ;
        RECT  2.230 -0.280 2.510 0.680 ;
        RECT  0.470 -0.280 2.230 0.340 ;
        RECT  0.190 -0.280 0.470 1.230 ;
        RECT  0.000 -0.280 0.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 3.320 2.800 3.880 ;
        RECT  0.180 3.260 1.230 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.430 2.520 2.710 2.860 ;
        RECT  1.710 2.700 2.430 2.860 ;
        RECT  1.520 2.520 1.710 2.860 ;
        RECT  0.540 2.520 1.520 2.680 ;
    END
END AOI32XLTR

MACRO AOI32X4TR
    CLASS CORE ;
    FOREIGN AOI32X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.040 4.320 2.030 ;
        RECT  4.100 1.040 4.240 3.160 ;
        RECT  4.080 0.440 4.100 3.160 ;
        RECT  3.840 0.440 4.080 1.310 ;
        RECT  4.000 1.790 4.080 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.840 2.720 1.430 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.130 1.950 1.560 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.180 0.650 1.560 ;
        RECT  0.080 1.180 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.540 1.130 1.830 ;
        RECT  0.880 1.540 1.120 2.010 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.240 1.520 2.360 ;
        RECT  1.280 2.040 1.360 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.280 4.800 0.280 ;
        RECT  4.290 -0.280 4.570 0.750 ;
        RECT  3.610 -0.280 4.290 0.280 ;
        RECT  3.330 -0.280 3.610 1.070 ;
        RECT  2.650 -0.280 3.330 0.280 ;
        RECT  2.370 -0.280 2.650 0.340 ;
        RECT  0.670 -0.280 2.370 0.280 ;
        RECT  0.380 -0.280 0.670 0.980 ;
        RECT  0.000 -0.280 0.380 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 3.320 4.800 3.880 ;
        RECT  4.480 2.430 4.700 3.880 ;
        RECT  3.670 3.320 4.480 3.880 ;
        RECT  2.020 3.260 3.670 3.880 ;
        RECT  1.510 3.320 2.020 3.880 ;
        RECT  1.230 2.840 1.510 3.880 ;
        RECT  0.500 3.320 1.230 3.880 ;
        RECT  0.230 2.540 0.500 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.670 1.470 3.890 1.630 ;
        RECT  3.510 1.230 3.670 2.750 ;
        RECT  3.130 1.230 3.510 1.390 ;
        RECT  2.710 2.590 3.510 2.750 ;
        RECT  3.100 1.590 3.260 1.930 ;
        RECT  2.970 0.520 3.130 1.390 ;
        RECT  2.390 1.770 3.100 1.930 ;
        RECT  2.850 0.520 2.970 0.680 ;
        RECT  2.590 2.120 2.870 2.340 ;
        RECT  1.850 2.180 2.590 2.340 ;
        RECT  2.270 1.770 2.390 2.020 ;
        RECT  2.110 0.810 2.270 2.020 ;
        RECT  1.530 0.810 2.110 0.970 ;
        RECT  1.690 2.060 1.850 2.680 ;
        RECT  0.940 2.520 1.690 2.680 ;
        RECT  0.770 2.300 0.940 2.680 ;
    END
END AOI32X4TR

MACRO AOI32X2TR
    CLASS CORE ;
    FOREIGN AOI32X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 0.710 4.630 2.890 ;
        RECT  4.400 0.710 4.440 1.080 ;
        RECT  4.260 2.040 4.440 2.890 ;
        RECT  2.950 0.920 4.400 1.080 ;
        RECT  3.610 2.040 4.260 2.360 ;
        RECT  3.340 2.040 3.610 2.840 ;
        RECT  2.790 0.440 2.950 1.080 ;
        RECT  0.190 0.920 2.790 1.080 ;
        END
        ANTENNADIFFAREA 6.964 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.240 3.960 1.560 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.120 1.380 4.280 1.880 ;
        RECT  3.250 1.720 4.120 1.880 ;
        RECT  3.080 1.240 3.250 1.880 ;
        RECT  2.880 1.240 3.080 1.560 ;
        END
        ANTENNAGATEAREA 0.3264 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.730 1.600 ;
        END
        ANTENNAGATEAREA 0.3696 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.610 2.350 1.960 ;
        RECT  1.120 1.800 2.190 1.960 ;
        RECT  0.850 1.640 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.3696 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.760 2.900 1.920 ;
        RECT  2.590 1.760 2.750 2.280 ;
        RECT  0.370 2.120 2.590 2.280 ;
        RECT  0.370 1.580 0.650 1.860 ;
        RECT  0.360 1.580 0.370 2.280 ;
        RECT  0.330 1.240 0.360 2.280 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.3696 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.850 -0.280 4.800 0.280 ;
        RECT  3.570 -0.280 3.850 0.760 ;
        RECT  1.850 -0.280 3.570 0.280 ;
        RECT  1.570 -0.280 1.850 0.760 ;
        RECT  0.000 -0.280 1.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 3.320 4.800 3.880 ;
        RECT  2.330 3.260 2.610 3.880 ;
        RECT  1.810 3.320 2.330 3.880 ;
        RECT  1.530 3.260 1.810 3.880 ;
        RECT  0.770 3.320 1.530 3.880 ;
        RECT  0.490 3.260 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 2.620 4.090 3.160 ;
        RECT  3.070 3.000 3.810 3.160 ;
        RECT  2.910 2.080 3.070 3.160 ;
        RECT  0.990 2.440 2.910 2.720 ;
        RECT  0.090 2.520 0.990 2.720 ;
    END
END AOI32X2TR

MACRO AOI32X1TR
    CLASS CORE ;
    FOREIGN AOI32X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.840 2.320 1.160 ;
        RECT  2.110 0.840 2.270 2.620 ;
        RECT  1.350 0.840 2.110 1.160 ;
        RECT  1.950 2.290 2.110 2.620 ;
        END
        ANTENNADIFFAREA 2.904 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        RECT  2.430 1.720 2.480 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.600 1.950 1.980 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.410 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.720 0.970 2.360 ;
        RECT  0.480 2.040 0.810 2.360 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.400 1.430 1.680 ;
        RECT  1.150 1.240 1.190 1.680 ;
        RECT  0.880 1.240 1.150 1.560 ;
        END
        ANTENNAGATEAREA 0.1872 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.280 2.800 0.280 ;
        RECT  2.230 -0.280 2.510 0.680 ;
        RECT  0.470 -0.280 2.230 0.340 ;
        RECT  0.190 -0.280 0.470 1.230 ;
        RECT  0.000 -0.280 0.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 3.320 2.800 3.880 ;
        RECT  0.180 3.260 1.230 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.430 2.590 2.710 2.950 ;
        RECT  1.750 2.790 2.430 2.950 ;
        RECT  1.470 2.160 1.750 2.950 ;
        RECT  0.850 2.780 1.470 2.950 ;
        RECT  0.540 2.610 0.850 2.950 ;
    END
END AOI32X1TR

MACRO AOI31XLTR
    CLASS CORE ;
    FOREIGN AOI31XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.230 2.320 2.630 ;
        RECT  2.080 0.920 2.240 2.630 ;
        RECT  1.660 0.920 2.080 1.080 ;
        RECT  2.010 2.330 2.080 2.630 ;
        RECT  1.380 0.800 1.660 1.080 ;
        END
        ANTENNADIFFAREA 1.568 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.700 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.200 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.580 1.050 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.240 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1104 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  1.940 -0.280 2.220 0.760 ;
        RECT  0.530 -0.280 1.940 0.340 ;
        RECT  0.250 -0.280 0.530 0.930 ;
        RECT  0.000 -0.280 0.250 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 3.320 2.400 3.880 ;
        RECT  1.050 2.530 1.330 3.880 ;
        RECT  0.370 3.260 1.050 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 2.210 1.810 2.600 ;
        RECT  0.850 2.210 1.530 2.370 ;
        RECT  0.570 2.210 0.850 2.630 ;
    END
END AOI31XLTR

MACRO AOI31X4TR
    CLASS CORE ;
    FOREIGN AOI31X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.040 3.920 1.940 ;
        RECT  3.700 1.040 3.830 3.160 ;
        RECT  3.610 0.440 3.700 3.160 ;
        RECT  3.420 0.440 3.610 1.310 ;
        RECT  3.550 1.910 3.610 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.190 2.080 1.570 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.280 0.660 1.570 ;
        RECT  0.320 1.190 0.360 1.570 ;
        RECT  0.080 1.190 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.600 1.200 1.880 ;
        RECT  0.920 1.600 1.120 2.000 ;
        RECT  0.880 1.640 0.920 2.000 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.260 1.520 2.360 ;
        RECT  1.280 2.040 1.360 2.360 ;
        END
        ANTENNAGATEAREA 0.12 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.180 -0.280 4.400 0.280 ;
        RECT  3.900 -0.280 4.180 0.840 ;
        RECT  3.180 -0.280 3.900 0.280 ;
        RECT  2.900 -0.280 3.180 0.400 ;
        RECT  2.320 -0.280 2.900 0.280 ;
        RECT  2.040 -0.280 2.320 0.400 ;
        RECT  0.660 -0.280 2.040 0.340 ;
        RECT  0.380 -0.280 0.660 1.030 ;
        RECT  0.000 -0.280 0.380 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.300 3.320 4.400 3.880 ;
        RECT  4.020 2.170 4.300 3.880 ;
        RECT  3.250 3.320 4.020 3.880 ;
        RECT  1.710 3.200 3.250 3.880 ;
        RECT  1.400 3.320 1.710 3.880 ;
        RECT  1.140 2.840 1.400 3.880 ;
        RECT  0.490 3.260 1.140 3.880 ;
        RECT  0.180 2.520 0.490 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.960 1.470 3.450 1.750 ;
        RECT  2.800 0.980 2.960 2.750 ;
        RECT  2.560 0.980 2.800 1.260 ;
        RECT  2.730 2.590 2.800 2.750 ;
        RECT  2.450 2.590 2.730 2.870 ;
        RECT  2.440 1.530 2.640 1.810 ;
        RECT  2.400 1.530 2.440 2.400 ;
        RECT  2.240 0.870 2.400 2.400 ;
        RECT  1.780 0.870 2.240 1.030 ;
        RECT  2.160 2.120 2.240 2.400 ;
        RECT  1.840 2.120 1.960 2.400 ;
        RECT  1.680 2.120 1.840 2.680 ;
        RECT  1.500 0.750 1.780 1.030 ;
        RECT  1.000 2.520 1.680 2.680 ;
        RECT  0.840 2.190 1.000 2.680 ;
        RECT  0.720 2.190 0.840 2.470 ;
    END
END AOI31X4TR

MACRO AOI31X2TR
    CLASS CORE ;
    FOREIGN AOI31X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.150 3.920 2.320 ;
        RECT  2.950 1.150 3.680 1.310 ;
        RECT  3.670 2.160 3.680 2.320 ;
        RECT  3.510 2.160 3.670 2.840 ;
        RECT  2.790 0.580 2.950 1.310 ;
        RECT  0.590 0.920 2.790 1.080 ;
        RECT  0.430 0.740 0.590 1.080 ;
        END
        ANTENNADIFFAREA 4.24 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.470 3.520 1.960 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.360 1.580 ;
        RECT  1.720 1.360 2.080 1.580 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.760 2.490 1.920 ;
        RECT  1.280 1.240 1.520 1.920 ;
        RECT  0.890 1.760 1.280 1.920 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.770 2.910 2.050 ;
        RECT  2.710 1.770 2.870 2.240 ;
        RECT  0.670 2.080 2.710 2.240 ;
        RECT  0.670 1.240 0.720 1.560 ;
        RECT  0.510 1.240 0.670 2.240 ;
        RECT  0.470 1.240 0.510 1.700 ;
        END
        ANTENNAGATEAREA 0.3744 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.540 -0.280 4.400 0.280 ;
        RECT  3.250 -0.280 3.540 0.990 ;
        RECT  1.810 -0.280 3.250 0.280 ;
        RECT  1.530 -0.280 1.810 0.760 ;
        RECT  0.000 -0.280 1.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.770 3.320 4.400 3.880 ;
        RECT  2.490 2.720 2.770 3.880 ;
        RECT  1.770 3.320 2.490 3.880 ;
        RECT  1.490 3.260 1.770 3.880 ;
        RECT  0.890 3.320 1.490 3.880 ;
        RECT  0.610 2.720 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.990 2.610 4.150 3.160 ;
        RECT  3.190 3.000 3.990 3.160 ;
        RECT  3.030 2.210 3.190 3.160 ;
        RECT  2.230 2.400 3.030 2.560 ;
        RECT  2.070 2.400 2.230 2.680 ;
        RECT  1.310 2.400 2.070 2.560 ;
        RECT  1.150 2.400 1.310 2.680 ;
        RECT  0.350 2.400 1.150 2.560 ;
        RECT  0.190 2.100 0.350 2.940 ;
    END
END AOI31X2TR

MACRO AOI31X1TR
    CLASS CORE ;
    FOREIGN AOI31X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.640 2.320 2.760 ;
        RECT  2.080 0.920 2.240 2.760 ;
        RECT  1.660 0.920 2.080 1.080 ;
        RECT  2.010 2.080 2.080 2.760 ;
        RECT  1.380 0.800 1.660 1.080 ;
        END
        ANTENNADIFFAREA 2.584 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.700 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.200 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.580 1.050 1.960 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.440 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.18 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  1.940 -0.280 2.220 0.760 ;
        RECT  0.530 -0.280 1.940 0.340 ;
        RECT  0.250 -0.280 0.530 0.930 ;
        RECT  0.000 -0.280 0.250 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 3.320 2.400 3.880 ;
        RECT  1.050 2.440 1.330 3.880 ;
        RECT  0.370 3.260 1.050 3.880 ;
        RECT  0.090 2.560 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 2.120 1.810 2.820 ;
        RECT  0.850 2.120 1.530 2.280 ;
        RECT  0.570 2.120 0.850 2.800 ;
    END
END AOI31X1TR

MACRO AOI2BB2XLTR
    CLASS CORE ;
    FOREIGN AOI2BB2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.080 2.720 2.360 ;
        RECT  2.090 1.080 2.480 1.240 ;
        RECT  2.440 2.040 2.480 2.360 ;
        RECT  2.270 2.040 2.440 2.330 ;
        RECT  1.810 0.900 2.090 1.240 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 2.840 1.160 3.160 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 2.040 1.960 2.360 ;
        RECT  1.640 1.720 1.810 2.360 ;
        RECT  1.530 1.720 1.640 2.000 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.890 1.620 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.650 -0.280 2.800 0.280 ;
        RECT  2.370 -0.280 2.650 0.910 ;
        RECT  1.250 -0.280 2.370 0.280 ;
        RECT  0.970 -0.280 1.250 0.580 ;
        RECT  0.360 -0.280 0.970 0.280 ;
        RECT  0.090 -0.280 0.360 0.580 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.690 3.320 2.800 3.880 ;
        RECT  1.410 3.200 1.690 3.880 ;
        RECT  0.370 3.320 1.410 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 1.400 2.290 1.680 ;
        RECT  2.030 2.800 2.150 3.080 ;
        RECT  1.870 2.520 2.030 3.080 ;
        RECT  1.210 1.400 2.010 1.560 ;
        RECT  0.890 2.520 1.870 2.680 ;
        RECT  1.090 0.920 1.210 2.070 ;
        RECT  1.050 0.920 1.090 2.190 ;
        RECT  0.810 0.920 1.050 1.080 ;
        RECT  0.810 1.910 1.050 2.190 ;
        RECT  0.530 0.800 0.810 1.080 ;
    END
END AOI2BB2XLTR

MACRO AOI2BB2X4TR
    CLASS CORE ;
    FOREIGN AOI2BB2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.390 0.520 6.550 1.140 ;
        RECT  4.220 0.520 6.390 0.680 ;
        RECT  4.060 0.520 4.220 1.080 ;
        RECT  3.120 0.920 4.060 1.080 ;
        RECT  3.120 1.910 3.340 2.840 ;
        RECT  3.060 0.920 3.120 2.840 ;
        RECT  2.880 0.920 3.060 2.070 ;
        RECT  2.860 0.920 2.880 1.310 ;
        RECT  2.380 1.910 2.880 2.070 ;
        RECT  2.580 0.440 2.860 1.310 ;
        RECT  2.100 1.910 2.380 3.030 ;
        END
        ANTENNADIFFAREA 8.58 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.340 1.260 5.900 1.540 ;
        RECT  5.180 1.260 5.340 1.860 ;
        RECT  4.070 1.700 5.180 1.860 ;
        RECT  3.680 1.240 4.070 1.860 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.220 1.320 6.340 1.540 ;
        RECT  6.060 0.840 6.220 1.540 ;
        RECT  4.840 0.840 6.060 1.000 ;
        RECT  4.480 0.840 4.840 1.540 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 1.580 1.920 1.960 ;
        RECT  1.540 1.580 1.710 3.030 ;
        RECT  0.690 2.870 1.540 3.030 ;
        RECT  0.530 1.910 0.690 3.030 ;
        RECT  0.320 1.910 0.530 2.070 ;
        RECT  0.160 1.580 0.320 2.070 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.910 1.680 ;
        END
        ANTENNAGATEAREA 0.2952 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.700 -0.280 6.800 0.280 ;
        RECT  5.420 -0.280 5.700 0.360 ;
        RECT  3.900 -0.280 5.420 0.280 ;
        RECT  3.060 -0.280 3.900 0.760 ;
        RECT  2.380 -0.280 3.060 0.280 ;
        RECT  1.700 -0.280 2.380 0.800 ;
        RECT  0.960 -0.280 1.700 0.280 ;
        RECT  0.640 -0.280 0.960 0.800 ;
        RECT  0.000 -0.280 0.640 0.280 ;
        RECT  0.240 0.520 0.640 0.800 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.220 3.320 6.800 3.880 ;
        RECT  5.940 2.340 6.220 3.880 ;
        RECT  5.260 3.320 5.940 3.880 ;
        RECT  4.980 2.340 5.260 3.880 ;
        RECT  4.300 3.320 4.980 3.880 ;
        RECT  4.020 2.340 4.300 3.880 ;
        RECT  1.920 3.320 4.020 3.880 ;
        RECT  0.370 3.260 1.920 3.880 ;
        RECT  0.090 2.430 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.420 2.020 6.700 3.140 ;
        RECT  5.740 2.020 6.420 2.180 ;
        RECT  5.460 2.020 5.740 3.140 ;
        RECT  4.780 2.020 5.460 2.180 ;
        RECT  4.500 2.020 4.780 3.140 ;
        RECT  3.820 2.020 4.500 2.180 ;
        RECT  3.540 2.020 3.820 3.160 ;
        RECT  2.860 3.000 3.540 3.160 ;
        RECT  2.580 2.230 2.860 3.160 ;
        RECT  2.420 1.470 2.580 1.750 ;
        RECT  2.260 1.260 2.420 1.750 ;
        RECT  1.440 1.260 2.260 1.420 ;
        RECT  1.320 0.450 1.440 1.420 ;
        RECT  1.250 0.450 1.320 2.070 ;
        RECT  1.170 1.250 1.250 2.070 ;
        RECT  1.160 1.250 1.170 2.710 ;
        RECT  0.890 1.910 1.160 2.710 ;
    END
END AOI2BB2X4TR

MACRO AOI2BB2X2TR
    CLASS CORE ;
    FOREIGN AOI2BB2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 0.840 3.960 1.160 ;
        RECT  3.680 0.820 3.840 2.360 ;
        RECT  2.160 0.820 3.680 1.100 ;
        RECT  3.320 2.200 3.680 2.360 ;
        RECT  3.040 2.200 3.320 2.480 ;
        END
        ANTENNADIFFAREA 4.926 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.440 3.520 1.960 ;
        RECT  2.400 1.440 3.240 1.600 ;
        RECT  2.240 1.440 2.400 2.170 ;
        RECT  1.600 2.010 2.240 2.170 ;
        RECT  1.320 1.770 1.600 2.170 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 0.440 4.170 0.600 ;
        RECT  1.960 1.570 2.080 1.850 ;
        RECT  1.800 0.440 1.960 1.850 ;
        RECT  1.640 0.840 1.800 1.160 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.160 1.560 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.180 0.340 2.360 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 -0.280 4.400 0.280 ;
        RECT  1.120 -0.280 1.400 1.020 ;
        RECT  0.360 -0.280 1.120 0.340 ;
        RECT  0.140 -0.280 0.360 1.020 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.280 3.320 4.400 3.880 ;
        RECT  4.000 2.100 4.280 3.880 ;
        RECT  2.320 3.260 4.000 3.880 ;
        RECT  2.040 3.200 2.320 3.880 ;
        RECT  1.320 3.260 2.040 3.880 ;
        RECT  1.040 2.650 1.320 3.880 ;
        RECT  0.000 3.320 1.040 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.520 2.650 3.800 2.930 ;
        RECT  2.840 2.770 3.520 2.930 ;
        RECT  2.840 1.760 2.960 2.040 ;
        RECT  2.680 1.760 2.840 2.490 ;
        RECT  2.560 2.650 2.840 2.930 ;
        RECT  0.700 2.330 2.680 2.490 ;
        RECT  1.800 2.770 2.560 2.930 ;
        RECT  1.520 2.650 1.800 2.930 ;
        RECT  0.680 0.800 0.920 1.080 ;
        RECT  0.680 2.330 0.700 2.890 ;
        RECT  0.520 0.800 0.680 2.890 ;
        RECT  0.160 2.600 0.520 2.890 ;
    END
END AOI2BB2X2TR

MACRO AOI2BB2X1TR
    CLASS CORE ;
    FOREIGN AOI2BB2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.580 0.770 2.720 2.360 ;
        RECT  2.480 0.770 2.580 2.740 ;
        RECT  2.090 0.770 2.480 0.930 ;
        RECT  2.290 2.040 2.480 2.740 ;
        RECT  1.810 0.650 2.090 0.930 ;
        END
        ANTENNADIFFAREA 2.584 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.660 0.720 3.160 ;
        END
        ANTENNAGATEAREA 0.1584 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.640 1.960 1.960 ;
        RECT  1.660 1.410 1.850 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.180 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.210 1.120 1.560 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.280 2.800 0.280 ;
        RECT  0.970 -0.280 1.250 0.400 ;
        RECT  0.090 -0.280 0.970 0.340 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.680 3.320 2.800 3.880 ;
        RECT  1.400 3.170 1.680 3.880 ;
        RECT  0.310 3.320 1.400 3.880 ;
        RECT  0.120 2.600 0.310 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 1.090 2.290 1.440 ;
        RECT  1.800 2.130 2.090 2.770 ;
        RECT  1.500 1.090 2.010 1.250 ;
        RECT  1.150 2.490 1.800 2.770 ;
        RECT  1.340 0.860 1.500 2.190 ;
        RECT  0.810 0.860 1.340 1.020 ;
        RECT  0.820 1.930 1.340 2.190 ;
        RECT  0.880 2.490 1.150 3.110 ;
        RECT  0.530 0.740 0.810 1.020 ;
    END
END AOI2BB2X1TR

MACRO AOI2BB1XLTR
    CLASS CORE ;
    FOREIGN AOI2BB1XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.940 2.320 3.160 ;
        RECT  1.820 0.940 2.160 1.100 ;
        RECT  2.080 1.910 2.160 3.160 ;
        RECT  2.000 1.910 2.080 2.360 ;
        RECT  1.540 0.820 1.820 1.100 ;
        END
        ANTENNADIFFAREA 1.716 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.580 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.580 1.060 1.860 ;
        RECT  0.480 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  0.380 -0.280 2.220 0.340 ;
        RECT  0.100 -0.280 0.380 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.820 3.320 2.400 3.880 ;
        RECT  1.360 3.260 1.820 3.880 ;
        RECT  1.060 2.700 1.360 3.880 ;
        RECT  0.370 3.260 1.060 3.880 ;
        RECT  0.000 3.320 0.370 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.260 2.000 1.610 ;
        RECT  1.680 1.260 1.840 2.540 ;
        RECT  0.820 1.260 1.680 1.420 ;
        RECT  0.500 2.380 1.680 2.540 ;
        RECT  0.660 1.000 0.820 1.420 ;
        RECT  0.540 1.000 0.660 1.280 ;
        RECT  0.220 2.380 0.500 2.660 ;
    END
END AOI2BB1XLTR

MACRO AOI2BB1X4TR
    CLASS CORE ;
    FOREIGN AOI2BB1X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.920 4.260 3.160 ;
        RECT  3.810 0.920 4.000 1.160 ;
        RECT  3.960 2.120 4.000 3.160 ;
        RECT  3.680 2.120 3.960 2.990 ;
        RECT  3.530 0.440 3.810 1.160 ;
        RECT  2.690 2.120 3.680 2.360 ;
        RECT  2.850 0.920 3.530 1.160 ;
        RECT  2.570 0.440 2.850 1.160 ;
        RECT  2.410 2.120 2.690 2.950 ;
        END
        ANTENNADIFFAREA 7.12 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.700 3.290 1.960 ;
        RECT  2.840 1.640 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.624 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.640 1.960 1.960 ;
        RECT  1.410 1.640 1.570 2.800 ;
        RECT  0.320 2.640 1.410 2.800 ;
        RECT  0.160 1.710 0.320 2.800 ;
        RECT  0.100 1.710 0.160 1.990 ;
        END
        ANTENNAGATEAREA 0.2856 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.640 0.890 1.960 ;
        END
        ANTENNAGATEAREA 0.2856 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.280 4.400 0.280 ;
        RECT  4.010 -0.280 4.290 0.670 ;
        RECT  3.330 -0.280 4.010 0.280 ;
        RECT  3.050 -0.280 3.330 0.670 ;
        RECT  2.370 -0.280 3.050 0.280 ;
        RECT  2.090 -0.280 2.370 1.160 ;
        RECT  1.090 -0.280 2.090 0.280 ;
        RECT  0.810 -0.280 1.090 1.160 ;
        RECT  0.000 -0.280 0.810 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.490 3.320 4.400 3.880 ;
        RECT  3.210 2.520 3.490 3.880 ;
        RECT  1.850 3.320 3.210 3.880 ;
        RECT  1.570 3.200 1.850 3.880 ;
        RECT  0.370 3.260 1.570 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.560 1.320 3.840 1.650 ;
        RECT  2.490 1.320 3.560 1.480 ;
        RECT  2.210 1.320 2.490 1.960 ;
        RECT  1.570 1.320 2.210 1.480 ;
        RECT  1.290 0.520 1.570 1.480 ;
        RECT  1.210 1.320 1.290 1.480 ;
        RECT  1.050 1.320 1.210 2.450 ;
        RECT  0.610 1.320 1.050 1.480 ;
        RECT  0.810 2.120 1.050 2.450 ;
        RECT  0.330 0.520 0.610 1.480 ;
    END
END AOI2BB1X4TR

MACRO AOI2BB1X2TR
    CLASS CORE ;
    FOREIGN AOI2BB1X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.030 1.990 2.760 ;
        RECT  1.680 2.440 1.770 2.760 ;
        END
        ANTENNADIFFAREA 3.556 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.640 2.720 2.760 ;
        RECT  2.350 1.640 2.470 1.960 ;
        RECT  2.190 0.710 2.350 1.960 ;
        RECT  1.610 0.710 2.190 0.870 ;
        RECT  1.390 0.710 1.610 1.640 ;
        END
        ANTENNAGATEAREA 0.3024 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.520 0.910 1.960 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.440 0.320 1.740 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.280 2.800 0.280 ;
        RECT  2.230 -0.280 2.510 0.340 ;
        RECT  1.370 -0.280 2.230 0.280 ;
        RECT  1.090 -0.280 1.370 0.400 ;
        RECT  0.540 -0.280 1.090 0.340 ;
        RECT  0.000 -0.280 0.540 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.430 3.260 2.710 3.880 ;
        RECT  1.150 3.320 2.430 3.880 ;
        RECT  0.870 3.260 1.150 3.880 ;
        RECT  0.000 3.320 0.870 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.520 2.940 2.190 3.160 ;
        RECT  1.230 2.940 1.520 3.100 ;
        RECT  1.070 0.980 1.230 3.100 ;
        RECT  0.790 0.980 1.070 1.140 ;
        RECT  0.310 2.940 1.070 3.100 ;
        RECT  0.510 0.860 0.790 1.140 ;
        RECT  0.150 2.030 0.310 3.100 ;
        RECT  0.090 2.030 0.150 2.830 ;
    END
END AOI2BB1X2TR

MACRO AOI2BB1X1TR
    CLASS CORE ;
    FOREIGN AOI2BB1X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.940 2.320 3.160 ;
        RECT  1.820 0.940 2.160 1.100 ;
        RECT  2.070 1.910 2.160 3.160 ;
        RECT  2.000 1.910 2.070 2.770 ;
        RECT  1.540 0.820 1.820 1.100 ;
        END
        ANTENNADIFFAREA 2.508 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.580 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.580 1.120 2.360 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0744 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  0.420 -0.280 2.220 0.340 ;
        RECT  0.140 -0.280 0.420 0.750 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.820 3.320 2.400 3.880 ;
        RECT  1.360 3.260 1.820 3.880 ;
        RECT  1.060 2.860 1.360 3.880 ;
        RECT  0.370 3.260 1.060 3.880 ;
        RECT  0.000 3.320 0.370 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.260 2.000 1.610 ;
        RECT  1.680 1.260 1.840 2.680 ;
        RECT  1.040 1.260 1.680 1.420 ;
        RECT  0.500 2.520 1.680 2.680 ;
        RECT  0.880 1.000 1.040 1.420 ;
        RECT  0.580 1.000 0.880 1.280 ;
        RECT  0.220 2.120 0.500 2.680 ;
    END
END AOI2BB1X1TR

MACRO AOI22XLTR
    CLASS CORE ;
    FOREIGN AOI22XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 0.840 2.320 2.280 ;
        RECT  0.890 0.920 2.080 1.080 ;
        RECT  1.810 2.120 2.080 2.280 ;
        RECT  1.530 2.120 1.810 2.550 ;
        END
        ANTENNADIFFAREA 1.7195 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.840 0.510 1.480 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        RECT  0.480 1.640 0.880 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 -0.280 2.400 0.280 ;
        RECT  1.810 -0.280 2.090 0.350 ;
        RECT  0.370 -0.280 1.810 0.290 ;
        RECT  0.090 -0.280 0.370 0.370 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 3.320 2.400 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.170 2.440 2.290 2.690 ;
        RECT  2.010 2.440 2.170 3.100 ;
        RECT  1.330 2.940 2.010 3.100 ;
        RECT  1.170 2.120 1.330 3.100 ;
        RECT  1.050 2.120 1.170 2.550 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.580 ;
    END
END AOI22XLTR

MACRO AOI22X4TR
    CLASS CORE ;
    FOREIGN AOI22X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.820 0.590 5.920 1.360 ;
        RECT  5.580 0.590 5.820 2.840 ;
        RECT  5.460 0.590 5.580 1.160 ;
        RECT  5.480 2.120 5.580 2.840 ;
        RECT  4.800 2.120 5.480 2.360 ;
        RECT  4.000 0.920 5.460 1.160 ;
        RECT  4.520 2.120 4.800 2.840 ;
        RECT  3.840 2.120 4.520 2.360 ;
        RECT  3.720 0.440 4.000 1.160 ;
        RECT  3.560 2.120 3.840 2.840 ;
        RECT  2.310 0.580 3.720 0.820 ;
        RECT  2.030 0.500 2.310 1.060 ;
        RECT  0.640 0.580 2.030 0.820 ;
        RECT  0.630 0.510 0.640 0.820 ;
        RECT  0.350 0.510 0.630 1.070 ;
        END
        ANTENNADIFFAREA 12.062 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.220 2.920 1.560 ;
        RECT  1.550 1.220 2.440 1.380 ;
        RECT  1.390 1.220 1.550 1.560 ;
        RECT  0.950 1.280 1.390 1.560 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.540 2.280 1.820 ;
        RECT  1.830 1.540 1.990 1.880 ;
        RECT  0.760 1.720 1.830 1.880 ;
        RECT  0.390 1.240 0.760 1.880 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.720 1.320 5.000 1.600 ;
        RECT  3.560 1.320 4.720 1.480 ;
        RECT  3.200 1.240 3.560 1.880 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.260 1.380 5.420 1.960 ;
        RECT  4.520 1.800 5.260 1.960 ;
        RECT  3.840 1.640 4.520 1.960 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.840 -0.280 6.400 0.280 ;
        RECT  4.560 -0.280 4.840 0.680 ;
        RECT  3.160 -0.280 4.560 0.280 ;
        RECT  2.880 -0.280 3.160 0.400 ;
        RECT  1.470 -0.280 2.880 0.280 ;
        RECT  1.190 -0.280 1.470 0.400 ;
        RECT  0.000 -0.280 1.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.790 3.320 6.400 3.880 ;
        RECT  2.510 2.640 2.790 3.880 ;
        RECT  1.830 3.260 2.510 3.880 ;
        RECT  1.550 2.610 1.830 3.880 ;
        RECT  0.950 3.260 1.550 3.880 ;
        RECT  0.670 3.200 0.950 3.880 ;
        RECT  0.000 3.320 0.670 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.980 2.050 6.240 3.160 ;
        RECT  5.280 3.000 5.980 3.160 ;
        RECT  5.000 2.540 5.280 3.160 ;
        RECT  4.320 3.000 5.000 3.160 ;
        RECT  4.040 2.540 4.320 3.160 ;
        RECT  3.270 3.000 4.040 3.160 ;
        RECT  2.990 2.040 3.270 3.160 ;
        RECT  2.310 2.040 2.990 2.200 ;
        RECT  2.030 2.040 2.310 2.920 ;
        RECT  1.350 2.040 2.030 2.200 ;
        RECT  1.070 2.040 1.350 2.890 ;
        RECT  0.430 2.040 1.070 2.200 ;
        RECT  0.150 2.040 0.430 3.160 ;
    END
END AOI22X4TR

MACRO AOI22X2TR
    CLASS CORE ;
    FOREIGN AOI22X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.150 0.920 4.310 2.200 ;
        RECT  3.350 0.920 4.150 1.080 ;
        RECT  3.920 2.040 4.150 2.200 ;
        RECT  3.830 2.040 3.920 2.360 ;
        RECT  3.640 2.040 3.830 2.750 ;
        RECT  3.550 2.120 3.640 2.750 ;
        RECT  2.870 2.120 3.550 2.280 ;
        RECT  3.070 0.800 3.350 1.080 ;
        RECT  1.470 0.920 3.070 1.080 ;
        RECT  2.590 2.120 2.870 2.750 ;
        RECT  1.190 0.800 1.470 1.080 ;
        END
        ANTENNADIFFAREA 5.184 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.240 2.110 1.640 ;
        RECT  0.790 1.240 1.830 1.400 ;
        RECT  0.440 1.240 0.790 1.640 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.580 1.670 1.860 ;
        RECT  1.240 1.580 1.560 1.960 ;
        RECT  0.990 1.580 1.240 1.860 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.710 1.240 3.990 1.640 ;
        RECT  2.720 1.240 3.710 1.400 ;
        RECT  2.390 1.240 2.720 1.640 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.580 3.550 1.860 ;
        RECT  2.880 1.580 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.190 -0.280 4.400 0.280 ;
        RECT  3.910 -0.280 4.190 0.760 ;
        RECT  2.350 -0.280 3.910 0.340 ;
        RECT  2.070 -0.280 2.350 0.760 ;
        RECT  0.670 -0.280 2.070 0.340 ;
        RECT  0.390 -0.280 0.670 0.990 ;
        RECT  0.000 -0.280 0.390 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 3.320 4.400 3.880 ;
        RECT  1.590 3.200 1.870 3.880 ;
        RECT  0.990 3.260 1.590 3.880 ;
        RECT  0.710 2.470 0.990 3.880 ;
        RECT  0.000 3.320 0.710 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.250 2.470 4.310 2.750 ;
        RECT  4.090 2.470 4.250 3.070 ;
        RECT  3.350 2.910 4.090 3.070 ;
        RECT  3.070 2.470 3.350 3.070 ;
        RECT  2.390 2.910 3.070 3.070 ;
        RECT  2.230 2.120 2.390 3.070 ;
        RECT  2.110 2.120 2.230 2.750 ;
        RECT  1.470 2.120 2.110 2.280 ;
        RECT  1.190 2.120 1.470 2.750 ;
        RECT  0.510 2.120 1.190 2.280 ;
        RECT  0.230 2.120 0.510 2.750 ;
    END
END AOI22X2TR

MACRO AOI22X1TR
    CLASS CORE ;
    FOREIGN AOI22X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.240 2.320 2.360 ;
        RECT  2.080 0.840 2.240 2.360 ;
        RECT  0.890 0.840 2.080 1.000 ;
        RECT  1.810 2.120 2.080 2.280 ;
        RECT  1.530 2.120 1.810 2.780 ;
        END
        ANTENNADIFFAREA 2.802 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.720 0.590 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.640 ;
        RECT  0.480 1.240 0.880 1.560 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.850 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.280 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.080 -0.280 2.400 0.280 ;
        RECT  1.800 -0.280 2.080 0.680 ;
        RECT  0.370 -0.280 1.800 0.290 ;
        RECT  0.090 -0.280 0.370 0.970 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 3.320 2.400 3.880 ;
        RECT  0.570 3.250 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.170 2.570 2.290 2.850 ;
        RECT  2.010 2.570 2.170 3.100 ;
        RECT  1.330 2.940 2.010 3.100 ;
        RECT  1.170 2.120 1.330 3.100 ;
        RECT  1.050 2.120 1.170 2.850 ;
        RECT  0.640 2.120 1.050 2.280 ;
        RECT  0.480 2.120 0.640 2.680 ;
        RECT  0.370 2.520 0.480 2.680 ;
        RECT  0.090 2.520 0.370 2.850 ;
    END
END AOI22X1TR

MACRO AOI222XLTR
    CLASS CORE ;
    FOREIGN AOI222XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 0.800 3.400 1.080 ;
        RECT  3.120 2.650 3.390 2.930 ;
        RECT  3.060 0.920 3.120 1.080 ;
        RECT  3.060 2.040 3.120 2.930 ;
        RECT  2.880 0.920 3.060 2.930 ;
        RECT  1.620 0.920 2.880 1.080 ;
        RECT  1.310 0.800 1.620 1.080 ;
        END
        ANTENNADIFFAREA 3.6725 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.240 0.720 1.620 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.490 1.120 2.000 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.880 1.560 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 1.620 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.240 3.520 2.360 ;
        RECT  3.260 1.240 3.280 1.500 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 -0.280 3.600 0.280 ;
        RECT  2.280 -0.280 2.560 0.760 ;
        RECT  0.740 -0.280 2.280 0.280 ;
        RECT  0.460 -0.280 0.740 1.080 ;
        RECT  0.000 -0.280 0.460 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 3.320 3.600 3.880 ;
        RECT  0.920 3.240 1.230 3.880 ;
        RECT  0.370 3.320 0.920 3.880 ;
        RECT  0.090 2.890 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.410 2.770 2.680 3.050 ;
        RECT  0.860 2.160 2.090 2.320 ;
        RECT  0.590 2.160 0.860 2.440 ;
    END
END AOI222XLTR

MACRO AOI222X4TR
    CLASS CORE ;
    FOREIGN AOI222X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.030 1.040 5.120 2.070 ;
        RECT  4.770 0.440 5.030 3.160 ;
        RECT  4.750 0.440 4.770 1.310 ;
        RECT  4.750 1.910 4.770 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.270 0.550 1.560 ;
        RECT  0.320 1.240 0.360 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.160 1.870 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.240 1.920 1.560 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.790 1.870 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.440 3.560 0.760 ;
        RECT  2.890 0.480 3.240 0.760 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 -0.280 5.600 0.280 ;
        RECT  5.230 -0.280 5.510 0.760 ;
        RECT  4.550 -0.280 5.230 0.280 ;
        RECT  4.270 -0.280 4.550 0.850 ;
        RECT  2.530 -0.280 4.270 0.280 ;
        RECT  2.250 -0.280 2.530 0.760 ;
        RECT  0.800 -0.280 2.250 0.340 ;
        RECT  0.520 -0.280 0.800 1.080 ;
        RECT  0.000 -0.280 0.520 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 3.320 5.600 3.880 ;
        RECT  5.230 2.230 5.510 3.880 ;
        RECT  4.550 3.320 5.230 3.880 ;
        RECT  4.270 2.230 4.550 3.880 ;
        RECT  1.230 3.260 4.270 3.880 ;
        RECT  0.950 3.200 1.230 3.880 ;
        RECT  0.430 3.320 0.950 3.880 ;
        RECT  0.150 3.200 0.430 3.880 ;
        RECT  0.000 3.320 0.150 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.590 1.470 4.610 1.750 ;
        RECT  4.430 1.150 4.590 2.070 ;
        RECT  4.070 1.150 4.430 1.310 ;
        RECT  4.070 1.910 4.430 2.070 ;
        RECT  3.370 1.470 4.270 1.750 ;
        RECT  3.790 0.570 4.070 1.310 ;
        RECT  3.790 1.910 4.070 2.930 ;
        RECT  3.490 1.970 3.610 2.630 ;
        RECT  3.330 1.970 3.490 2.950 ;
        RECT  3.170 0.920 3.370 1.750 ;
        RECT  2.650 2.790 3.330 2.950 ;
        RECT  3.010 0.920 3.170 2.630 ;
        RECT  1.690 0.920 3.010 1.080 ;
        RECT  2.850 2.030 3.010 2.630 ;
        RECT  2.370 2.170 2.650 2.950 ;
        RECT  1.690 2.790 2.370 2.950 ;
        RECT  1.890 2.120 2.170 2.630 ;
        RECT  0.830 2.120 1.890 2.280 ;
        RECT  1.410 0.800 1.690 1.080 ;
        RECT  1.530 2.440 1.690 2.950 ;
        RECT  1.410 2.440 1.530 2.630 ;
        RECT  0.550 2.120 0.830 2.690 ;
    END
END AOI222X4TR

MACRO AOI222X2TR
    CLASS CORE ;
    FOREIGN AOI222X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.540 2.120 5.820 2.780 ;
        RECT  4.860 2.120 5.540 2.280 ;
        RECT  4.800 0.840 5.160 1.160 ;
        RECT  4.800 2.120 4.860 2.780 ;
        RECT  4.720 0.840 4.800 2.780 ;
        RECT  4.640 1.000 4.720 2.780 ;
        RECT  3.400 1.000 4.640 1.160 ;
        RECT  3.120 0.840 3.400 1.160 ;
        RECT  2.040 1.000 3.120 1.160 ;
        RECT  1.880 0.730 2.040 1.160 ;
        RECT  1.340 0.730 1.880 0.890 ;
        RECT  1.060 0.610 1.340 0.890 ;
        END
        ANTENNADIFFAREA 6.948 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.320 1.940 1.600 ;
        RECT  1.560 1.050 1.720 1.600 ;
        RECT  0.720 1.050 1.560 1.210 ;
        RECT  0.440 1.050 0.720 1.630 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.370 1.400 1.650 ;
        RECT  0.880 1.370 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.320 4.040 1.600 ;
        RECT  2.760 1.320 3.760 1.480 ;
        RECT  2.480 1.320 2.760 1.960 ;
        RECT  2.440 1.320 2.480 1.600 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.640 3.600 1.920 ;
        RECT  3.240 1.640 3.560 1.960 ;
        RECT  2.920 1.640 3.240 1.920 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.240 5.960 1.890 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.230 1.640 5.520 1.960 ;
        RECT  5.040 1.380 5.230 1.960 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.880 -0.280 6.400 0.280 ;
        RECT  5.600 -0.280 5.880 0.990 ;
        RECT  4.240 -0.280 5.600 0.280 ;
        RECT  3.960 -0.280 4.240 0.840 ;
        RECT  2.480 -0.280 3.960 0.280 ;
        RECT  2.200 -0.280 2.480 0.840 ;
        RECT  0.540 -0.280 2.200 0.280 ;
        RECT  0.260 -0.280 0.540 0.890 ;
        RECT  0.000 -0.280 0.260 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.320 6.400 3.880 ;
        RECT  1.940 2.990 2.220 3.880 ;
        RECT  1.380 3.320 1.940 3.880 ;
        RECT  1.100 3.240 1.380 3.880 ;
        RECT  0.380 3.320 1.100 3.880 ;
        RECT  0.100 2.090 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.020 2.100 6.300 3.100 ;
        RECT  5.340 2.940 6.020 3.100 ;
        RECT  5.060 2.470 5.340 3.100 ;
        RECT  4.360 2.940 5.060 3.100 ;
        RECT  4.080 2.120 4.360 3.100 ;
        RECT  3.400 2.120 4.080 2.280 ;
        RECT  3.600 2.440 3.880 3.100 ;
        RECT  2.920 2.940 3.600 3.100 ;
        RECT  3.120 2.120 3.400 2.780 ;
        RECT  2.320 2.120 3.120 2.280 ;
        RECT  2.760 2.470 2.920 3.100 ;
        RECT  2.640 2.470 2.760 2.770 ;
        RECT  1.740 2.610 2.640 2.770 ;
        RECT  2.160 1.720 2.320 2.280 ;
        RECT  2.100 1.720 2.160 2.000 ;
        RECT  1.460 2.120 1.740 2.770 ;
        RECT  0.860 2.120 1.460 2.280 ;
        RECT  0.580 2.120 0.860 3.160 ;
    END
END AOI222X2TR

MACRO AOI222X1TR
    CLASS CORE ;
    FOREIGN AOI222X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.800 3.720 1.080 ;
        RECT  3.280 0.800 3.440 2.780 ;
        RECT  2.000 0.800 3.280 0.960 ;
        RECT  3.120 2.160 3.280 2.780 ;
        RECT  1.680 0.800 2.000 1.160 ;
        END
        ANTENNADIFFAREA 3.876 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.410 0.720 1.660 ;
        RECT  0.080 0.440 0.330 1.660 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.720 1.140 1.960 ;
        RECT  0.880 1.530 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.210 2.720 1.640 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.400 2.200 1.680 ;
        RECT  1.520 1.400 1.920 1.560 ;
        RECT  1.280 1.240 1.520 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.370 3.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.240 3.920 2.360 ;
        RECT  3.600 1.240 3.680 1.670 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.880 -0.280 4.000 0.280 ;
        RECT  2.600 -0.280 2.880 0.640 ;
        RECT  1.200 -0.280 2.600 0.340 ;
        RECT  0.920 -0.280 1.200 0.990 ;
        RECT  0.000 -0.280 0.920 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 3.320 4.000 3.880 ;
        RECT  1.200 2.480 1.480 3.880 ;
        RECT  0.520 3.320 1.200 3.880 ;
        RECT  0.240 2.050 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.600 2.640 3.880 3.100 ;
        RECT  2.920 2.940 3.600 3.100 ;
        RECT  2.640 2.300 2.920 3.100 ;
        RECT  1.960 2.940 2.640 3.100 ;
        RECT  2.160 1.910 2.440 2.780 ;
        RECT  1.520 1.910 2.160 2.070 ;
        RECT  1.680 2.230 1.960 3.100 ;
        RECT  1.360 1.910 1.520 2.320 ;
        RECT  1.000 2.160 1.360 2.320 ;
        RECT  0.720 2.160 1.000 3.070 ;
    END
END AOI222X1TR

MACRO AOI221XLTR
    CLASS CORE ;
    FOREIGN AOI221XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.920 3.120 3.040 ;
        RECT  2.960 0.800 3.040 3.040 ;
        RECT  2.760 0.800 2.960 1.080 ;
        RECT  2.880 1.640 2.960 3.040 ;
        RECT  2.720 2.760 2.880 3.040 ;
        RECT  1.520 0.920 2.760 1.080 ;
        RECT  1.250 0.800 1.520 1.080 ;
        END
        ANTENNADIFFAREA 3.05 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 1.770 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.230 0.720 1.610 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.470 1.120 2.000 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.810 1.560 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 -0.280 3.200 0.280 ;
        RECT  2.200 -0.280 2.480 0.760 ;
        RECT  0.640 -0.280 2.200 0.280 ;
        RECT  0.360 -0.280 0.640 1.070 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 3.320 3.200 3.880 ;
        RECT  1.000 3.200 1.280 3.880 ;
        RECT  0.420 3.260 1.000 3.880 ;
        RECT  0.140 3.200 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.460 2.760 2.540 3.040 ;
        RECT  0.880 2.160 2.140 2.320 ;
        RECT  0.600 2.160 0.880 2.440 ;
    END
END AOI221XLTR

MACRO AOI221X4TR
    CLASS CORE ;
    FOREIGN AOI221X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.600 1.150 4.720 2.170 ;
        RECT  4.480 0.440 4.600 3.160 ;
        RECT  4.320 0.440 4.480 1.310 ;
        RECT  4.320 1.910 4.480 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.880 1.560 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.170 0.580 1.450 ;
        RECT  0.320 0.840 0.360 1.450 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.160 1.770 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.240 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.560 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.080 -0.280 5.200 0.280 ;
        RECT  4.800 -0.280 5.080 0.990 ;
        RECT  4.120 -0.280 4.800 0.280 ;
        RECT  3.840 -0.280 4.120 0.850 ;
        RECT  2.560 -0.280 3.840 0.340 ;
        RECT  2.280 -0.280 2.560 0.760 ;
        RECT  0.800 -0.280 2.280 0.340 ;
        RECT  0.520 -0.280 0.800 1.000 ;
        RECT  0.000 -0.280 0.520 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.080 3.320 5.200 3.880 ;
        RECT  4.800 2.510 5.080 3.880 ;
        RECT  4.120 3.320 4.800 3.880 ;
        RECT  3.840 2.230 4.120 3.880 ;
        RECT  1.260 3.260 3.840 3.880 ;
        RECT  0.980 3.200 1.260 3.880 ;
        RECT  0.460 3.320 0.980 3.880 ;
        RECT  0.180 3.200 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.160 1.470 4.320 1.750 ;
        RECT  4.000 1.150 4.160 2.070 ;
        RECT  3.640 1.150 4.000 1.310 ;
        RECT  3.640 1.910 4.000 2.070 ;
        RECT  3.200 1.470 3.840 1.750 ;
        RECT  3.360 0.570 3.640 1.310 ;
        RECT  3.360 1.910 3.640 2.930 ;
        RECT  3.040 0.800 3.200 2.400 ;
        RECT  2.800 0.800 3.040 1.080 ;
        RECT  2.880 2.040 3.040 2.400 ;
        RECT  1.720 0.920 2.800 1.080 ;
        RECT  2.400 2.120 2.680 2.570 ;
        RECT  1.720 2.120 2.400 2.280 ;
        RECT  1.920 2.440 2.200 2.890 ;
        RECT  0.860 2.730 1.920 2.890 ;
        RECT  1.440 0.800 1.720 1.080 ;
        RECT  1.440 2.120 1.720 2.570 ;
        RECT  0.580 2.140 0.860 2.890 ;
    END
END AOI221X4TR

MACRO AOI221X2TR
    CLASS CORE ;
    FOREIGN AOI221X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.950 1.910 5.120 2.840 ;
        RECT  4.750 0.920 4.950 2.840 ;
        RECT  4.670 0.920 4.750 1.200 ;
        RECT  3.590 0.920 4.670 1.080 ;
        RECT  3.310 0.800 3.590 1.080 ;
        RECT  1.400 0.920 3.310 1.080 ;
        RECT  1.120 0.800 1.400 1.080 ;
        END
        ANTENNADIFFAREA 4.842 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.240 5.520 2.360 ;
        RECT  5.110 1.240 5.280 1.610 ;
        END
        ANTENNAGATEAREA 0.3576 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.240 2.080 1.590 ;
        RECT  0.720 1.240 1.810 1.400 ;
        RECT  0.440 1.240 0.720 1.590 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.560 1.240 1.960 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.240 4.230 1.590 ;
        RECT  3.120 1.240 3.950 1.400 ;
        RECT  2.630 1.240 3.120 1.590 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.580 3.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.430 -0.280 5.600 0.280 ;
        RECT  5.150 -0.280 5.430 1.080 ;
        RECT  4.430 -0.280 5.150 0.280 ;
        RECT  4.150 -0.280 4.430 0.760 ;
        RECT  2.670 -0.280 4.150 0.280 ;
        RECT  2.040 -0.280 2.670 0.760 ;
        RECT  0.600 -0.280 2.040 0.280 ;
        RECT  0.320 -0.280 0.600 0.940 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 3.320 5.600 3.880 ;
        RECT  2.000 2.530 2.280 3.880 ;
        RECT  1.440 3.260 2.000 3.880 ;
        RECT  1.160 3.200 1.440 3.880 ;
        RECT  0.440 3.320 1.160 3.880 ;
        RECT  0.160 1.920 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.450 2.630 5.510 2.940 ;
        RECT  5.290 2.630 5.450 3.160 ;
        RECT  4.550 3.000 5.290 3.160 ;
        RECT  4.270 1.910 4.550 3.160 ;
        RECT  3.590 3.000 4.270 3.160 ;
        RECT  3.790 2.120 4.070 2.840 ;
        RECT  3.110 2.120 3.790 2.280 ;
        RECT  3.310 2.440 3.590 3.160 ;
        RECT  2.630 3.000 3.310 3.160 ;
        RECT  2.990 2.120 3.110 2.840 ;
        RECT  2.830 1.750 2.990 2.840 ;
        RECT  1.800 1.750 2.830 1.910 ;
        RECT  2.470 2.070 2.630 3.160 ;
        RECT  2.350 2.070 2.470 2.350 ;
        RECT  1.640 1.750 1.800 2.730 ;
        RECT  1.520 2.120 1.640 2.730 ;
        RECT  0.920 2.120 1.520 2.280 ;
        RECT  0.640 2.120 0.920 3.160 ;
    END
END AOI221X2TR

MACRO AOI221X1TR
    CLASS CORE ;
    FOREIGN AOI221X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.920 3.120 2.870 ;
        RECT  1.670 0.920 2.880 1.080 ;
        RECT  0.990 0.800 1.670 1.080 ;
        END
        ANTENNADIFFAREA 4.648 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 1.010 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.240 2.320 1.650 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.810 1.560 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 -0.280 3.200 0.280 ;
        RECT  2.260 -0.280 2.540 0.740 ;
        RECT  0.430 -0.280 2.260 0.280 ;
        RECT  0.150 -0.280 0.430 0.550 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 3.320 3.200 3.880 ;
        RECT  1.050 2.760 1.330 3.880 ;
        RECT  0.350 3.260 1.050 3.880 ;
        RECT  0.090 2.200 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 2.120 2.630 2.740 ;
        RECT  1.610 2.440 2.350 2.600 ;
        RECT  1.990 2.120 2.150 2.280 ;
        RECT  1.830 1.810 1.990 2.280 ;
        RECT  0.850 1.810 1.830 1.970 ;
        RECT  1.450 2.130 1.610 2.600 ;
        RECT  0.570 1.810 0.850 2.820 ;
    END
END AOI221X1TR

MACRO AOI21XLTR
    CLASS CORE ;
    FOREIGN AOI21XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.840 1.920 1.960 ;
        RECT  1.680 0.840 1.840 2.560 ;
        RECT  1.370 0.920 1.680 1.080 ;
        RECT  1.530 2.280 1.680 2.560 ;
        RECT  0.970 0.800 1.370 1.080 ;
        END
        ANTENNADIFFAREA 1.44 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.460 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.0816 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.590 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.240 1.120 1.870 ;
        END
        ANTENNAGATEAREA 0.1008 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.280 2.000 0.280 ;
        RECT  1.530 -0.280 1.810 0.680 ;
        RECT  0.390 -0.280 1.530 0.280 ;
        RECT  0.100 -0.280 0.390 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 3.320 2.000 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 2.120 1.330 2.560 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.560 ;
    END
END AOI21XLTR

MACRO AOI21X4TR
    CLASS CORE ;
    FOREIGN AOI21X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 0.930 4.700 3.040 ;
        RECT  4.320 0.930 4.400 2.160 ;
        RECT  3.440 2.750 4.400 3.040 ;
        RECT  4.080 1.090 4.320 2.160 ;
        RECT  3.640 1.090 4.080 1.330 ;
        RECT  3.360 0.840 3.640 1.330 ;
        RECT  2.260 0.840 3.360 1.080 ;
        RECT  1.960 0.440 2.260 1.080 ;
        RECT  0.530 0.840 1.960 1.080 ;
        RECT  0.260 0.500 0.530 1.210 ;
        END
        ANTENNADIFFAREA 8.64 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.560 3.920 1.960 ;
        RECT  3.280 1.640 3.320 1.960 ;
        END
        ANTENNAGATEAREA 0.624 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.240 2.840 1.560 ;
        RECT  1.550 1.240 2.470 1.400 ;
        RECT  0.880 1.240 1.550 1.560 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.580 2.210 1.880 ;
        RECT  0.720 1.720 1.920 1.880 ;
        RECT  0.440 1.470 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.6984 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 -0.280 4.800 0.280 ;
        RECT  3.860 -0.280 4.140 0.920 ;
        RECT  3.110 -0.280 3.860 0.280 ;
        RECT  2.830 -0.280 3.110 0.670 ;
        RECT  1.380 -0.280 2.830 0.280 ;
        RECT  1.100 -0.280 1.380 0.660 ;
        RECT  0.000 -0.280 1.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.760 3.320 4.800 3.880 ;
        RECT  2.480 3.200 2.760 3.880 ;
        RECT  1.720 3.320 2.480 3.880 ;
        RECT  1.440 3.200 1.720 3.880 ;
        RECT  0.800 3.320 1.440 3.880 ;
        RECT  0.520 3.200 0.800 3.880 ;
        RECT  0.000 3.320 0.520 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.200 2.430 4.220 2.590 ;
        RECT  2.970 2.120 3.200 2.890 ;
        RECT  2.240 2.120 2.970 2.280 ;
        RECT  1.960 2.120 2.240 2.940 ;
        RECT  1.320 2.120 1.960 2.280 ;
        RECT  1.040 2.120 1.320 2.890 ;
        RECT  0.410 2.120 1.040 2.280 ;
        RECT  0.130 2.120 0.410 2.770 ;
    END
END AOI21X4TR

MACRO AOI21X2TR
    CLASS CORE ;
    FOREIGN AOI21X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 0.980 3.400 1.400 ;
        RECT  3.040 1.240 3.120 1.560 ;
        RECT  2.880 1.240 3.040 2.570 ;
        RECT  2.440 1.240 2.880 1.400 ;
        RECT  2.750 2.170 2.880 2.570 ;
        RECT  2.280 0.840 2.440 1.400 ;
        RECT  2.160 0.840 2.280 1.120 ;
        RECT  0.760 0.960 2.160 1.120 ;
        RECT  0.480 0.840 0.760 1.120 ;
        END
        ANTENNADIFFAREA 4.212 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.560 2.720 1.960 ;
        END
        ANTENNAGATEAREA 0.312 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.600 1.790 1.960 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.560 2.240 1.840 ;
        RECT  1.960 1.280 2.120 1.840 ;
        RECT  0.830 1.280 1.960 1.440 ;
        RECT  0.760 1.280 0.830 1.880 ;
        RECT  0.670 1.280 0.760 1.960 ;
        RECT  0.440 1.600 0.670 1.960 ;
        END
        ANTENNAGATEAREA 0.3456 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.920 -0.280 3.600 0.280 ;
        RECT  2.640 -0.280 2.920 1.080 ;
        RECT  1.600 -0.280 2.640 0.280 ;
        RECT  1.320 -0.280 1.600 0.800 ;
        RECT  0.000 -0.280 1.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 3.320 3.600 3.880 ;
        RECT  1.790 2.490 2.070 3.880 ;
        RECT  1.110 3.260 1.790 3.880 ;
        RECT  0.830 2.490 1.110 3.880 ;
        RECT  0.000 3.320 0.830 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 2.060 3.510 2.890 ;
        RECT  2.550 2.730 3.230 2.890 ;
        RECT  2.270 2.120 2.550 2.890 ;
        RECT  1.590 2.120 2.270 2.280 ;
        RECT  1.310 2.120 1.590 2.770 ;
        RECT  0.630 2.120 1.310 2.280 ;
        RECT  0.350 2.120 0.630 2.770 ;
    END
END AOI21X2TR

MACRO AOI21X1TR
    CLASS CORE ;
    FOREIGN AOI21X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.840 1.920 1.960 ;
        RECT  1.680 0.840 1.840 2.560 ;
        RECT  1.370 0.920 1.680 1.080 ;
        RECT  1.530 2.280 1.680 2.560 ;
        RECT  0.970 0.800 1.370 1.080 ;
        END
        ANTENNADIFFAREA 2.488 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.460 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.156 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.430 0.590 1.740 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.240 1.120 1.870 ;
        END
        ANTENNAGATEAREA 0.1728 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.280 2.000 0.280 ;
        RECT  1.530 -0.280 1.810 0.680 ;
        RECT  0.390 -0.280 1.530 0.280 ;
        RECT  0.100 -0.280 0.390 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 3.320 2.000 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 2.120 1.330 2.560 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.560 ;
    END
END AOI21X1TR

MACRO AOI211XLTR
    CLASS CORE ;
    FOREIGN AOI211XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.860 2.320 2.760 ;
        RECT  2.020 0.860 2.160 1.080 ;
        RECT  2.080 1.640 2.160 2.760 ;
        RECT  1.960 2.040 2.080 2.760 ;
        RECT  1.300 0.920 2.020 1.080 ;
        RECT  1.020 0.870 1.300 1.080 ;
        END
        ANTENNADIFFAREA 2.172 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.550 1.520 2.360 ;
        RECT  1.280 2.040 1.300 2.360 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.750 ;
        END
        ANTENNAGATEAREA 0.0936 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.640 1.770 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.330 1.120 2.360 ;
        RECT  0.480 2.040 0.880 2.360 ;
        END
        ANTENNAGATEAREA 0.1128 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.280 2.400 0.280 ;
        RECT  1.440 -0.280 1.720 0.400 ;
        RECT  0.500 -0.280 1.440 0.340 ;
        RECT  0.220 -0.280 0.500 1.080 ;
        RECT  0.000 -0.280 0.220 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 3.320 2.400 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.090 2.520 1.440 2.740 ;
    END
END AOI211XLTR

MACRO AOI211X4TR
    CLASS CORE ;
    FOREIGN AOI211X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.040 3.920 1.760 ;
        RECT  3.560 0.440 3.800 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.240 1.520 1.880 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.520 1.920 2.100 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.510 1.010 1.960 ;
        END
        ANTENNAGATEAREA 0.1248 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.280 -0.280 4.400 0.280 ;
        RECT  4.000 -0.280 4.280 0.680 ;
        RECT  3.320 -0.280 4.000 0.280 ;
        RECT  3.040 -0.280 3.320 1.310 ;
        RECT  1.720 -0.280 3.040 0.340 ;
        RECT  1.440 -0.280 1.720 0.750 ;
        RECT  0.370 -0.280 1.440 0.340 ;
        RECT  0.090 -0.280 0.370 0.450 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.280 3.320 4.400 3.880 ;
        RECT  4.000 1.950 4.280 3.880 ;
        RECT  3.320 3.320 4.000 3.880 ;
        RECT  3.040 1.910 3.320 3.880 ;
        RECT  0.850 3.320 3.040 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.880 1.470 3.400 1.750 ;
        RECT  2.800 1.150 2.880 2.070 ;
        RECT  2.720 0.570 2.800 2.930 ;
        RECT  2.520 0.570 2.720 1.310 ;
        RECT  2.520 1.910 2.720 2.930 ;
        RECT  2.360 1.470 2.560 1.750 ;
        RECT  2.200 0.910 2.360 2.550 ;
        RECT  0.920 0.910 2.200 1.080 ;
        RECT  2.130 2.390 2.200 2.550 ;
        RECT  1.850 2.390 2.130 2.720 ;
        RECT  1.050 2.120 1.330 2.720 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.720 ;
    END
END AOI211X4TR

MACRO AOI211X2TR
    CLASS CORE ;
    FOREIGN AOI211X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 0.840 3.920 1.960 ;
        RECT  3.640 0.840 3.800 2.280 ;
        RECT  3.570 0.840 3.640 1.080 ;
        RECT  3.090 2.120 3.640 2.280 ;
        RECT  3.290 0.620 3.570 1.080 ;
        RECT  2.680 0.920 3.290 1.080 ;
        RECT  2.810 2.120 3.090 2.840 ;
        RECT  1.840 0.800 2.680 1.080 ;
        RECT  0.680 0.920 1.840 1.080 ;
        RECT  0.520 0.460 0.680 1.080 ;
        RECT  0.210 0.460 0.520 0.680 ;
        END
        ANTENNADIFFAREA 8.174 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.240 3.480 1.640 ;
        RECT  2.430 1.240 3.320 1.400 ;
        RECT  2.270 1.240 2.430 1.880 ;
        RECT  2.040 1.240 2.270 1.560 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.640 3.160 1.960 ;
        END
        ANTENNAGATEAREA 0.36 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.240 1.240 1.560 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.600 1.790 1.880 ;
        RECT  0.680 1.720 1.500 1.880 ;
        RECT  0.520 1.240 0.680 1.880 ;
        RECT  0.320 1.240 0.520 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.090 -0.280 4.000 0.280 ;
        RECT  2.800 -0.280 3.090 0.670 ;
        RECT  1.330 -0.280 2.800 0.280 ;
        RECT  1.050 -0.280 1.330 0.760 ;
        RECT  0.000 -0.280 1.050 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 3.320 4.000 3.880 ;
        RECT  1.530 2.520 1.810 3.880 ;
        RECT  0.850 3.260 1.530 3.880 ;
        RECT  0.570 2.570 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.610 2.440 3.890 3.160 ;
        RECT  2.290 3.000 3.610 3.160 ;
        RECT  2.130 2.040 2.290 3.160 ;
        RECT  2.010 2.040 2.130 2.970 ;
        RECT  1.330 2.040 2.010 2.200 ;
        RECT  1.050 2.040 1.330 2.950 ;
        RECT  0.660 2.040 1.050 2.200 ;
        RECT  0.500 2.040 0.660 2.280 ;
        RECT  0.370 2.120 0.500 2.280 ;
        RECT  0.090 2.120 0.370 2.970 ;
    END
END AOI211X2TR

MACRO AOI211X1TR
    CLASS CORE ;
    FOREIGN AOI211X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.920 2.320 2.760 ;
        RECT  2.160 0.800 2.240 2.930 ;
        RECT  1.960 0.800 2.160 1.080 ;
        RECT  2.080 1.640 2.160 2.930 ;
        RECT  1.960 1.910 2.080 2.930 ;
        RECT  1.300 0.920 1.960 1.080 ;
        RECT  1.020 0.800 1.300 1.080 ;
        END
        ANTENNADIFFAREA 3.378 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.490 1.520 2.360 ;
        RECT  1.280 2.040 1.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.750 ;
        END
        ANTENNAGATEAREA 0.1776 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.640 1.770 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.330 1.120 2.360 ;
        RECT  0.480 1.980 0.880 2.360 ;
        END
        ANTENNAGATEAREA 0.1944 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.280 2.400 0.280 ;
        RECT  1.440 -0.280 1.720 0.400 ;
        RECT  0.500 -0.280 1.440 0.340 ;
        RECT  0.220 -0.280 0.500 1.030 ;
        RECT  0.000 -0.280 0.220 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 3.320 2.400 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.160 2.650 1.440 2.930 ;
        RECT  0.370 2.650 1.160 2.890 ;
        RECT  0.090 2.590 0.370 2.890 ;
    END
END AOI211X1TR

MACRO AO22XLTR
    CLASS CORE ;
    FOREIGN AO22XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.030 2.720 3.000 ;
        RECT  2.430 1.030 2.480 1.310 ;
        RECT  1.890 2.720 2.480 3.000 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.490 1.030 1.670 ;
        RECT  0.480 1.490 0.790 1.960 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.220 1.960 1.660 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 0.490 1.400 0.710 ;
        RECT  0.840 0.440 1.200 0.870 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.280 2.800 0.280 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.370 -0.280 1.860 0.280 ;
        RECT  0.090 -0.280 0.370 0.680 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 3.320 2.800 3.880 ;
        RECT  1.750 3.200 2.030 3.880 ;
        RECT  0.830 3.260 1.750 3.880 ;
        RECT  0.550 2.800 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 0.590 2.470 0.870 ;
        RECT  2.060 0.590 2.250 1.030 ;
        RECT  2.080 1.930 2.200 2.210 ;
        RECT  1.920 1.930 2.080 2.510 ;
        RECT  1.520 0.870 2.060 1.030 ;
        RECT  1.180 2.350 1.920 2.510 ;
        RECT  1.520 1.910 1.720 2.190 ;
        RECT  1.360 0.870 1.520 2.190 ;
        RECT  1.000 1.030 1.360 1.310 ;
        RECT  1.020 1.930 1.180 2.510 ;
        RECT  0.370 2.350 1.020 2.510 ;
        RECT  0.210 2.350 0.370 2.800 ;
        RECT  0.090 2.520 0.210 2.800 ;
    END
END AO22XLTR

MACRO AO22X4TR
    CLASS CORE ;
    FOREIGN AO22X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.440 3.240 2.830 ;
        RECT  2.880 1.440 2.940 2.160 ;
        RECT  2.780 1.440 2.880 1.670 ;
        RECT  2.540 0.450 2.780 1.670 ;
        RECT  2.440 0.450 2.540 1.090 ;
        END
        ANTENNADIFFAREA 3.788 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.360 0.640 1.650 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.390 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.360 1.960 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.690 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.280 4.000 0.280 ;
        RECT  2.980 -0.280 3.140 1.100 ;
        RECT  2.200 -0.280 2.980 0.280 ;
        RECT  1.920 -0.280 2.200 0.760 ;
        RECT  0.390 -0.280 1.920 0.280 ;
        RECT  0.100 -0.280 0.390 0.650 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 3.320 4.000 3.880 ;
        RECT  3.440 2.110 3.720 3.880 ;
        RECT  2.750 3.320 3.440 3.880 ;
        RECT  2.480 2.520 2.750 3.880 ;
        RECT  0.860 3.320 2.480 3.880 ;
        RECT  0.580 2.590 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 1.320 2.380 1.670 ;
        RECT  2.120 0.920 2.280 2.280 ;
        RECT  2.080 2.440 2.240 3.160 ;
        RECT  1.260 0.920 2.120 1.080 ;
        RECT  1.830 2.120 2.120 2.280 ;
        RECT  1.280 3.000 2.080 3.160 ;
        RECT  1.530 2.120 1.830 2.840 ;
        RECT  1.120 2.270 1.280 3.160 ;
        RECT  1.000 0.520 1.260 1.080 ;
        RECT  0.380 2.270 1.120 2.430 ;
        RECT  0.120 2.270 0.380 3.160 ;
    END
END AO22X4TR

MACRO AO22X2TR
    CLASS CORE ;
    FOREIGN AO22X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 0.440 2.850 1.250 ;
        RECT  2.570 0.440 2.760 3.000 ;
        RECT  2.440 2.440 2.570 3.000 ;
        RECT  2.030 2.760 2.440 3.000 ;
        END
        ANTENNADIFFAREA 3.118 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.210 0.510 1.590 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.970 1.600 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.440 1.560 0.760 ;
        END
        ANTENNAGATEAREA 0.132 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 -0.280 3.200 0.280 ;
        RECT  2.090 -0.280 2.370 0.670 ;
        RECT  0.370 -0.280 2.090 0.280 ;
        RECT  0.090 -0.280 0.370 0.390 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.800 3.320 3.200 3.880 ;
        RECT  1.520 3.200 2.800 3.880 ;
        RECT  0.770 3.260 1.520 3.880 ;
        RECT  0.490 3.200 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.130 0.920 2.410 1.580 ;
        RECT  2.130 1.910 2.250 2.190 ;
        RECT  1.480 0.920 2.130 1.080 ;
        RECT  1.970 1.910 2.130 2.510 ;
        RECT  1.290 2.350 1.970 2.510 ;
        RECT  1.490 1.910 1.770 2.190 ;
        RECT  1.480 1.910 1.490 2.070 ;
        RECT  1.320 0.920 1.480 2.070 ;
        RECT  1.010 0.920 1.320 1.080 ;
        RECT  1.010 2.230 1.290 2.510 ;
        RECT  0.370 2.230 1.010 2.390 ;
        RECT  0.090 2.230 0.370 2.510 ;
    END
END AO22X2TR

MACRO AO22X1TR
    CLASS CORE ;
    FOREIGN AO22X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.990 2.720 3.000 ;
        RECT  2.430 0.990 2.480 1.270 ;
        RECT  1.650 2.720 2.480 3.000 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.480 0.880 1.750 ;
        RECT  0.480 1.480 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.180 1.960 1.620 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.440 1.200 0.870 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 -0.280 2.800 0.280 ;
        RECT  1.790 -0.280 2.070 0.400 ;
        RECT  0.370 -0.280 1.790 0.280 ;
        RECT  0.090 -0.280 0.370 0.580 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.040 3.320 2.800 3.880 ;
        RECT  1.660 3.200 2.040 3.880 ;
        RECT  0.830 3.260 1.660 3.880 ;
        RECT  0.550 2.680 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.230 0.480 2.510 0.760 ;
        RECT  1.520 0.600 2.230 0.760 ;
        RECT  2.080 1.970 2.200 2.250 ;
        RECT  1.920 1.970 2.080 2.510 ;
        RECT  1.170 2.350 1.920 2.510 ;
        RECT  1.520 1.910 1.720 2.190 ;
        RECT  1.360 0.600 1.520 2.190 ;
        RECT  0.920 1.030 1.360 1.310 ;
        RECT  0.950 1.970 1.170 2.510 ;
        RECT  0.370 2.350 0.950 2.510 ;
        RECT  0.210 2.350 0.370 2.840 ;
        RECT  0.090 2.560 0.210 2.840 ;
    END
END AO22X1TR

MACRO AO21XLTR
    CLASS CORE ;
    FOREIGN AO21XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.030 2.320 2.760 ;
        RECT  2.040 1.030 2.080 1.560 ;
        RECT  1.930 2.600 2.080 2.760 ;
        RECT  2.030 1.030 2.040 1.310 ;
        RECT  1.650 2.600 1.930 2.880 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.200 1.520 1.640 ;
        END
        ANTENNAGATEAREA 0.06 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 2.350 1.160 2.760 ;
        END
        ANTENNAGATEAREA 0.0672 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.280 2.400 0.280 ;
        RECT  1.480 -0.280 1.760 0.400 ;
        RECT  0.390 -0.280 1.480 0.340 ;
        RECT  0.100 -0.280 0.390 1.050 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 3.320 2.400 3.880 ;
        RECT  1.510 3.200 1.790 3.880 ;
        RECT  0.830 3.260 1.510 3.880 ;
        RECT  0.550 3.200 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.590 2.070 0.870 ;
        RECT  1.680 0.590 1.840 2.190 ;
        RECT  1.270 0.590 1.680 0.800 ;
        RECT  1.080 1.910 1.360 2.190 ;
        RECT  0.990 0.520 1.270 0.800 ;
        RECT  0.430 1.970 1.080 2.190 ;
        RECT  0.160 1.910 0.430 2.190 ;
    END
END AO21XLTR

MACRO AO21X4TR
    CLASS CORE ;
    FOREIGN AO21X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.780 1.020 2.820 2.070 ;
        RECT  2.580 0.440 2.780 3.080 ;
        RECT  2.500 0.440 2.580 1.310 ;
        RECT  2.480 1.910 2.580 3.080 ;
        END
        ANTENNADIFFAREA 3.94 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.240 1.960 1.640 ;
        END
        ANTENNAGATEAREA 0.2424 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.840 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.160 1.640 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.280 3.600 0.280 ;
        RECT  2.980 -0.280 3.260 1.310 ;
        RECT  2.300 -0.280 2.980 0.280 ;
        RECT  1.580 -0.280 2.300 0.760 ;
        RECT  0.520 -0.280 1.580 0.280 ;
        RECT  0.240 -0.280 0.520 0.610 ;
        RECT  0.000 -0.280 0.240 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 3.320 3.600 3.880 ;
        RECT  2.980 1.910 3.260 3.880 ;
        RECT  2.300 3.320 2.980 3.880 ;
        RECT  2.020 2.930 2.300 3.880 ;
        RECT  1.000 3.320 2.020 3.880 ;
        RECT  0.720 2.120 1.000 3.880 ;
        RECT  0.000 3.320 0.720 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 1.470 2.420 1.750 ;
        RECT  2.120 0.920 2.280 2.070 ;
        RECT  1.340 0.920 2.120 1.080 ;
        RECT  1.990 1.910 2.120 2.070 ;
        RECT  1.680 1.910 1.990 2.750 ;
        RECT  1.200 1.800 1.480 3.160 ;
        RECT  1.060 0.590 1.340 1.080 ;
        RECT  0.520 1.800 1.200 1.960 ;
        RECT  0.240 1.800 0.520 3.100 ;
    END
END AO21X4TR

MACRO AO21X2TR
    CLASS CORE ;
    FOREIGN AO21X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 0.440 2.680 1.260 ;
        RECT  2.460 0.440 2.620 2.600 ;
        RECT  2.360 2.440 2.460 2.600 ;
        RECT  2.110 2.440 2.360 2.760 ;
        RECT  1.850 2.440 2.110 3.000 ;
        END
        ANTENNADIFFAREA 2.848 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.240 1.920 1.620 ;
        RECT  1.490 1.340 1.680 1.620 ;
        END
        ANTENNAGATEAREA 0.1224 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.330 0.810 1.610 ;
        RECT  0.440 1.240 0.720 1.610 ;
        END
        ANTENNAGATEAREA 0.1392 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.440 1.320 0.730 ;
        RECT  0.880 0.440 1.120 0.760 ;
        END
        ANTENNAGATEAREA 0.1368 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.280 2.800 0.280 ;
        RECT  1.850 -0.280 2.130 0.670 ;
        RECT  0.680 -0.280 1.850 0.280 ;
        RECT  0.400 -0.280 0.680 0.800 ;
        RECT  0.000 -0.280 0.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 3.320 2.800 3.880 ;
        RECT  1.090 3.200 2.130 3.880 ;
        RECT  0.810 2.250 1.090 3.880 ;
        RECT  0.000 3.320 0.810 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.080 0.900 2.240 2.140 ;
        RECT  1.460 0.900 2.080 1.060 ;
        RECT  1.770 1.860 2.080 2.140 ;
        RECT  1.290 1.910 1.570 2.220 ;
        RECT  1.300 0.900 1.460 1.180 ;
        RECT  0.610 1.910 1.290 2.070 ;
        RECT  0.330 1.910 0.610 2.230 ;
    END
END AO21X2TR

MACRO AO21X1TR
    CLASS CORE ;
    FOREIGN AO21X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.240 2.320 2.880 ;
        RECT  2.160 1.030 2.310 2.880 ;
        RECT  2.030 1.030 2.160 2.360 ;
        RECT  1.900 2.720 2.160 2.880 ;
        RECT  1.610 2.720 1.900 3.000 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.200 1.520 1.640 ;
        END
        ANTENNAGATEAREA 0.0648 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.240 0.760 1.640 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 2.350 1.180 2.760 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 -0.280 2.400 0.280 ;
        RECT  1.500 -0.280 1.780 0.360 ;
        RECT  0.370 -0.280 1.500 0.340 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 3.320 2.400 3.880 ;
        RECT  1.580 3.200 1.910 3.880 ;
        RECT  0.720 3.320 1.580 3.880 ;
        RECT  0.450 2.560 0.720 3.880 ;
        RECT  0.000 3.320 0.450 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.520 2.110 0.800 ;
        RECT  1.680 0.520 1.840 2.190 ;
        RECT  1.630 0.520 1.680 1.030 ;
        RECT  0.980 0.810 1.630 1.030 ;
        RECT  0.100 1.910 1.380 2.190 ;
    END
END AO21X1TR

MACRO ANTENNATR
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNATR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.870 0.570 1.030 ;
        RECT  0.080 0.440 0.320 1.560 ;
        END
        ANTENNAGATEAREA 2.449 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
END ANTENNATR

MACRO AND4XLTR
    CLASS CORE ;
    FOREIGN AND4XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.890 2.720 2.760 ;
        RECT  2.360 0.890 2.560 1.050 ;
        RECT  2.480 1.640 2.560 2.760 ;
        END
        ANTENNADIFFAREA 1.209 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.600 1.940 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.580 1.480 1.860 ;
        RECT  0.880 1.240 1.120 1.860 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.410 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.280 2.800 0.280 ;
        RECT  1.820 -0.280 2.130 1.050 ;
        RECT  0.000 -0.280 1.820 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 3.320 2.800 3.880 ;
        RECT  1.890 2.520 2.170 3.880 ;
        RECT  1.220 3.320 1.890 3.880 ;
        RECT  0.460 2.840 1.220 3.880 ;
        RECT  0.000 3.320 0.460 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 1.220 2.400 1.440 ;
        RECT  2.100 1.220 2.260 2.280 ;
        RECT  1.530 1.220 2.100 1.380 ;
        RECT  1.680 2.120 2.100 2.280 ;
        RECT  1.400 2.120 1.680 2.800 ;
        RECT  1.370 0.920 1.530 1.380 ;
        RECT  0.750 2.120 1.400 2.280 ;
        RECT  0.580 0.920 1.370 1.080 ;
        RECT  0.530 2.120 0.750 2.400 ;
        RECT  0.300 0.800 0.580 1.080 ;
    END
END AND4XLTR

MACRO AND4X8TR
    CLASS CORE ;
    FOREIGN AND4X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.910 0.650 6.220 3.160 ;
        RECT  5.900 1.030 5.910 3.160 ;
        RECT  5.270 1.030 5.900 1.760 ;
        RECT  5.200 0.440 5.270 1.760 ;
        RECT  5.040 0.440 5.200 3.160 ;
        END
        ANTENNADIFFAREA 7.776 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.240 4.560 2.680 ;
        RECT  4.300 1.240 4.400 1.520 ;
        RECT  1.920 2.520 4.400 2.680 ;
        RECT  1.600 1.900 1.920 2.680 ;
        END
        ANTENNAGATEAREA 0.5184 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.020 1.920 4.240 2.360 ;
        RECT  2.320 2.200 4.020 2.360 ;
        RECT  2.080 1.580 2.320 2.360 ;
        RECT  1.240 1.580 2.080 1.740 ;
        RECT  1.020 1.580 1.240 1.860 ;
        END
        ANTENNAGATEAREA 0.5184 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.540 1.580 3.820 1.860 ;
        RECT  2.760 1.700 3.540 1.860 ;
        RECT  2.600 1.240 2.760 1.860 ;
        RECT  0.800 1.240 2.600 1.400 ;
        RECT  0.500 1.240 0.800 1.960 ;
        RECT  0.480 1.640 0.500 1.960 ;
        END
        ANTENNAGATEAREA 0.5184 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 0.920 3.290 1.540 ;
        RECT  0.320 0.920 3.120 1.080 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.5184 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.710 -0.280 6.800 0.280 ;
        RECT  6.430 -0.280 6.710 1.310 ;
        RECT  5.750 -0.280 6.430 0.340 ;
        RECT  5.470 -0.280 5.750 0.870 ;
        RECT  4.790 -0.280 5.470 0.280 ;
        RECT  4.500 -0.280 4.790 0.670 ;
        RECT  1.860 -0.280 4.500 0.280 ;
        RECT  1.580 -0.280 1.860 0.400 ;
        RECT  0.000 -0.280 1.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.700 3.320 6.800 3.880 ;
        RECT  6.420 1.910 6.700 3.880 ;
        RECT  5.740 3.320 6.420 3.880 ;
        RECT  5.460 2.010 5.740 3.880 ;
        RECT  4.700 3.320 5.460 3.880 ;
        RECT  4.420 3.200 4.700 3.880 ;
        RECT  3.660 3.320 4.420 3.880 ;
        RECT  3.380 3.200 3.660 3.880 ;
        RECT  2.620 3.320 3.380 3.880 ;
        RECT  2.340 3.200 2.620 3.880 ;
        RECT  1.580 3.320 2.340 3.880 ;
        RECT  1.300 3.200 1.580 3.880 ;
        RECT  0.580 3.260 1.300 3.880 ;
        RECT  0.300 2.530 0.580 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.720 0.830 4.880 3.000 ;
        RECT  4.030 0.830 4.720 0.990 ;
        RECT  4.180 2.840 4.720 3.000 ;
        RECT  3.900 2.840 4.180 3.120 ;
        RECT  3.870 0.600 4.030 0.990 ;
        RECT  3.140 2.840 3.900 3.000 ;
        RECT  3.380 0.600 3.870 0.760 ;
        RECT  3.040 0.480 3.380 0.760 ;
        RECT  2.860 2.840 3.140 3.120 ;
        RECT  0.650 0.600 3.040 0.760 ;
        RECT  2.100 2.840 2.860 3.000 ;
        RECT  1.820 2.840 2.100 3.120 ;
        RECT  1.060 2.840 1.820 3.000 ;
        RECT  0.900 2.330 1.060 3.000 ;
        RECT  0.780 2.330 0.900 2.950 ;
        RECT  0.490 0.440 0.650 0.760 ;
        RECT  0.100 0.440 0.490 0.680 ;
    END
END AND4X8TR

MACRO AND4X6TR
    CLASS CORE ;
    FOREIGN AND4X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.160 0.770 5.440 3.160 ;
        RECT  4.480 1.040 5.160 1.910 ;
        RECT  4.300 0.530 4.480 3.160 ;
        RECT  4.200 0.530 4.300 1.310 ;
        RECT  4.200 1.910 4.300 3.160 ;
        END
        ANTENNADIFFAREA 7.064 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.770 3.720 2.050 ;
        RECT  3.440 1.770 3.600 2.370 ;
        RECT  0.610 2.210 3.440 2.370 ;
        RECT  0.320 1.450 0.610 2.370 ;
        RECT  0.080 1.240 0.320 2.370 ;
        END
        ANTENNAGATEAREA 0.4008 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.640 3.280 1.980 ;
        RECT  2.880 0.920 3.040 1.980 ;
        RECT  1.090 0.920 2.880 1.080 ;
        RECT  0.930 0.920 1.090 2.050 ;
        RECT  0.810 1.770 0.930 2.050 ;
        END
        ANTENNAGATEAREA 0.4008 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.240 2.720 2.000 ;
        RECT  1.530 1.800 2.480 1.960 ;
        RECT  1.250 1.770 1.530 2.050 ;
        END
        ANTENNAGATEAREA 0.4008 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 2.090 1.640 ;
        END
        ANTENNAGATEAREA 0.4008 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.960 -0.280 5.600 0.280 ;
        RECT  4.680 -0.280 4.960 0.870 ;
        RECT  4.000 -0.280 4.680 0.280 ;
        RECT  3.720 -0.280 4.000 1.200 ;
        RECT  0.610 -0.280 3.720 0.280 ;
        RECT  0.330 -0.280 0.610 1.080 ;
        RECT  0.000 -0.280 0.330 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.960 3.320 5.600 3.880 ;
        RECT  4.680 2.230 4.960 3.880 ;
        RECT  3.960 3.320 4.680 3.880 ;
        RECT  3.680 3.200 3.960 3.880 ;
        RECT  3.050 3.320 3.680 3.880 ;
        RECT  2.770 3.200 3.050 3.880 ;
        RECT  2.130 3.320 2.770 3.880 ;
        RECT  1.850 3.200 2.130 3.880 ;
        RECT  1.330 3.320 1.850 3.880 ;
        RECT  1.050 3.200 1.330 3.880 ;
        RECT  0.370 3.260 1.050 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.040 1.470 4.140 1.750 ;
        RECT  3.880 1.360 4.040 2.690 ;
        RECT  3.560 1.360 3.880 1.520 ;
        RECT  3.570 2.530 3.880 2.690 ;
        RECT  3.290 2.530 3.570 2.810 ;
        RECT  3.400 0.600 3.560 1.520 ;
        RECT  2.330 0.600 3.400 0.760 ;
        RECT  2.650 2.530 3.290 2.690 ;
        RECT  2.370 2.530 2.650 2.810 ;
        RECT  1.730 2.530 2.370 2.690 ;
        RECT  1.770 0.480 2.330 0.760 ;
        RECT  1.450 2.530 1.730 2.810 ;
        RECT  0.810 2.530 1.450 2.690 ;
        RECT  0.530 2.530 0.810 2.810 ;
    END
END AND4X6TR

MACRO AND4X4TR
    CLASS CORE ;
    FOREIGN AND4X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.040 4.320 2.150 ;
        RECT  4.040 1.040 4.080 1.310 ;
        RECT  4.040 1.910 4.080 2.150 ;
        RECT  3.760 0.440 4.040 1.310 ;
        RECT  3.760 1.910 4.040 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.420 3.280 2.430 ;
        RECT  3.000 1.420 3.120 1.700 ;
        RECT  2.510 2.270 3.120 2.430 ;
        RECT  2.350 2.270 2.510 2.680 ;
        RECT  0.720 2.520 2.350 2.680 ;
        RECT  0.560 1.360 0.720 2.680 ;
        RECT  0.440 1.360 0.560 1.960 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.820 2.880 2.100 ;
        RECT  2.600 1.640 2.760 2.100 ;
        RECT  2.440 1.150 2.600 2.100 ;
        RECT  1.120 1.150 2.440 1.310 ;
        RECT  0.960 1.150 1.120 1.980 ;
        RECT  0.900 1.700 0.960 1.980 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.820 2.280 2.100 ;
        RECT  1.960 1.940 2.000 2.100 ;
        RECT  1.680 1.940 1.960 2.360 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.470 1.760 1.750 ;
        RECT  1.480 1.470 1.520 1.960 ;
        RECT  1.280 1.590 1.480 1.960 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.560 -0.280 4.800 0.280 ;
        RECT  4.280 -0.280 4.560 0.770 ;
        RECT  3.520 -0.280 4.280 0.280 ;
        RECT  3.190 -0.280 3.520 0.870 ;
        RECT  0.510 -0.280 3.190 0.340 ;
        RECT  0.240 -0.280 0.510 1.070 ;
        RECT  0.000 -0.280 0.240 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 3.320 4.800 3.880 ;
        RECT  4.240 2.330 4.520 3.880 ;
        RECT  3.560 3.320 4.240 3.880 ;
        RECT  3.280 2.910 3.560 3.880 ;
        RECT  2.520 3.320 3.280 3.880 ;
        RECT  2.240 3.200 2.520 3.880 ;
        RECT  1.440 3.320 2.240 3.880 ;
        RECT  1.160 2.840 1.440 3.880 ;
        RECT  0.000 3.320 1.160 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.600 1.470 3.780 1.750 ;
        RECT  3.440 1.100 3.600 2.750 ;
        RECT  2.920 1.100 3.440 1.260 ;
        RECT  3.080 2.590 3.440 2.750 ;
        RECT  2.800 2.590 3.080 3.000 ;
        RECT  2.760 0.710 2.920 1.260 ;
        RECT  2.000 2.840 2.800 3.000 ;
        RECT  1.680 0.710 2.760 0.990 ;
        RECT  1.720 2.840 2.000 3.120 ;
    END
END AND4X4TR

MACRO AND4X2TR
    CLASS CORE ;
    FOREIGN AND4X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.500 3.120 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.640 2.360 1.960 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.960 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.680 1.300 1.960 ;
        RECT  0.960 1.240 1.120 1.960 ;
        RECT  0.880 1.240 0.960 1.560 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.630 0.680 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1344 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.500 -0.280 3.200 0.280 ;
        RECT  2.220 -0.280 2.500 0.680 ;
        RECT  0.000 -0.280 2.220 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 3.320 3.200 3.880 ;
        RECT  2.300 2.440 2.580 3.880 ;
        RECT  1.540 3.260 2.300 3.880 ;
        RECT  1.260 2.440 1.540 3.880 ;
        RECT  0.540 3.260 1.260 3.880 ;
        RECT  0.260 2.230 0.540 3.880 ;
        RECT  0.000 3.320 0.260 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.520 0.920 2.680 2.280 ;
        RECT  0.880 0.920 2.520 1.080 ;
        RECT  2.060 2.120 2.520 2.280 ;
        RECT  1.780 2.120 2.060 2.400 ;
        RECT  1.020 2.120 1.780 2.280 ;
        RECT  0.740 2.120 1.020 2.400 ;
        RECT  0.600 0.800 0.880 1.080 ;
    END
END AND4X2TR

MACRO AND4X1TR
    CLASS CORE ;
    FOREIGN AND4X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.650 2.720 2.760 ;
        RECT  2.410 0.650 2.560 0.930 ;
        RECT  2.480 1.640 2.560 2.760 ;
        END
        ANTENNADIFFAREA 1.792 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.600 1.940 1.960 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.580 1.480 1.860 ;
        RECT  0.880 1.240 1.120 1.860 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.410 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.072 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.210 -0.280 2.800 0.280 ;
        RECT  1.930 -0.280 2.210 0.930 ;
        RECT  0.000 -0.280 1.930 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 3.320 2.800 3.880 ;
        RECT  1.890 2.520 2.170 3.880 ;
        RECT  1.220 3.320 1.890 3.880 ;
        RECT  0.480 2.840 1.220 3.880 ;
        RECT  0.000 3.320 0.480 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 1.160 2.400 1.440 ;
        RECT  2.100 1.160 2.260 2.280 ;
        RECT  1.770 1.160 2.100 1.320 ;
        RECT  1.680 2.120 2.100 2.280 ;
        RECT  1.610 0.920 1.770 1.320 ;
        RECT  1.400 2.120 1.680 2.800 ;
        RECT  0.780 0.920 1.610 1.080 ;
        RECT  0.750 2.120 1.400 2.280 ;
        RECT  0.330 0.800 0.780 1.080 ;
        RECT  0.530 2.120 0.750 2.400 ;
    END
END AND4X1TR

MACRO AND3XLTR
    CLASS CORE ;
    FOREIGN AND3XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.090 2.320 2.760 ;
        RECT  2.000 1.090 2.160 1.250 ;
        RECT  2.080 1.640 2.160 2.760 ;
        RECT  2.030 2.010 2.080 2.760 ;
        END
        ANTENNADIFFAREA 1.2875 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.240 1.520 1.750 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.440 1.120 0.760 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.280 2.400 0.280 ;
        RECT  1.320 -0.280 1.630 0.760 ;
        RECT  0.000 -0.280 1.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 3.320 2.400 3.880 ;
        RECT  1.480 2.260 1.760 3.880 ;
        RECT  0.830 3.320 1.480 3.880 ;
        RECT  0.550 2.500 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.440 1.900 1.690 ;
        RECT  1.680 0.920 1.840 2.090 ;
        RECT  0.400 0.920 1.680 1.080 ;
        RECT  1.180 1.910 1.680 2.090 ;
        RECT  1.020 1.910 1.180 2.280 ;
        RECT  0.370 2.120 1.020 2.280 ;
        RECT  0.120 0.920 0.400 1.290 ;
        RECT  0.210 2.120 0.370 2.780 ;
        RECT  0.090 2.500 0.210 2.780 ;
    END
END AND3XLTR

MACRO AND3X8TR
    CLASS CORE ;
    FOREIGN AND3X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.610 1.650 4.690 3.160 ;
        RECT  4.410 0.440 4.610 3.160 ;
        RECT  4.330 0.440 4.410 1.760 ;
        RECT  3.730 1.040 4.330 1.760 ;
        RECT  3.490 1.040 3.730 3.160 ;
        RECT  3.450 0.440 3.490 3.160 ;
        RECT  3.210 0.440 3.450 1.250 ;
        END
        ANTENNADIFFAREA 7.488 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.850 2.970 2.130 ;
        RECT  2.690 1.850 2.850 2.440 ;
        RECT  0.720 2.280 2.690 2.440 ;
        RECT  0.570 1.860 0.720 2.440 ;
        RECT  0.560 1.740 0.570 2.440 ;
        RECT  0.480 1.740 0.560 2.360 ;
        RECT  0.290 1.740 0.480 2.020 ;
        END
        ANTENNAGATEAREA 0.468 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.840 2.490 2.120 ;
        RECT  1.160 1.960 2.210 2.120 ;
        RECT  0.880 1.640 1.160 2.120 ;
        END
        ANTENNAGATEAREA 0.468 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 2.010 1.780 ;
        RECT  1.330 1.500 1.640 1.780 ;
        END
        ANTENNAGATEAREA 0.468 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.280 6.000 0.280 ;
        RECT  4.850 -0.280 5.130 1.310 ;
        RECT  4.050 -0.280 4.850 0.280 ;
        RECT  3.770 -0.280 4.050 0.670 ;
        RECT  3.010 -0.280 3.770 0.280 ;
        RECT  2.730 -0.280 3.010 1.250 ;
        RECT  0.690 -0.280 2.730 0.280 ;
        RECT  0.410 -0.280 0.690 1.110 ;
        RECT  0.000 -0.280 0.410 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.210 3.320 6.000 3.880 ;
        RECT  4.930 2.050 5.210 3.880 ;
        RECT  4.210 3.320 4.930 3.880 ;
        RECT  3.930 2.050 4.210 3.880 ;
        RECT  3.250 3.320 3.930 3.880 ;
        RECT  2.970 2.930 3.250 3.880 ;
        RECT  2.290 3.320 2.970 3.880 ;
        RECT  2.010 2.930 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.930 1.330 3.880 ;
        RECT  0.310 3.320 1.050 3.880 ;
        RECT  0.090 2.420 0.310 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 1.410 3.290 2.760 ;
        RECT  3.010 1.410 3.130 1.690 ;
        RECT  2.770 2.600 3.130 2.760 ;
        RECT  2.330 1.410 3.010 1.570 ;
        RECT  2.490 2.600 2.770 2.880 ;
        RECT  1.810 2.600 2.490 2.760 ;
        RECT  2.170 0.920 2.330 1.570 ;
        RECT  1.810 0.920 2.170 1.080 ;
        RECT  1.530 0.520 1.810 1.080 ;
        RECT  1.530 2.600 1.810 2.880 ;
        RECT  0.850 2.600 1.530 2.760 ;
        RECT  0.570 2.600 0.850 2.880 ;
    END
END AND3X8TR

MACRO AND3X6TR
    CLASS CORE ;
    FOREIGN AND3X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.340 0.500 4.620 3.160 ;
        RECT  3.700 1.440 4.340 2.160 ;
        RECT  3.660 0.440 3.700 2.160 ;
        RECT  3.430 0.440 3.660 3.160 ;
        RECT  3.380 0.440 3.430 1.310 ;
        RECT  3.380 1.910 3.430 3.160 ;
        END
        ANTENNADIFFAREA 7.48 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.150 2.900 1.630 ;
        RECT  2.240 1.150 2.620 1.310 ;
        RECT  2.080 0.920 2.240 1.310 ;
        RECT  1.180 0.920 2.080 1.080 ;
        RECT  1.020 0.920 1.180 1.400 ;
        RECT  0.760 1.240 1.020 1.400 ;
        RECT  0.440 1.240 0.760 1.560 ;
        RECT  0.400 1.240 0.440 1.540 ;
        END
        ANTENNAGATEAREA 0.3648 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.680 2.460 1.960 ;
        RECT  2.080 1.640 2.360 1.960 ;
        RECT  2.040 1.720 2.080 1.960 ;
        RECT  1.200 1.720 2.040 1.880 ;
        RECT  0.920 1.580 1.200 1.880 ;
        END
        ANTENNAGATEAREA 0.3648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.240 1.920 1.560 ;
        END
        ANTENNAGATEAREA 0.3648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 -0.280 4.800 0.280 ;
        RECT  3.860 -0.280 4.140 1.190 ;
        RECT  3.100 -0.280 3.860 0.280 ;
        RECT  2.820 -0.280 3.100 0.670 ;
        RECT  0.860 -0.280 2.820 0.280 ;
        RECT  0.580 -0.280 0.860 1.080 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 3.320 4.800 3.880 ;
        RECT  3.860 2.560 4.140 3.880 ;
        RECT  3.140 3.320 3.860 3.880 ;
        RECT  2.860 3.200 3.140 3.880 ;
        RECT  2.200 3.320 2.860 3.880 ;
        RECT  1.920 3.200 2.200 3.880 ;
        RECT  1.280 3.320 1.920 3.880 ;
        RECT  1.000 3.200 1.280 3.880 ;
        RECT  0.400 3.310 1.000 3.880 ;
        RECT  0.120 2.170 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.220 1.470 3.270 1.750 ;
        RECT  3.060 0.830 3.220 2.330 ;
        RECT  2.560 0.830 3.060 0.990 ;
        RECT  2.720 2.170 3.060 2.330 ;
        RECT  2.440 2.170 2.720 2.890 ;
        RECT  2.400 0.600 2.560 0.990 ;
        RECT  1.800 2.170 2.440 2.330 ;
        RECT  1.980 0.600 2.400 0.760 ;
        RECT  1.700 0.480 1.980 0.760 ;
        RECT  1.520 2.170 1.800 2.890 ;
        RECT  0.880 2.170 1.520 2.330 ;
        RECT  0.600 2.170 0.880 2.890 ;
    END
END AND3X6TR

MACRO AND3X4TR
    CLASS CORE ;
    FOREIGN AND3X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.040 2.730 1.760 ;
        RECT  2.280 1.040 2.360 3.160 ;
        RECT  2.110 0.600 2.280 3.160 ;
        RECT  2.040 0.600 2.110 1.280 ;
        RECT  2.080 2.020 2.110 3.160 ;
        RECT  1.920 0.600 2.040 0.760 ;
        END
        ANTENNADIFFAREA 3.897 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.560 1.750 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.520 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.240 0.720 1.670 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.280 3.200 0.280 ;
        RECT  2.440 -0.280 2.710 0.820 ;
        RECT  1.720 -0.280 2.440 0.280 ;
        RECT  1.440 -0.280 1.720 0.650 ;
        RECT  0.000 -0.280 1.440 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.920 3.320 3.200 3.880 ;
        RECT  2.640 2.020 2.920 3.880 ;
        RECT  1.880 3.320 2.640 3.880 ;
        RECT  1.600 2.440 1.880 3.880 ;
        RECT  0.920 3.320 1.600 3.880 ;
        RECT  0.640 2.440 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.880 1.490 1.940 1.770 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  0.520 0.920 1.720 1.080 ;
        RECT  1.400 2.120 1.720 2.280 ;
        RECT  1.120 2.120 1.400 2.950 ;
        RECT  0.440 2.120 1.120 2.280 ;
        RECT  0.240 0.740 0.520 1.080 ;
        RECT  0.160 2.120 0.440 2.950 ;
    END
END AND3X4TR

MACRO AND3X2TR
    CLASS CORE ;
    FOREIGN AND3X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.500 2.320 3.160 ;
        RECT  2.000 0.500 2.160 1.310 ;
        RECT  2.080 1.640 2.160 3.160 ;
        RECT  2.000 1.910 2.080 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.480 1.520 1.960 ;
        RECT  1.280 1.640 1.300 1.960 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.580 1.120 2.410 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.580 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1296 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.280 2.400 0.280 ;
        RECT  1.480 -0.280 1.760 0.800 ;
        RECT  0.000 -0.280 1.480 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 3.320 2.400 3.880 ;
        RECT  1.480 3.260 1.760 3.880 ;
        RECT  0.890 3.320 1.480 3.880 ;
        RECT  0.580 3.040 0.890 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.470 1.920 1.750 ;
        RECT  1.680 1.130 1.840 2.880 ;
        RECT  0.520 1.130 1.680 1.290 ;
        RECT  1.340 2.720 1.680 2.880 ;
        RECT  1.060 2.720 1.340 3.000 ;
        RECT  0.550 2.720 1.060 2.880 ;
        RECT  0.390 2.190 0.550 2.880 ;
        RECT  0.240 1.010 0.520 1.290 ;
        RECT  0.200 2.190 0.390 2.350 ;
    END
END AND3X2TR

MACRO AND3X1TR
    CLASS CORE ;
    FOREIGN AND3X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.920 2.320 2.760 ;
        RECT  2.000 0.920 2.160 1.200 ;
        RECT  2.080 1.640 2.160 2.760 ;
        RECT  2.030 2.070 2.080 2.760 ;
        END
        ANTENNADIFFAREA 2.036 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.520 1.750 ;
        RECT  1.200 1.450 1.280 1.750 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.830 1.120 1.230 ;
        RECT  0.760 0.830 1.040 1.480 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.640 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.0696 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.890 -0.280 2.400 0.280 ;
        RECT  1.600 -0.280 1.890 0.340 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 3.320 2.400 3.880 ;
        RECT  1.520 2.260 1.810 3.880 ;
        RECT  0.830 3.320 1.520 3.880 ;
        RECT  0.550 2.500 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 1.440 1.900 1.760 ;
        RECT  1.680 0.850 1.840 2.090 ;
        RECT  1.440 0.850 1.680 1.010 ;
        RECT  1.180 1.910 1.680 2.090 ;
        RECT  1.280 0.440 1.440 1.010 ;
        RECT  0.440 0.440 1.280 0.600 ;
        RECT  1.020 1.910 1.180 2.280 ;
        RECT  0.370 2.120 1.020 2.280 ;
        RECT  0.160 0.440 0.440 1.210 ;
        RECT  0.210 2.120 0.370 2.780 ;
        RECT  0.090 2.500 0.210 2.780 ;
    END
END AND3X1TR

MACRO AND2XLTR
    CLASS CORE ;
    FOREIGN AND2XLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.840 1.920 2.440 ;
        RECT  1.600 0.840 1.680 1.130 ;
        RECT  1.600 2.120 1.680 2.440 ;
        END
        ANTENNADIFFAREA 1.174 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.240 1.120 1.690 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.610 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.280 2.000 0.280 ;
        RECT  1.020 -0.280 1.290 0.760 ;
        RECT  0.000 -0.280 1.020 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 2.000 3.880 ;
        RECT  1.120 2.200 1.400 3.880 ;
        RECT  0.380 3.320 1.120 3.880 ;
        RECT  0.100 2.120 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.360 1.520 1.640 ;
        RECT  1.280 0.920 1.440 2.030 ;
        RECT  0.670 0.920 1.280 1.080 ;
        RECT  0.860 1.870 1.280 2.030 ;
        RECT  0.580 1.870 0.860 2.300 ;
        RECT  0.510 0.520 0.670 1.080 ;
        RECT  0.090 0.520 0.510 0.680 ;
    END
END AND2XLTR

MACRO AND2X8TR
    CLASS CORE ;
    FOREIGN AND2X8TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.040 3.730 1.760 ;
        RECT  3.410 0.580 3.690 3.160 ;
        RECT  2.730 0.980 3.410 1.760 ;
        RECT  2.450 0.980 2.730 3.160 ;
        END
        ANTENNADIFFAREA 7.712 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.580 1.850 1.860 ;
        RECT  1.570 1.580 1.730 1.960 ;
        RECT  0.640 1.800 1.570 1.960 ;
        RECT  0.320 1.420 0.640 1.960 ;
        RECT  0.080 1.420 0.320 2.760 ;
        END
        ANTENNAGATEAREA 0.4536 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.200 1.160 1.640 ;
        END
        ANTENNAGATEAREA 0.4536 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 -0.280 4.400 0.280 ;
        RECT  3.890 -0.280 4.170 1.310 ;
        RECT  3.210 -0.280 3.890 0.280 ;
        RECT  2.930 -0.280 3.210 0.670 ;
        RECT  2.050 -0.280 2.930 0.340 ;
        RECT  1.770 -0.280 2.050 0.930 ;
        RECT  0.450 -0.280 1.770 0.280 ;
        RECT  0.170 -0.280 0.450 1.080 ;
        RECT  0.000 -0.280 0.170 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 3.320 4.400 3.880 ;
        RECT  3.890 1.910 4.170 3.880 ;
        RECT  3.210 3.320 3.890 3.880 ;
        RECT  2.930 2.120 3.210 3.880 ;
        RECT  2.250 3.320 2.930 3.880 ;
        RECT  1.970 2.440 2.250 3.880 ;
        RECT  1.250 3.260 1.970 3.880 ;
        RECT  0.970 2.600 1.250 3.880 ;
        RECT  0.370 3.260 0.970 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.170 1.360 2.290 1.640 ;
        RECT  2.010 1.090 2.170 2.280 ;
        RECT  1.480 1.090 2.010 1.250 ;
        RECT  1.730 2.120 2.010 2.280 ;
        RECT  1.450 2.120 1.730 2.880 ;
        RECT  1.320 0.880 1.480 1.250 ;
        RECT  0.770 2.120 1.450 2.280 ;
        RECT  1.250 0.880 1.320 1.040 ;
        RECT  0.970 0.760 1.250 1.040 ;
        RECT  0.490 2.120 0.770 2.880 ;
    END
END AND2X8TR

MACRO AND2X6TR
    CLASS CORE ;
    FOREIGN AND2X6TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.440 3.730 3.160 ;
        RECT  2.770 1.040 3.450 1.760 ;
        RECT  2.690 1.040 2.770 3.160 ;
        RECT  2.510 0.440 2.690 3.160 ;
        RECT  2.410 0.440 2.510 1.310 ;
        RECT  2.490 1.910 2.510 3.160 ;
        END
        ANTENNADIFFAREA 7.48 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.640 1.930 1.960 ;
        RECT  0.720 1.800 1.650 1.960 ;
        RECT  0.470 1.320 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.310 1.470 1.640 ;
        RECT  0.880 1.240 1.130 1.640 ;
        END
        ANTENNAGATEAREA 0.3408 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.210 -0.280 4.000 0.280 ;
        RECT  2.930 -0.280 3.210 0.800 ;
        RECT  2.170 -0.280 2.930 0.280 ;
        RECT  1.890 -0.280 2.170 0.800 ;
        RECT  0.520 -0.280 1.890 0.280 ;
        RECT  0.240 -0.280 0.520 1.050 ;
        RECT  0.000 -0.280 0.240 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.250 3.320 4.000 3.880 ;
        RECT  2.970 2.080 3.250 3.880 ;
        RECT  2.290 3.320 2.970 3.880 ;
        RECT  2.010 2.450 2.290 3.880 ;
        RECT  1.330 3.320 2.010 3.880 ;
        RECT  1.050 2.450 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.120 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 1.470 2.350 1.750 ;
        RECT  2.090 0.960 2.250 2.280 ;
        RECT  1.730 0.960 2.090 1.120 ;
        RECT  1.810 2.120 2.090 2.280 ;
        RECT  1.530 2.120 1.810 2.730 ;
        RECT  1.570 0.920 1.730 1.120 ;
        RECT  1.350 0.920 1.570 1.080 ;
        RECT  0.850 2.120 1.530 2.280 ;
        RECT  1.040 0.800 1.350 1.080 ;
        RECT  0.570 2.120 0.850 2.730 ;
    END
END AND2X6TR

MACRO AND2X4TR
    CLASS CORE ;
    FOREIGN AND2X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.440 2.320 2.160 ;
        RECT  1.950 1.440 2.120 3.160 ;
        RECT  1.840 0.960 1.950 3.160 ;
        RECT  1.790 0.960 1.840 1.610 ;
        RECT  1.710 0.440 1.790 1.610 ;
        RECT  1.510 0.440 1.710 1.120 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.600 1.170 1.960 ;
        END
        ANTENNAGATEAREA 0.2256 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.600 0.620 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2256 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.280 2.800 0.280 ;
        RECT  2.120 -0.280 2.400 1.260 ;
        RECT  1.310 -0.280 2.120 0.280 ;
        RECT  1.030 -0.280 1.310 1.120 ;
        RECT  0.000 -0.280 1.030 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.640 3.320 2.800 3.880 ;
        RECT  2.360 2.440 2.640 3.880 ;
        RECT  1.640 3.320 2.360 3.880 ;
        RECT  1.360 2.440 1.640 3.880 ;
        RECT  0.510 3.260 1.360 3.880 ;
        RECT  0.230 2.590 0.510 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.380 1.280 1.540 2.280 ;
        RECT  0.680 1.280 1.380 1.440 ;
        RECT  0.990 2.120 1.380 2.280 ;
        RECT  0.710 2.120 0.990 2.890 ;
        RECT  0.520 0.900 0.680 1.440 ;
        RECT  0.220 0.520 0.520 1.080 ;
    END
END AND2X4TR

MACRO AND2X2TR
    CLASS CORE ;
    FOREIGN AND2X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.500 1.920 3.160 ;
        RECT  1.600 0.500 1.760 1.310 ;
        RECT  1.680 1.640 1.760 3.160 ;
        RECT  1.600 1.910 1.680 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
        ANTENNAGATEAREA 0.1176 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.380 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.1176 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 -0.280 2.000 0.280 ;
        RECT  1.110 -0.280 1.410 0.760 ;
        RECT  0.000 -0.280 1.110 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 2.000 3.880 ;
        RECT  1.120 2.560 1.400 3.880 ;
        RECT  0.390 3.290 1.120 3.880 ;
        RECT  0.130 2.160 0.390 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.470 1.520 1.750 ;
        RECT  1.280 0.920 1.440 2.340 ;
        RECT  0.430 0.920 1.280 1.080 ;
        RECT  0.830 2.180 1.280 2.340 ;
        RECT  0.670 2.180 0.830 3.000 ;
        RECT  0.550 2.720 0.670 3.000 ;
        RECT  0.150 0.920 0.430 1.220 ;
    END
END AND2X2TR

MACRO AND2X1TR
    CLASS CORE ;
    FOREIGN AND2X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.840 1.920 2.420 ;
        RECT  1.600 0.840 1.680 1.130 ;
        RECT  1.600 2.050 1.680 2.420 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.240 1.120 1.840 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.610 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.0624 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.280 2.000 0.280 ;
        RECT  1.020 -0.280 1.290 0.760 ;
        RECT  0.000 -0.280 1.020 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.320 2.000 3.880 ;
        RECT  1.120 2.320 1.400 3.880 ;
        RECT  0.380 3.320 1.120 3.880 ;
        RECT  0.100 2.120 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 1.360 1.520 1.640 ;
        RECT  1.280 0.920 1.440 2.160 ;
        RECT  0.670 0.920 1.280 1.080 ;
        RECT  0.860 2.000 1.280 2.160 ;
        RECT  0.580 2.000 0.860 2.300 ;
        RECT  0.510 0.520 0.670 1.080 ;
        RECT  0.090 0.520 0.510 0.680 ;
    END
END AND2X1TR

MACRO AHHCONX4TR
    CLASS CORE ;
    FOREIGN AHHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 2.560 3.730 2.840 ;
        RECT  2.770 2.680 3.550 2.840 ;
        RECT  2.720 2.240 2.770 2.840 ;
        RECT  2.640 1.160 2.720 2.840 ;
        RECT  2.450 0.980 2.640 2.840 ;
        RECT  2.380 0.980 2.450 2.250 ;
        RECT  1.860 1.970 2.380 2.250 ;
        RECT  1.590 1.970 1.860 2.520 ;
        END
        ANTENNADIFFAREA 5.646 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.520 1.150 6.760 2.360 ;
        RECT  6.280 1.150 6.520 1.310 ;
        RECT  6.160 2.120 6.520 2.360 ;
        RECT  6.040 0.710 6.280 1.310 ;
        RECT  5.880 2.120 6.160 3.160 ;
        RECT  4.440 0.710 6.040 0.990 ;
        RECT  5.240 2.120 5.880 2.360 ;
        RECT  4.880 2.120 5.240 3.160 ;
        END
        ANTENNADIFFAREA 6.624 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 1.470 6.360 1.960 ;
        RECT  6.040 1.640 6.080 1.960 ;
        RECT  4.920 1.800 6.040 1.960 ;
        RECT  4.620 1.470 4.920 1.960 ;
        RECT  4.460 1.470 4.620 2.700 ;
        RECT  4.110 2.540 4.460 2.700 ;
        RECT  3.950 2.540 4.110 3.160 ;
        RECT  1.050 3.000 3.950 3.160 ;
        END
        ANTENNAGATEAREA 0.936 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.240 1.360 5.480 1.640 ;
        RECT  5.080 1.150 5.240 1.640 ;
        RECT  4.120 1.150 5.080 1.310 ;
        RECT  3.840 1.150 4.120 1.850 ;
        RECT  3.640 1.150 3.840 1.560 ;
        END
        ANTENNAGATEAREA 0.8328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.080 -0.280 7.200 0.280 ;
        RECT  6.800 -0.280 7.080 0.990 ;
        RECT  5.440 -0.280 6.800 0.280 ;
        RECT  5.160 -0.280 5.440 0.400 ;
        RECT  3.790 -0.280 5.160 0.340 ;
        RECT  3.420 -0.280 3.790 0.990 ;
        RECT  0.610 -0.280 3.420 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.640 3.320 7.200 3.880 ;
        RECT  6.360 2.590 6.640 3.880 ;
        RECT  5.680 3.320 6.360 3.880 ;
        RECT  5.400 2.590 5.680 3.880 ;
        RECT  4.720 3.320 5.400 3.880 ;
        RECT  4.440 2.930 4.720 3.880 ;
        RECT  0.890 3.320 4.440 3.880 ;
        RECT  0.610 3.180 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.960 2.100 4.240 2.380 ;
        RECT  3.320 2.220 3.960 2.380 ;
        RECT  3.100 2.220 3.320 2.520 ;
        RECT  2.930 0.660 3.100 2.520 ;
        RECT  2.800 0.660 2.930 0.990 ;
        RECT  2.220 0.660 2.800 0.820 ;
        RECT  2.110 2.560 2.290 2.840 ;
        RECT  2.060 0.660 2.220 1.370 ;
        RECT  1.390 1.530 2.220 1.810 ;
        RECT  0.370 2.680 2.110 2.840 ;
        RECT  1.070 1.210 2.060 1.370 ;
        RECT  1.680 0.500 1.900 1.050 ;
        RECT  0.370 0.500 1.680 0.660 ;
        RECT  1.230 1.530 1.390 2.520 ;
        RECT  0.690 0.830 1.290 1.050 ;
        RECT  1.090 1.960 1.230 2.520 ;
        RECT  0.690 1.960 1.090 2.120 ;
        RECT  0.850 1.210 1.070 1.800 ;
        RECT  0.530 0.830 0.690 2.120 ;
        RECT  0.090 0.500 0.370 3.160 ;
    END
END AHHCONX4TR

MACRO AHHCONX2TR
    CLASS CORE ;
    FOREIGN AHHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.530 2.560 3.810 2.840 ;
        RECT  2.850 2.680 3.530 2.840 ;
        RECT  2.760 2.240 2.850 2.840 ;
        RECT  2.660 2.040 2.760 2.840 ;
        RECT  2.570 0.970 2.660 2.840 ;
        RECT  2.440 0.970 2.570 2.400 ;
        RECT  1.890 2.240 2.440 2.400 ;
        RECT  1.610 2.240 1.890 2.520 ;
        END
        ANTENNADIFFAREA 5.178 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.760 0.920 5.920 1.940 ;
        RECT  4.920 0.920 5.760 1.080 ;
        RECT  5.520 1.780 5.760 1.940 ;
        RECT  5.400 1.780 5.520 2.360 ;
        RECT  5.360 1.780 5.400 3.160 ;
        RECT  5.280 2.040 5.360 3.160 ;
        RECT  5.120 2.120 5.280 3.160 ;
        RECT  4.640 0.800 4.920 1.080 ;
        END
        ANTENNADIFFAREA 3.312 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.960 1.560 5.120 1.960 ;
        RECT  4.800 1.560 4.960 2.610 ;
        RECT  4.130 2.450 4.800 2.610 ;
        RECT  3.970 2.450 4.130 3.160 ;
        RECT  2.290 3.000 3.970 3.160 ;
        END
        ANTENNAGATEAREA 0.6504 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 1.340 5.600 1.620 ;
        RECT  5.320 1.240 5.480 1.620 ;
        RECT  4.360 1.240 5.320 1.400 ;
        RECT  4.040 1.240 4.360 1.850 ;
        END
        ANTENNAGATEAREA 0.5448 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.760 -0.280 6.000 0.280 ;
        RECT  5.480 -0.280 5.760 0.600 ;
        RECT  4.120 -0.280 5.480 0.340 ;
        RECT  3.340 -0.280 4.120 0.990 ;
        RECT  0.610 -0.280 3.340 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.900 3.320 6.000 3.880 ;
        RECT  5.680 2.100 5.900 3.880 ;
        RECT  4.920 3.320 5.680 3.880 ;
        RECT  4.640 2.930 4.920 3.880 ;
        RECT  0.890 3.320 4.640 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.160 2.010 4.440 2.290 ;
        RECT  3.330 2.130 4.160 2.290 ;
        RECT  3.210 2.130 3.330 2.520 ;
        RECT  3.140 1.150 3.210 2.520 ;
        RECT  3.050 0.650 3.140 2.520 ;
        RECT  2.860 0.650 3.050 1.310 ;
        RECT  2.280 0.650 2.860 0.810 ;
        RECT  2.090 2.560 2.370 2.840 ;
        RECT  2.120 0.650 2.280 1.410 ;
        RECT  1.450 1.570 2.280 1.850 ;
        RECT  1.130 1.250 2.120 1.410 ;
        RECT  0.370 2.680 2.090 2.840 ;
        RECT  1.740 0.500 1.960 0.950 ;
        RECT  0.370 0.500 1.740 0.660 ;
        RECT  0.690 0.870 1.560 1.090 ;
        RECT  1.290 1.570 1.450 2.510 ;
        RECT  1.150 2.000 1.290 2.510 ;
        RECT  0.690 2.000 1.150 2.160 ;
        RECT  0.850 1.250 1.130 1.840 ;
        RECT  0.530 0.870 0.690 2.160 ;
        RECT  0.090 0.500 0.370 3.160 ;
    END
END AHHCONX2TR

MACRO AHHCINX4TR
    CLASS CORE ;
    FOREIGN AHHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.840 2.720 2.720 ;
        RECT  2.420 1.010 2.510 2.720 ;
        RECT  2.270 1.010 2.420 2.340 ;
        RECT  2.230 1.010 2.270 1.290 ;
        RECT  1.740 2.100 2.270 2.340 ;
        RECT  1.460 2.100 1.740 2.400 ;
        END
        ANTENNADIFFAREA 5.636 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.000 0.980 7.120 2.380 ;
        RECT  6.900 0.980 7.000 3.150 ;
        RECT  5.880 0.980 6.900 1.220 ;
        RECT  6.480 2.140 6.900 3.150 ;
        RECT  5.400 2.140 6.480 2.370 ;
        RECT  5.600 0.440 5.880 1.220 ;
        RECT  4.920 0.980 5.600 1.220 ;
        RECT  5.120 2.140 5.400 3.150 ;
        RECT  4.640 0.440 4.920 1.220 ;
        END
        ANTENNADIFFAREA 7.12 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.720 1.700 6.360 1.980 ;
        RECT  4.760 1.820 5.720 1.980 ;
        RECT  4.720 1.820 4.760 2.580 ;
        RECT  4.440 1.700 4.720 2.580 ;
        RECT  3.170 2.420 4.440 2.580 ;
        RECT  3.010 2.420 3.170 3.100 ;
        RECT  1.340 2.880 3.010 3.100 ;
        END
        ANTENNAGATEAREA 0.9816 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.240 3.860 1.560 ;
        END
        ANTENNAGATEAREA 0.5016 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.400 -0.280 7.200 0.280 ;
        RECT  6.120 -0.280 6.400 0.800 ;
        RECT  5.400 -0.280 6.120 0.280 ;
        RECT  5.120 -0.280 5.400 0.800 ;
        RECT  4.440 -0.280 5.120 0.280 ;
        RECT  4.160 -0.280 4.440 0.670 ;
        RECT  3.470 -0.280 4.160 0.280 ;
        RECT  3.190 -0.280 3.470 0.900 ;
        RECT  0.000 -0.280 3.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.200 3.320 7.200 3.880 ;
        RECT  5.920 2.530 6.200 3.880 ;
        RECT  4.600 3.320 5.920 3.880 ;
        RECT  4.320 2.870 4.600 3.880 ;
        RECT  3.660 3.320 4.320 3.880 ;
        RECT  3.380 2.900 3.660 3.880 ;
        RECT  0.890 3.260 3.380 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.520 1.380 6.740 1.980 ;
        RECT  5.560 1.380 6.520 1.540 ;
        RECT  4.920 1.380 5.560 1.660 ;
        RECT  4.180 1.380 4.920 1.540 ;
        RECT  4.020 0.920 4.180 2.260 ;
        RECT  3.950 0.920 4.020 1.080 ;
        RECT  3.860 1.980 4.020 2.260 ;
        RECT  3.670 0.440 3.950 1.080 ;
        RECT  2.990 1.320 3.120 2.260 ;
        RECT  2.960 0.500 2.990 2.260 ;
        RECT  2.710 0.500 2.960 1.480 ;
        RECT  2.070 0.500 2.710 0.660 ;
        RECT  1.940 2.500 2.220 2.720 ;
        RECT  1.910 0.500 2.070 1.520 ;
        RECT  1.740 1.680 2.020 1.940 ;
        RECT  0.370 2.560 1.940 2.720 ;
        RECT  0.950 1.360 1.910 1.520 ;
        RECT  1.470 0.500 1.750 1.200 ;
        RECT  1.280 1.780 1.740 1.940 ;
        RECT  0.310 0.500 1.470 0.660 ;
        RECT  0.630 0.820 1.290 1.040 ;
        RECT  1.110 1.780 1.280 2.400 ;
        RECT  1.000 1.870 1.110 2.400 ;
        RECT  0.630 1.870 1.000 2.030 ;
        RECT  0.790 1.360 0.950 1.710 ;
        RECT  0.470 0.820 0.630 2.030 ;
        RECT  0.310 2.190 0.370 3.160 ;
        RECT  0.090 0.500 0.310 3.160 ;
    END
END AHHCINX4TR

MACRO AHHCINX2TR
    CLASS CORE ;
    FOREIGN AHHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.840 2.720 1.160 ;
        RECT  2.420 0.880 2.440 1.160 ;
        RECT  2.260 0.880 2.420 2.720 ;
        END
        ANTENNADIFFAREA 5.864 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.320 1.930 4.760 2.720 ;
        RECT  4.280 0.920 4.320 2.720 ;
        RECT  4.160 0.920 4.280 2.360 ;
        RECT  3.880 0.800 4.160 1.080 ;
        END
        ANTENNADIFFAREA 3.168 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.920 1.580 5.200 3.040 ;
        RECT  3.960 2.880 4.920 3.040 ;
        RECT  3.680 1.330 3.960 3.040 ;
        RECT  2.800 2.880 3.680 3.040 ;
        RECT  2.740 1.680 2.800 3.040 ;
        RECT  2.580 1.680 2.740 3.100 ;
        RECT  1.050 2.880 2.580 3.100 ;
        END
        ANTENNAGATEAREA 0.6696 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.480 5.410 0.640 ;
        RECT  3.360 0.480 3.520 1.640 ;
        RECT  3.280 1.240 3.360 1.640 ;
        END
        ANTENNAGATEAREA 0.3912 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 -0.280 6.000 0.280 ;
        RECT  4.400 -0.280 4.680 0.320 ;
        RECT  3.640 -0.280 4.400 0.280 ;
        RECT  3.360 -0.280 3.640 0.320 ;
        RECT  0.890 -0.280 3.360 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.280 3.320 6.000 3.880 ;
        RECT  0.890 3.260 5.280 3.880 ;
        RECT  0.610 3.200 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.630 1.260 5.910 2.490 ;
        RECT  5.610 1.260 5.630 1.420 ;
        RECT  5.330 0.910 5.610 1.420 ;
        RECT  4.760 1.260 5.330 1.420 ;
        RECT  4.600 1.260 4.760 1.770 ;
        RECT  4.480 1.490 4.600 1.770 ;
        RECT  3.120 2.030 3.240 2.720 ;
        RECT  3.100 1.150 3.120 2.720 ;
        RECT  2.960 0.440 3.100 2.720 ;
        RECT  2.880 0.440 2.960 1.310 ;
        RECT  2.100 0.440 2.880 0.600 ;
        RECT  1.940 0.440 2.100 1.540 ;
        RECT  1.720 2.140 2.000 2.720 ;
        RECT  1.070 1.380 1.940 1.540 ;
        RECT  1.510 1.700 1.790 1.980 ;
        RECT  1.500 0.500 1.780 1.220 ;
        RECT  0.370 2.560 1.720 2.720 ;
        RECT  1.420 1.820 1.510 1.980 ;
        RECT  0.310 0.500 1.500 0.660 ;
        RECT  1.230 1.820 1.420 2.400 ;
        RECT  0.690 0.840 1.290 1.060 ;
        RECT  1.140 1.890 1.230 2.400 ;
        RECT  0.690 1.890 1.140 2.050 ;
        RECT  0.850 1.380 1.070 1.730 ;
        RECT  0.530 0.840 0.690 2.050 ;
        RECT  0.310 1.910 0.370 3.160 ;
        RECT  0.090 0.500 0.310 3.160 ;
    END
END AHHCINX2TR

MACRO AHCSHCONX4TR
    CLASS CORE ;
    FOREIGN AHCSHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 0.440 7.920 3.160 ;
        RECT  7.640 0.440 7.680 1.230 ;
        RECT  7.600 1.840 7.680 3.160 ;
        RECT  7.280 1.840 7.600 2.560 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.720 2.380 7.120 2.760 ;
        END
        ANTENNAGATEAREA 0.2784 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 2.160 1.750 3.160 ;
        RECT  0.790 2.160 1.590 2.320 ;
        RECT  1.270 0.440 1.430 1.240 ;
        RECT  0.510 1.080 1.270 1.240 ;
        RECT  0.510 2.160 0.790 3.160 ;
        RECT  0.480 1.080 0.510 3.160 ;
        RECT  0.350 1.080 0.480 2.320 ;
        END
        ANTENNADIFFAREA 5.148 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.680 3.030 2.600 ;
        RECT  2.870 1.560 2.910 2.600 ;
        RECT  2.750 1.560 2.870 1.840 ;
        RECT  2.720 2.440 2.870 2.600 ;
        RECT  2.480 2.440 2.720 2.760 ;
        RECT  2.070 2.440 2.480 2.600 ;
        RECT  1.910 1.840 2.070 2.600 ;
        RECT  1.630 1.840 1.910 2.000 ;
        RECT  1.070 1.720 1.630 2.000 ;
        END
        ANTENNAGATEAREA 0.7872 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.420 2.090 1.580 ;
        RECT  1.810 1.240 1.920 1.580 ;
        RECT  1.680 1.240 1.810 1.560 ;
        RECT  0.830 1.400 1.680 1.560 ;
        RECT  0.670 1.400 0.830 1.680 ;
        END
        ANTENNAGATEAREA 0.7176 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.870 -0.280 8.000 0.280 ;
        RECT  4.590 -0.280 4.870 0.610 ;
        RECT  2.230 -0.280 4.590 0.280 ;
        RECT  2.070 -0.280 2.230 1.080 ;
        RECT  0.590 -0.280 2.070 0.280 ;
        RECT  0.430 -0.280 0.590 0.800 ;
        RECT  0.000 -0.280 0.430 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.300 3.320 8.000 3.880 ;
        RECT  7.020 3.100 7.300 3.880 ;
        RECT  4.630 3.320 7.020 3.880 ;
        RECT  4.350 3.020 4.630 3.880 ;
        RECT  2.230 3.320 4.350 3.880 ;
        RECT  2.070 2.910 2.230 3.880 ;
        RECT  1.270 3.320 2.070 3.880 ;
        RECT  1.110 2.480 1.270 3.880 ;
        RECT  0.310 3.320 1.110 3.880 ;
        RECT  0.150 2.480 0.310 3.880 ;
        RECT  0.000 3.320 0.150 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.480 1.400 7.520 1.680 ;
        RECT  7.320 0.440 7.480 1.680 ;
        RECT  5.940 0.440 7.320 0.600 ;
        RECT  6.820 0.850 6.940 1.010 ;
        RECT  6.820 1.970 6.940 2.130 ;
        RECT  6.660 0.850 6.820 2.130 ;
        RECT  6.420 1.520 6.660 1.680 ;
        RECT  6.260 0.790 6.420 1.080 ;
        RECT  6.260 1.910 6.420 3.160 ;
        RECT  6.100 0.790 6.260 2.200 ;
        RECT  4.950 3.000 6.260 3.160 ;
        RECT  5.780 0.440 5.940 2.740 ;
        RECT  5.360 0.440 5.520 2.840 ;
        RECT  5.300 0.440 5.360 0.930 ;
        RECT  5.240 2.680 5.360 2.840 ;
        RECT  4.430 0.770 5.300 0.930 ;
        RECT  4.970 1.090 5.090 1.250 ;
        RECT  4.970 1.910 5.030 2.190 ;
        RECT  4.810 1.090 4.970 2.450 ;
        RECT  4.790 2.700 4.950 3.160 ;
        RECT  3.670 2.290 4.810 2.450 ;
        RECT  3.350 2.700 4.790 2.860 ;
        RECT  4.270 0.440 4.430 1.640 ;
        RECT  2.710 0.440 4.270 0.600 ;
        RECT  3.950 0.850 4.110 2.130 ;
        RECT  3.830 1.970 3.950 2.130 ;
        RECT  3.510 1.580 3.670 2.450 ;
        RECT  3.350 0.850 3.510 1.130 ;
        RECT  3.190 0.970 3.350 2.860 ;
        RECT  2.590 0.440 2.710 1.310 ;
        RECT  2.590 2.000 2.710 2.280 ;
        RECT  2.550 0.440 2.590 2.280 ;
        RECT  2.430 1.150 2.550 2.160 ;
    END
END AHCSHCONX4TR

MACRO AHCSHCONX2TR
    CLASS CORE ;
    FOREIGN AHCSHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 0.440 7.120 3.160 ;
        RECT  6.720 0.440 6.960 1.150 ;
        RECT  6.720 1.910 6.960 3.160 ;
        END
        ANTENNADIFFAREA 3.458 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 2.440 6.080 2.760 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 2.170 0.850 3.160 ;
        RECT  0.320 2.170 0.570 2.360 ;
        RECT  0.320 0.440 0.530 1.280 ;
        RECT  0.250 0.440 0.320 2.360 ;
        RECT  0.080 1.120 0.250 2.360 ;
        END
        ANTENNADIFFAREA 3.136 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.550 2.070 2.720 ;
        RECT  1.680 1.550 1.910 1.960 ;
        RECT  1.170 2.560 1.910 2.720 ;
        RECT  1.010 1.850 1.170 2.720 ;
        RECT  0.710 1.850 1.010 2.010 ;
        RECT  0.490 1.730 0.710 2.010 ;
        END
        ANTENNAGATEAREA 0.5496 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.220 1.160 1.560 ;
        RECT  0.840 1.220 1.130 1.620 ;
        END
        ANTENNAGATEAREA 0.4752 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.480 -0.280 7.200 0.280 ;
        RECT  3.970 -0.280 6.480 0.340 ;
        RECT  3.690 -0.280 3.970 0.580 ;
        RECT  1.330 -0.280 3.690 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.000 -0.280 1.050 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.520 3.320 7.200 3.880 ;
        RECT  6.240 1.910 6.520 3.880 ;
        RECT  6.200 3.200 6.240 3.880 ;
        RECT  3.790 3.260 6.200 3.880 ;
        RECT  3.510 2.960 3.790 3.880 ;
        RECT  1.330 3.320 3.510 3.880 ;
        RECT  1.050 2.880 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 2.540 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.440 1.390 6.720 1.670 ;
        RECT  6.300 1.390 6.440 1.550 ;
        RECT  6.140 0.500 6.300 1.550 ;
        RECT  5.040 0.500 6.140 0.660 ;
        RECT  5.860 1.000 5.980 1.280 ;
        RECT  5.860 1.920 5.980 2.200 ;
        RECT  5.700 1.000 5.860 2.200 ;
        RECT  5.520 1.520 5.700 1.800 ;
        RECT  5.360 0.850 5.520 1.130 ;
        RECT  5.360 1.960 5.520 2.890 ;
        RECT  5.200 0.850 5.360 3.100 ;
        RECT  4.110 2.940 5.200 3.100 ;
        RECT  4.880 0.500 5.040 2.780 ;
        RECT  4.760 0.500 4.880 1.130 ;
        RECT  4.760 2.110 4.880 2.780 ;
        RECT  4.400 0.500 4.560 2.780 ;
        RECT  4.280 0.500 4.400 0.900 ;
        RECT  4.280 2.500 4.400 2.780 ;
        RECT  3.590 0.740 4.280 0.900 ;
        RECT  4.070 1.060 4.190 1.280 ;
        RECT  4.070 1.880 4.190 2.200 ;
        RECT  3.950 2.640 4.110 3.100 ;
        RECT  3.910 1.060 4.070 2.480 ;
        RECT  2.450 2.640 3.950 2.800 ;
        RECT  2.830 2.320 3.910 2.480 ;
        RECT  3.530 0.740 3.590 1.610 ;
        RECT  3.370 0.440 3.530 1.610 ;
        RECT  1.810 0.440 3.370 0.600 ;
        RECT  3.210 1.980 3.270 2.160 ;
        RECT  2.990 0.850 3.210 2.160 ;
        RECT  2.610 1.590 2.830 2.480 ;
        RECT  2.450 0.850 2.610 1.130 ;
        RECT  2.330 0.850 2.450 2.800 ;
        RECT  2.230 0.970 2.330 2.800 ;
        RECT  1.530 0.440 1.810 1.280 ;
        RECT  1.530 2.120 1.750 2.400 ;
        RECT  1.520 1.120 1.530 1.280 ;
        RECT  1.520 2.120 1.530 2.280 ;
        RECT  1.360 1.120 1.520 2.280 ;
    END
END AHCSHCONX2TR

MACRO AHCSHCINX4TR
    CLASS CORE ;
    FOREIGN AHCSHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.600 0.440 7.760 3.160 ;
        RECT  7.440 0.440 7.600 1.230 ;
        RECT  7.440 1.840 7.600 3.160 ;
        RECT  7.280 1.840 7.440 2.560 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.480 2.350 6.760 3.100 ;
        END
        ANTENNAGATEAREA 0.2784 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.710 1.820 0.990 ;
        RECT  0.860 0.830 1.540 0.990 ;
        RECT  0.880 1.910 1.120 3.160 ;
        RECT  0.360 1.910 0.880 2.070 ;
        RECT  0.580 0.710 0.860 0.990 ;
        RECT  0.360 0.830 0.580 0.990 ;
        RECT  0.080 0.830 0.360 2.070 ;
        END
        ANTENNADIFFAREA 4.896 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 2.350 2.720 2.630 ;
        RECT  1.520 2.350 2.440 2.510 ;
        RECT  1.280 1.470 1.520 2.510 ;
        RECT  1.100 1.470 1.280 1.750 ;
        END
        ANTENNAGATEAREA 0.8136 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.470 2.400 1.750 ;
        RECT  1.960 1.590 2.120 1.750 ;
        RECT  1.680 1.590 1.960 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.200 -0.280 8.000 0.280 ;
        RECT  6.920 -0.280 7.200 0.400 ;
        RECT  4.380 -0.280 6.920 0.280 ;
        RECT  4.100 -0.280 4.380 0.610 ;
        RECT  2.300 -0.280 4.100 0.280 ;
        RECT  2.020 -0.280 2.300 0.670 ;
        RECT  1.340 -0.280 2.020 0.280 ;
        RECT  1.060 -0.280 1.340 0.670 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 0.670 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.200 3.320 8.000 3.880 ;
        RECT  6.920 2.800 7.200 3.880 ;
        RECT  4.540 3.260 6.920 3.880 ;
        RECT  4.260 2.990 4.540 3.880 ;
        RECT  1.980 3.320 4.260 3.880 ;
        RECT  1.700 2.930 1.980 3.880 ;
        RECT  0.380 3.320 1.700 3.880 ;
        RECT  0.100 2.230 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.280 1.470 7.440 1.650 ;
        RECT  7.120 0.560 7.280 1.650 ;
        RECT  6.560 0.560 7.120 0.720 ;
        RECT  6.500 1.030 6.720 2.190 ;
        RECT  6.400 0.440 6.560 0.720 ;
        RECT  6.440 1.030 6.500 1.740 ;
        RECT  6.400 1.460 6.440 1.740 ;
        RECT  5.760 0.440 6.400 0.600 ;
        RECT  6.240 1.910 6.320 2.860 ;
        RECT  6.200 0.790 6.240 2.860 ;
        RECT  6.040 0.790 6.200 3.100 ;
        RECT  5.960 0.790 6.040 1.070 ;
        RECT  4.860 2.940 6.040 3.100 ;
        RECT  5.760 2.050 5.840 2.780 ;
        RECT  5.560 0.440 5.760 2.780 ;
        RECT  5.480 0.440 5.560 1.070 ;
        RECT  5.280 2.050 5.360 2.330 ;
        RECT  5.080 0.520 5.280 2.330 ;
        RECT  5.000 0.520 5.080 0.930 ;
        RECT  4.180 0.770 5.000 0.930 ;
        RECT  4.780 1.090 4.900 1.310 ;
        RECT  4.780 1.910 4.900 2.190 ;
        RECT  4.700 2.670 4.860 3.100 ;
        RECT  4.620 1.090 4.780 2.510 ;
        RECT  3.540 2.670 4.700 2.830 ;
        RECT  3.420 2.350 4.620 2.510 ;
        RECT  4.180 1.380 4.300 1.660 ;
        RECT  4.020 0.770 4.180 1.660 ;
        RECT  3.580 0.770 4.020 0.930 ;
        RECT  3.740 1.910 4.020 2.190 ;
        RECT  3.740 1.090 3.860 1.310 ;
        RECT  3.580 1.090 3.740 2.190 ;
        RECT  3.420 0.710 3.580 0.930 ;
        RECT  3.260 2.670 3.540 2.950 ;
        RECT  2.780 0.710 3.420 0.870 ;
        RECT  3.200 1.560 3.420 2.510 ;
        RECT  3.040 1.030 3.260 1.310 ;
        RECT  3.040 2.670 3.260 2.830 ;
        RECT  2.980 1.030 3.040 2.830 ;
        RECT  2.880 1.150 2.980 2.830 ;
        RECT  2.720 0.440 2.780 0.870 ;
        RECT  2.560 0.440 2.720 2.070 ;
        RECT  2.500 0.440 2.560 1.310 ;
        RECT  2.460 1.910 2.560 2.070 ;
        RECT  1.960 1.150 2.500 1.310 ;
        RECT  2.180 1.910 2.460 2.190 ;
        RECT  1.680 1.150 1.960 1.430 ;
        RECT  0.740 1.150 1.680 1.310 ;
        RECT  0.520 1.150 0.740 1.430 ;
    END
END AHCSHCINX4TR

MACRO AHCSHCINX2TR
    CLASS CORE ;
    FOREIGN AHCSHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.730 0.440 6.890 3.160 ;
        RECT  6.570 0.440 6.730 1.230 ;
        RECT  6.480 1.910 6.730 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.200 2.040 6.320 2.360 ;
        RECT  6.040 2.040 6.200 2.510 ;
        RECT  5.860 2.350 6.040 2.510 ;
        RECT  5.580 2.350 5.860 3.100 ;
        END
        ANTENNAGATEAREA 0.2784 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.720 0.850 1.000 ;
        RECT  0.240 0.840 0.570 1.000 ;
        RECT  0.240 1.910 0.320 3.160 ;
        RECT  0.080 0.840 0.240 3.160 ;
        END
        ANTENNADIFFAREA 3.376 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 2.360 1.810 2.640 ;
        RECT  0.720 2.360 1.590 2.520 ;
        RECT  0.680 1.640 0.720 2.520 ;
        RECT  0.480 1.240 0.680 2.520 ;
        RECT  0.400 1.240 0.480 1.520 ;
        END
        ANTENNAGATEAREA 0.576 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.480 1.490 1.760 ;
        RECT  1.160 1.600 1.270 1.760 ;
        RECT  0.880 1.600 1.160 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.330 -0.280 7.200 0.280 ;
        RECT  6.050 -0.280 6.330 0.400 ;
        RECT  3.430 -0.280 6.050 0.280 ;
        RECT  3.150 -0.280 3.430 0.610 ;
        RECT  1.330 -0.280 3.150 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.300 3.320 7.200 3.880 ;
        RECT  6.020 2.800 6.300 3.880 ;
        RECT  3.630 3.260 6.020 3.880 ;
        RECT  3.350 2.990 3.630 3.880 ;
        RECT  1.180 3.320 3.350 3.880 ;
        RECT  0.900 2.930 1.180 3.880 ;
        RECT  0.000 3.320 0.900 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.410 1.470 6.570 1.750 ;
        RECT  6.250 0.560 6.410 1.750 ;
        RECT  5.690 0.560 6.250 0.720 ;
        RECT  5.600 1.030 5.880 2.190 ;
        RECT  5.530 0.440 5.690 0.720 ;
        RECT  5.530 1.460 5.600 1.740 ;
        RECT  4.890 0.440 5.530 0.600 ;
        RECT  5.370 1.910 5.420 2.860 ;
        RECT  5.300 0.790 5.370 2.860 ;
        RECT  5.140 0.790 5.300 3.100 ;
        RECT  5.090 0.790 5.140 1.070 ;
        RECT  3.950 2.940 5.140 3.100 ;
        RECT  4.890 2.050 4.940 2.780 ;
        RECT  4.660 0.440 4.890 2.780 ;
        RECT  4.610 0.440 4.660 1.070 ;
        RECT  4.410 2.050 4.460 2.780 ;
        RECT  4.180 0.770 4.410 2.780 ;
        RECT  4.130 0.770 4.180 1.050 ;
        RECT  3.310 0.770 4.130 0.930 ;
        RECT  3.950 1.910 3.990 2.190 ;
        RECT  3.870 1.090 3.950 2.190 ;
        RECT  3.790 2.670 3.950 3.100 ;
        RECT  3.710 1.090 3.870 2.510 ;
        RECT  2.630 2.670 3.790 2.830 ;
        RECT  3.670 1.090 3.710 1.310 ;
        RECT  2.510 2.350 3.710 2.510 ;
        RECT  3.030 0.770 3.310 1.660 ;
        RECT  2.870 1.910 3.110 2.190 ;
        RECT  2.610 0.770 3.030 0.930 ;
        RECT  2.710 1.090 2.870 2.190 ;
        RECT  2.590 1.090 2.710 1.310 ;
        RECT  2.350 2.670 2.630 2.950 ;
        RECT  2.450 0.440 2.610 0.930 ;
        RECT  2.290 1.560 2.510 2.510 ;
        RECT  1.810 0.440 2.450 0.600 ;
        RECT  2.130 2.670 2.350 2.830 ;
        RECT  2.130 1.030 2.290 1.310 ;
        RECT  1.970 1.030 2.130 2.830 ;
        RECT  1.660 0.440 1.810 2.080 ;
        RECT  1.650 0.440 1.660 2.200 ;
        RECT  1.530 0.440 1.650 1.320 ;
        RECT  1.380 1.920 1.650 2.200 ;
        RECT  1.080 1.160 1.530 1.320 ;
        RECT  0.860 1.160 1.080 1.440 ;
    END
END AHCSHCINX2TR

MACRO AFHCONX4TR
    CLASS CORE ;
    FOREIGN AFHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.920 0.470 13.100 3.160 ;
        RECT  12.820 0.470 12.920 1.310 ;
        RECT  12.820 1.910 12.920 3.160 ;
        RECT  12.480 2.240 12.820 2.960 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.480 1.020 7.660 1.300 ;
        RECT  7.480 2.040 7.640 2.320 ;
        RECT  7.320 0.760 7.480 2.320 ;
        RECT  6.540 0.760 7.320 0.920 ;
        RECT  6.460 0.760 6.540 1.200 ;
        RECT  6.300 0.760 6.460 2.780 ;
        RECT  6.080 1.840 6.300 2.780 ;
        END
        ANTENNADIFFAREA 7.724 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.720 1.380 9.020 1.660 ;
        RECT  8.480 1.240 8.720 1.660 ;
        RECT  8.320 1.380 8.480 1.660 ;
        END
        ANTENNAGATEAREA 1.0656 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.560 5.120 1.960 ;
        END
        ANTENNAGATEAREA 1.0224 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.720 1.580 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.620 -0.280 13.200 0.280 ;
        RECT  12.340 -0.280 12.620 1.200 ;
        RECT  10.300 -0.280 12.340 0.280 ;
        RECT  10.020 -0.280 10.300 0.320 ;
        RECT  9.320 -0.280 10.020 0.280 ;
        RECT  9.040 -0.280 9.320 0.320 ;
        RECT  8.280 -0.280 9.040 0.280 ;
        RECT  8.000 -0.280 8.280 0.320 ;
        RECT  5.360 -0.280 8.000 0.280 ;
        RECT  5.080 -0.280 5.360 0.400 ;
        RECT  0.890 -0.280 5.080 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.580 3.320 13.200 3.880 ;
        RECT  12.300 3.240 12.580 3.880 ;
        RECT  9.990 3.320 12.300 3.880 ;
        RECT  9.710 2.990 9.990 3.880 ;
        RECT  9.030 3.320 9.710 3.880 ;
        RECT  8.750 2.990 9.030 3.880 ;
        RECT  5.400 3.260 8.750 3.880 ;
        RECT  5.120 2.940 5.400 3.880 ;
        RECT  0.850 3.320 5.120 3.880 ;
        RECT  0.570 2.070 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.660 1.470 12.760 1.750 ;
        RECT  12.500 1.470 12.660 1.960 ;
        RECT  12.180 1.800 12.500 1.960 ;
        RECT  12.020 0.770 12.180 1.640 ;
        RECT  12.020 1.800 12.180 3.120 ;
        RECT  10.940 0.770 12.020 0.930 ;
        RECT  11.420 2.960 12.020 3.120 ;
        RECT  11.740 1.090 11.860 1.250 ;
        RECT  11.740 2.110 11.860 2.800 ;
        RECT  11.580 1.090 11.740 2.800 ;
        RECT  10.620 0.440 11.590 0.600 ;
        RECT  11.260 1.090 11.420 3.120 ;
        RECT  11.100 1.090 11.260 1.310 ;
        RECT  11.100 2.190 11.260 2.350 ;
        RECT  10.880 2.670 11.100 3.160 ;
        RECT  10.780 0.770 10.940 2.390 ;
        RECT  8.550 2.670 10.880 2.830 ;
        RECT  9.500 0.800 10.780 1.080 ;
        RECT  10.470 2.230 10.780 2.390 ;
        RECT  10.460 0.440 10.620 0.640 ;
        RECT  10.400 1.240 10.620 1.980 ;
        RECT  10.190 2.230 10.470 2.510 ;
        RECT  9.340 0.480 10.460 0.640 ;
        RECT  9.340 1.240 10.400 1.400 ;
        RECT  8.270 2.290 10.190 2.510 ;
        RECT  7.990 1.910 9.510 2.130 ;
        RECT  9.180 0.480 9.340 1.400 ;
        RECT  7.760 0.480 9.180 0.640 ;
        RECT  7.990 0.860 8.800 1.080 ;
        RECT  8.390 2.670 8.550 3.100 ;
        RECT  6.840 2.940 8.390 3.100 ;
        RECT  7.830 0.860 7.990 2.780 ;
        RECT  7.160 2.620 7.830 2.780 ;
        RECT  7.600 0.440 7.760 0.640 ;
        RECT  6.140 0.440 7.600 0.600 ;
        RECT  7.000 1.080 7.160 2.780 ;
        RECT  6.840 1.080 7.000 1.300 ;
        RECT  6.680 1.610 6.840 3.100 ;
        RECT  5.720 2.940 6.680 3.100 ;
        RECT  5.980 0.440 6.140 1.480 ;
        RECT  4.500 0.560 5.980 0.720 ;
        RECT  5.940 1.320 5.980 1.480 ;
        RECT  5.780 1.320 5.940 1.650 ;
        RECT  5.440 2.300 5.880 2.460 ;
        RECT  5.600 0.880 5.820 1.160 ;
        RECT  5.560 2.620 5.720 3.100 ;
        RECT  5.440 1.000 5.600 1.160 ;
        RECT  4.930 2.620 5.560 2.780 ;
        RECT  5.280 1.000 5.440 2.460 ;
        RECT  4.770 2.620 4.930 3.150 ;
        RECT  4.720 2.120 4.920 2.370 ;
        RECT  4.720 1.040 4.800 1.310 ;
        RECT  2.420 2.990 4.770 3.150 ;
        RECT  4.560 1.040 4.720 2.370 ;
        RECT  4.360 2.670 4.580 2.830 ;
        RECT  4.140 1.300 4.560 1.480 ;
        RECT  4.220 0.550 4.500 0.850 ;
        RECT  4.200 1.640 4.360 2.830 ;
        RECT  3.540 0.550 4.220 0.710 ;
        RECT  3.980 1.640 4.200 1.800 ;
        RECT  2.800 2.670 4.200 2.830 ;
        RECT  3.880 1.960 4.040 2.240 ;
        RECT  3.820 0.870 3.980 1.800 ;
        RECT  3.660 1.960 3.880 2.120 ;
        RECT  3.700 0.870 3.820 1.150 ;
        RECT  3.540 1.310 3.660 2.120 ;
        RECT  3.500 0.550 3.540 2.120 ;
        RECT  3.380 0.550 3.500 1.470 ;
        RECT  3.280 0.730 3.380 1.010 ;
        RECT  3.120 2.350 3.240 2.510 ;
        RECT  2.960 0.450 3.120 2.510 ;
        RECT  1.210 0.450 2.960 0.610 ;
        RECT  2.640 0.770 2.800 2.830 ;
        RECT  1.930 0.770 2.640 0.930 ;
        RECT  2.200 1.090 2.420 3.150 ;
        RECT  1.720 2.390 2.200 3.150 ;
        RECT  1.770 0.770 1.930 1.250 ;
        RECT  1.460 0.880 1.770 1.250 ;
        RECT  1.250 0.880 1.460 3.160 ;
        RECT  1.050 2.450 1.250 3.160 ;
        RECT  1.050 0.450 1.210 0.660 ;
        RECT  0.910 0.920 1.070 1.910 ;
        RECT  0.370 0.500 1.050 0.660 ;
        RECT  0.370 0.920 0.910 1.080 ;
        RECT  0.370 1.750 0.910 1.910 ;
        RECT  0.090 0.500 0.370 1.080 ;
        RECT  0.090 1.750 0.370 3.160 ;
    END
END AFHCONX4TR

MACRO AFHCONX2TR
    CLASS CORE ;
    FOREIGN AFHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.940 0.470 11.100 3.160 ;
        RECT  10.820 0.470 10.940 1.310 ;
        RECT  10.880 1.910 10.940 3.160 ;
        RECT  10.820 2.240 10.880 3.160 ;
        RECT  10.480 2.240 10.820 2.960 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.460 0.760 6.540 1.200 ;
        RECT  6.300 0.760 6.460 2.780 ;
        RECT  6.080 1.840 6.300 2.780 ;
        END
        ANTENNADIFFAREA 4.426 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.520 1.380 7.650 1.660 ;
        RECT  7.280 1.240 7.520 1.660 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.560 5.120 1.960 ;
        END
        ANTENNAGATEAREA 1.0224 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.240 0.720 1.580 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.620 -0.280 11.200 0.280 ;
        RECT  10.340 -0.280 10.620 0.610 ;
        RECT  8.020 -0.280 10.340 0.280 ;
        RECT  7.740 -0.280 8.020 0.320 ;
        RECT  5.360 -0.280 7.740 0.280 ;
        RECT  5.080 -0.280 5.360 0.400 ;
        RECT  0.890 -0.280 5.080 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.580 3.320 11.200 3.880 ;
        RECT  10.300 3.240 10.580 3.880 ;
        RECT  8.200 3.320 10.300 3.880 ;
        RECT  7.920 2.990 8.200 3.880 ;
        RECT  5.400 3.320 7.920 3.880 ;
        RECT  5.120 2.940 5.400 3.880 ;
        RECT  0.850 3.320 5.120 3.880 ;
        RECT  0.570 2.070 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.720 1.470 10.780 1.750 ;
        RECT  10.560 1.470 10.720 1.960 ;
        RECT  10.320 1.800 10.560 1.960 ;
        RECT  10.220 0.770 10.380 1.640 ;
        RECT  10.160 1.800 10.320 2.720 ;
        RECT  9.060 0.770 10.220 0.930 ;
        RECT  9.520 2.560 10.160 2.720 ;
        RECT  10.000 1.090 10.040 1.250 ;
        RECT  9.840 1.090 10.000 2.400 ;
        RECT  9.760 1.090 9.840 1.250 ;
        RECT  8.620 0.440 9.710 0.600 ;
        RECT  9.360 1.090 9.520 2.720 ;
        RECT  9.140 3.000 9.370 3.160 ;
        RECT  9.220 1.090 9.360 1.310 ;
        RECT  9.060 1.470 9.200 2.510 ;
        RECT  8.980 2.670 9.140 3.160 ;
        RECT  9.040 0.770 9.060 2.510 ;
        RECT  8.900 0.770 9.040 1.630 ;
        RECT  8.400 2.350 9.040 2.510 ;
        RECT  7.520 2.670 8.980 2.830 ;
        RECT  8.800 0.770 8.900 1.080 ;
        RECT  8.660 1.810 8.840 2.140 ;
        RECT  8.340 0.800 8.800 1.080 ;
        RECT  8.040 1.860 8.660 2.140 ;
        RECT  8.460 0.440 8.620 0.640 ;
        RECT  8.040 0.480 8.460 0.640 ;
        RECT  7.880 0.480 8.040 2.140 ;
        RECT  7.170 0.480 7.880 0.640 ;
        RECT  7.100 2.100 7.660 2.260 ;
        RECT  7.360 2.670 7.520 3.100 ;
        RECT  6.780 2.940 7.360 3.100 ;
        RECT  7.010 0.440 7.170 0.640 ;
        RECT  6.940 1.020 7.100 2.780 ;
        RECT  6.140 0.440 7.010 0.600 ;
        RECT  6.930 1.020 6.940 1.300 ;
        RECT  6.620 1.610 6.780 3.100 ;
        RECT  5.720 2.940 6.620 3.100 ;
        RECT  5.980 0.440 6.140 1.480 ;
        RECT  4.500 0.560 5.980 0.720 ;
        RECT  5.940 1.320 5.980 1.480 ;
        RECT  5.780 1.320 5.940 1.650 ;
        RECT  5.440 2.300 5.880 2.460 ;
        RECT  5.600 0.880 5.820 1.160 ;
        RECT  5.560 2.620 5.720 3.100 ;
        RECT  5.440 1.000 5.600 1.160 ;
        RECT  4.930 2.620 5.560 2.780 ;
        RECT  5.280 1.000 5.440 2.460 ;
        RECT  4.770 2.620 4.930 3.150 ;
        RECT  4.720 2.120 4.920 2.370 ;
        RECT  4.720 1.040 4.800 1.310 ;
        RECT  2.390 2.990 4.770 3.150 ;
        RECT  4.560 1.040 4.720 2.370 ;
        RECT  4.360 2.670 4.580 2.830 ;
        RECT  4.140 1.300 4.560 1.480 ;
        RECT  4.220 0.550 4.500 0.850 ;
        RECT  4.200 1.640 4.360 2.830 ;
        RECT  3.540 0.550 4.220 0.710 ;
        RECT  3.980 1.640 4.200 1.800 ;
        RECT  2.800 2.670 4.200 2.830 ;
        RECT  3.880 1.960 4.040 2.240 ;
        RECT  3.820 0.870 3.980 1.800 ;
        RECT  3.660 1.960 3.880 2.120 ;
        RECT  3.700 0.870 3.820 1.150 ;
        RECT  3.540 1.310 3.660 2.120 ;
        RECT  3.500 0.550 3.540 2.120 ;
        RECT  3.380 0.550 3.500 1.470 ;
        RECT  3.280 0.730 3.380 1.010 ;
        RECT  3.120 2.350 3.240 2.510 ;
        RECT  2.960 0.450 3.120 2.510 ;
        RECT  1.210 0.450 2.960 0.610 ;
        RECT  2.640 0.770 2.800 2.830 ;
        RECT  1.850 0.770 2.640 0.930 ;
        RECT  2.170 1.090 2.390 3.150 ;
        RECT  1.720 2.450 2.170 3.150 ;
        RECT  1.520 0.770 1.850 1.120 ;
        RECT  1.400 0.880 1.520 1.120 ;
        RECT  1.230 0.880 1.400 3.160 ;
        RECT  1.110 2.450 1.230 3.160 ;
        RECT  1.050 0.450 1.210 0.660 ;
        RECT  0.910 0.920 1.070 1.910 ;
        RECT  0.370 0.500 1.050 0.660 ;
        RECT  0.370 0.920 0.910 1.080 ;
        RECT  0.370 1.750 0.910 1.910 ;
        RECT  0.090 0.500 0.370 1.080 ;
        RECT  0.090 1.750 0.370 3.160 ;
    END
END AFHCONX2TR

MACRO AFHCINX4TR
    CLASS CORE ;
    FOREIGN AFHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.400 0.880 10.620 2.090 ;
        RECT  10.340 0.880 10.400 2.560 ;
        RECT  10.080 1.840 10.340 2.560 ;
        END
        ANTENNADIFFAREA 2.57 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.600 1.020 9.860 1.240 ;
        RECT  9.580 1.020 9.600 2.230 ;
        RECT  9.280 1.080 9.580 2.230 ;
        RECT  9.020 2.010 9.280 2.230 ;
        RECT  8.680 2.010 9.020 2.290 ;
        RECT  8.430 0.760 8.680 2.290 ;
        RECT  7.820 0.760 8.430 0.920 ;
        RECT  8.000 2.010 8.430 2.290 ;
        RECT  7.680 1.840 8.000 2.560 ;
        RECT  7.660 0.760 7.820 1.330 ;
        RECT  7.270 2.010 7.680 2.290 ;
        RECT  7.500 1.070 7.660 1.330 ;
        RECT  6.940 2.010 7.270 2.720 ;
        END
        ANTENNADIFFAREA 8.996 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.440 1.240 14.760 1.620 ;
        END
        ANTENNAGATEAREA 1.056 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.680 1.570 5.920 1.960 ;
        END
        ANTENNAGATEAREA 0.7968 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.490 2.360 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.720 -0.280 16.000 0.280 ;
        RECT  15.440 -0.280 15.720 1.130 ;
        RECT  14.760 -0.280 15.440 0.280 ;
        RECT  14.480 -0.280 14.760 1.010 ;
        RECT  13.760 -0.280 14.480 0.280 ;
        RECT  13.480 -0.280 13.760 0.400 ;
        RECT  10.330 -0.280 13.480 0.280 ;
        RECT  10.050 -0.280 10.330 0.400 ;
        RECT  0.890 -0.280 10.050 0.280 ;
        RECT  0.610 -0.280 0.890 0.370 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.720 3.320 16.000 3.880 ;
        RECT  15.440 2.050 15.720 3.880 ;
        RECT  14.760 3.320 15.440 3.880 ;
        RECT  14.480 2.990 14.760 3.880 ;
        RECT  13.800 3.320 14.480 3.880 ;
        RECT  13.520 2.990 13.800 3.880 ;
        RECT  10.880 3.320 13.520 3.880 ;
        RECT  10.600 2.710 10.880 3.880 ;
        RECT  9.840 3.320 10.600 3.880 ;
        RECT  9.560 2.790 9.840 3.880 ;
        RECT  6.280 3.320 9.560 3.880 ;
        RECT  6.000 2.190 6.280 3.880 ;
        RECT  0.850 3.260 6.000 3.880 ;
        RECT  0.570 2.990 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.080 0.550 15.240 2.920 ;
        RECT  14.960 0.550 15.080 1.290 ;
        RECT  14.960 2.240 15.080 2.920 ;
        RECT  13.680 2.640 14.960 2.800 ;
        RECT  14.160 0.560 14.280 1.210 ;
        RECT  14.160 1.910 14.280 2.360 ;
        RECT  14.000 0.560 14.160 2.360 ;
        RECT  13.000 0.560 14.000 0.720 ;
        RECT  13.520 1.580 13.680 2.800 ;
        RECT  13.400 1.580 13.520 1.860 ;
        RECT  12.320 2.640 13.520 2.800 ;
        RECT  13.240 2.260 13.280 2.480 ;
        RECT  12.960 1.010 13.240 2.480 ;
        RECT  12.840 0.440 13.000 0.720 ;
        RECT  10.650 0.440 12.840 0.600 ;
        RECT  12.680 0.880 12.800 2.480 ;
        RECT  12.520 0.760 12.680 2.480 ;
        RECT  12.400 0.760 12.520 0.960 ;
        RECT  11.720 0.760 12.400 0.920 ;
        RECT  12.200 2.510 12.320 2.800 ;
        RECT  12.040 1.080 12.200 2.800 ;
        RECT  11.920 1.080 12.040 1.300 ;
        RECT  11.080 2.510 12.040 2.800 ;
        RECT  11.720 1.990 11.840 2.270 ;
        RECT  11.560 0.760 11.720 2.270 ;
        RECT  11.040 0.760 11.560 0.960 ;
        RECT  10.810 1.990 11.560 2.270 ;
        RECT  10.490 0.440 10.650 0.720 ;
        RECT  10.180 0.560 10.490 0.720 ;
        RECT  10.020 0.560 10.180 1.560 ;
        RECT  9.320 0.560 10.020 0.720 ;
        RECT  9.920 1.400 10.020 1.560 ;
        RECT  9.760 1.400 9.920 2.550 ;
        RECT  9.340 2.390 9.760 2.550 ;
        RECT  9.180 2.390 9.340 2.730 ;
        RECT  9.160 0.560 9.320 0.840 ;
        RECT  8.540 2.570 9.180 2.730 ;
        RECT  9.000 1.630 9.120 1.850 ;
        RECT  8.840 0.440 9.000 1.850 ;
        RECT  7.180 0.440 8.840 0.600 ;
        RECT  8.260 2.450 8.540 2.730 ;
        RECT  7.980 1.080 8.260 1.660 ;
        RECT  7.300 1.500 7.980 1.660 ;
        RECT  7.440 2.880 7.720 3.160 ;
        RECT  6.760 3.000 7.440 3.160 ;
        RECT  7.020 1.080 7.300 1.660 ;
        RECT  7.020 0.440 7.180 0.920 ;
        RECT  4.690 0.760 7.020 0.920 ;
        RECT  6.680 1.500 7.020 1.660 ;
        RECT  4.350 0.440 6.860 0.600 ;
        RECT  6.680 2.050 6.760 3.160 ;
        RECT  6.680 1.090 6.740 1.250 ;
        RECT  6.520 1.090 6.680 3.160 ;
        RECT  6.460 1.090 6.520 1.250 ;
        RECT  6.480 2.040 6.520 3.160 ;
        RECT  6.300 1.430 6.340 1.730 ;
        RECT  6.140 1.090 6.300 1.730 ;
        RECT  5.470 1.090 6.140 1.280 ;
        RECT  5.520 2.440 5.800 3.070 ;
        RECT  5.430 2.440 5.520 2.730 ;
        RECT  5.430 1.090 5.470 1.740 ;
        RECT  5.310 1.090 5.430 2.730 ;
        RECT  5.270 1.540 5.310 2.730 ;
        RECT  5.110 1.080 5.130 1.240 ;
        RECT  4.950 1.080 5.110 3.100 ;
        RECT  4.910 1.080 4.950 1.700 ;
        RECT  1.330 2.940 4.950 3.100 ;
        RECT  4.850 1.080 4.910 1.240 ;
        RECT  4.690 1.860 4.790 2.780 ;
        RECT  4.630 0.760 4.690 2.780 ;
        RECT  4.530 0.760 4.630 2.020 ;
        RECT  2.770 2.620 4.630 2.780 ;
        RECT  4.350 2.180 4.470 2.460 ;
        RECT  4.190 0.440 4.350 2.460 ;
        RECT  3.290 0.440 4.190 0.600 ;
        RECT  3.430 1.970 4.190 2.130 ;
        RECT  3.870 0.770 4.030 1.110 ;
        RECT  3.230 0.950 3.870 1.110 ;
        RECT  3.110 0.950 3.230 2.190 ;
        RECT  3.070 0.550 3.110 2.190 ;
        RECT  2.950 0.550 3.070 1.110 ;
        RECT  2.950 1.910 3.070 2.190 ;
        RECT  2.230 0.550 2.950 0.710 ;
        RECT  2.290 2.030 2.950 2.190 ;
        RECT  2.490 2.360 2.770 2.780 ;
        RECT  2.470 0.890 2.750 1.170 ;
        RECT  1.810 2.620 2.490 2.780 ;
        RECT  1.890 1.010 2.470 1.170 ;
        RECT  2.010 2.030 2.290 2.310 ;
        RECT  0.870 0.550 2.230 0.770 ;
        RECT  1.810 1.010 1.890 1.290 ;
        RECT  1.650 1.010 1.810 2.780 ;
        RECT  1.610 1.010 1.650 2.420 ;
        RECT  1.530 2.140 1.610 2.420 ;
        RECT  1.330 0.990 1.410 1.270 ;
        RECT  1.130 0.990 1.330 3.100 ;
        RECT  1.050 1.930 1.130 3.100 ;
        RECT  0.870 1.380 0.970 1.660 ;
        RECT  0.710 0.550 0.870 2.690 ;
        RECT  0.370 0.550 0.710 0.720 ;
        RECT  0.370 2.530 0.710 2.690 ;
        RECT  0.090 0.440 0.370 0.720 ;
        RECT  0.090 2.530 0.370 2.820 ;
    END
END AFHCINX4TR

MACRO AFHCINX2TR
    CLASS CORE ;
    FOREIGN AFHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.760 0.820 9.050 1.100 ;
        RECT  8.720 0.820 8.760 1.160 ;
        RECT  8.440 0.820 8.720 2.890 ;
        RECT  8.240 0.820 8.440 1.100 ;
        END
        ANTENNADIFFAREA 2.534 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.400 2.470 7.720 2.750 ;
        RECT  6.760 2.590 7.400 2.750 ;
        RECT  7.200 0.760 7.360 1.440 ;
        RECT  7.080 0.760 7.200 1.800 ;
        RECT  7.040 1.280 7.080 1.800 ;
        RECT  6.760 1.640 7.040 1.800 ;
        RECT  6.480 1.640 6.760 2.750 ;
        END
        ANTENNADIFFAREA 4.767 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.880 1.240 13.120 2.360 ;
        RECT  12.650 1.480 12.880 1.760 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.260 1.640 5.560 1.960 ;
        END
        ANTENNAGATEAREA 0.7464 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.240 0.720 1.640 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.110 -0.280 13.200 0.280 ;
        RECT  12.830 -0.280 13.110 1.080 ;
        RECT  11.490 -0.280 12.830 0.280 ;
        RECT  11.210 -0.280 11.490 0.340 ;
        RECT  8.850 -0.280 11.210 0.280 ;
        RECT  8.500 -0.280 8.850 0.340 ;
        RECT  5.800 -0.280 8.500 0.280 ;
        RECT  0.900 -0.280 5.800 0.340 ;
        RECT  0.620 -0.280 0.900 0.390 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.110 3.320 13.200 3.880 ;
        RECT  12.830 2.530 13.110 3.880 ;
        RECT  11.690 3.320 12.830 3.880 ;
        RECT  11.410 2.930 11.690 3.880 ;
        RECT  9.200 3.320 11.410 3.880 ;
        RECT  8.920 2.610 9.200 3.880 ;
        RECT  8.200 3.320 8.920 3.880 ;
        RECT  7.920 2.610 8.200 3.880 ;
        RECT  5.760 3.320 7.920 3.880 ;
        RECT  5.480 2.420 5.760 3.880 ;
        RECT  0.860 3.260 5.480 3.880 ;
        RECT  0.580 2.120 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.490 0.440 12.630 1.310 ;
        RECT  12.490 1.920 12.630 3.160 ;
        RECT  12.350 0.440 12.490 3.160 ;
        RECT  12.330 0.440 12.350 2.770 ;
        RECT  11.530 2.610 12.330 2.770 ;
        RECT  12.010 1.920 12.170 2.450 ;
        RECT  11.850 0.500 12.010 2.450 ;
        RECT  11.730 0.500 11.850 1.320 ;
        RECT  10.810 0.500 11.730 0.660 ;
        RECT  11.410 1.720 11.530 2.770 ;
        RECT  11.370 1.600 11.410 2.770 ;
        RECT  11.130 1.600 11.370 1.880 ;
        RECT  10.170 2.610 11.370 2.770 ;
        RECT  10.970 2.170 11.210 2.450 ;
        RECT  10.810 1.000 10.970 2.450 ;
        RECT  10.650 0.450 10.810 0.660 ;
        RECT  10.690 1.000 10.810 1.320 ;
        RECT  9.170 0.450 10.650 0.610 ;
        RECT  10.490 1.480 10.650 2.450 ;
        RECT  10.370 0.770 10.490 2.450 ;
        RECT  10.330 0.770 10.370 1.640 ;
        RECT  10.130 0.770 10.330 1.060 ;
        RECT  9.930 1.220 10.170 2.770 ;
        RECT  9.490 0.770 10.130 0.930 ;
        RECT  9.890 1.090 9.930 2.770 ;
        RECT  9.650 1.090 9.890 1.380 ;
        RECT  9.490 2.150 9.690 2.710 ;
        RECT  9.410 0.770 9.490 2.710 ;
        RECT  9.330 0.770 9.410 2.310 ;
        RECT  9.210 0.820 9.330 1.100 ;
        RECT  9.130 2.030 9.330 2.310 ;
        RECT  9.010 0.450 9.170 0.660 ;
        RECT  8.060 0.500 9.010 0.660 ;
        RECT  7.840 0.500 8.060 2.310 ;
        RECT  7.240 2.150 7.840 2.310 ;
        RECT  7.520 0.440 7.680 1.990 ;
        RECT  6.920 0.440 7.520 0.600 ;
        RECT  7.360 1.710 7.520 1.990 ;
        RECT  6.960 2.150 7.240 2.430 ;
        RECT  6.760 0.440 6.920 0.980 ;
        RECT  6.320 1.220 6.880 1.440 ;
        RECT  4.220 0.820 6.760 0.980 ;
        RECT  3.900 0.500 6.600 0.660 ;
        RECT  6.240 1.220 6.320 2.530 ;
        RECT  6.160 1.220 6.240 3.160 ;
        RECT  6.040 1.220 6.160 1.430 ;
        RECT  5.960 2.370 6.160 3.160 ;
        RECT  5.880 1.590 6.000 1.870 ;
        RECT  5.720 1.140 5.880 1.870 ;
        RECT  5.020 1.140 5.720 1.300 ;
        RECT  5.020 2.230 5.280 3.100 ;
        RECT  5.000 1.140 5.020 3.100 ;
        RECT  4.860 1.140 5.000 2.390 ;
        RECT  4.440 1.170 4.700 3.100 ;
        RECT  1.280 2.940 4.440 3.100 ;
        RECT  4.060 0.820 4.220 2.720 ;
        RECT  1.820 2.560 4.060 2.720 ;
        RECT  3.820 0.500 3.900 1.430 ;
        RECT  3.620 0.500 3.820 2.400 ;
        RECT  3.540 1.200 3.620 2.400 ;
        RECT  3.200 0.570 3.360 2.250 ;
        RECT  2.420 0.570 3.200 0.730 ;
        RECT  2.020 2.090 3.200 2.250 ;
        RECT  2.660 0.910 2.940 1.190 ;
        RECT  2.080 1.030 2.660 1.190 ;
        RECT  1.040 0.570 2.420 0.850 ;
        RECT  1.820 1.030 2.080 1.310 ;
        RECT  1.660 1.030 1.820 2.720 ;
        RECT  1.540 2.000 1.660 2.720 ;
        RECT  1.360 1.030 1.480 1.310 ;
        RECT  1.280 1.030 1.360 2.500 ;
        RECT  1.200 1.030 1.280 3.100 ;
        RECT  1.120 2.340 1.200 3.100 ;
        RECT  0.880 0.570 1.040 1.960 ;
        RECT  0.380 0.570 0.880 0.730 ;
        RECT  0.380 1.800 0.880 1.960 ;
        RECT  0.100 0.440 0.380 1.080 ;
        RECT  0.100 1.800 0.380 3.160 ;
    END
END AFHCINX2TR

MACRO AFCSIHCONX4TR
    CLASS CORE ;
    FOREIGN AFCSIHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.160 0.440 10.320 3.160 ;
        RECT  10.030 0.440 10.160 1.260 ;
        RECT  10.000 1.840 10.160 3.160 ;
        RECT  9.680 1.840 10.000 2.560 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.160 0.480 9.240 0.760 ;
        RECT  8.840 0.440 9.160 0.760 ;
        END
        ANTENNAGATEAREA 0.2976 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.710 1.810 0.990 ;
        RECT  0.850 0.830 1.530 0.990 ;
        RECT  0.880 1.910 1.170 3.160 ;
        RECT  0.320 1.910 0.880 2.070 ;
        RECT  0.570 0.710 0.850 0.990 ;
        RECT  0.320 0.830 0.570 0.990 ;
        RECT  0.080 0.830 0.320 2.070 ;
        END
        ANTENNADIFFAREA 4.896 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 2.110 3.710 2.390 ;
        RECT  3.010 0.990 3.250 1.220 ;
        RECT  2.850 0.990 3.010 2.390 ;
        RECT  2.720 1.840 2.850 2.390 ;
        RECT  2.480 1.840 2.720 2.560 ;
        RECT  2.390 1.840 2.480 2.390 ;
        END
        ANTENNADIFFAREA 5.553 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.770 1.350 3.890 1.630 ;
        RECT  3.610 0.620 3.770 1.630 ;
        RECT  2.610 0.620 3.610 0.780 ;
        RECT  2.450 0.620 2.610 1.480 ;
        RECT  2.210 1.320 2.450 1.480 ;
        RECT  1.810 1.320 2.210 1.600 ;
        RECT  1.650 1.150 1.810 1.480 ;
        RECT  0.760 1.150 1.650 1.310 ;
        RECT  0.480 1.150 0.760 1.560 ;
        END
        ANTENNAGATEAREA 1.1736 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.320 1.520 4.330 1.950 ;
        RECT  4.200 1.520 4.320 2.360 ;
        RECT  4.050 1.520 4.200 2.710 ;
        RECT  4.040 1.790 4.050 2.710 ;
        RECT  3.450 1.790 4.040 1.950 ;
        RECT  3.540 2.550 4.040 2.710 ;
        RECT  3.380 2.550 3.540 2.880 ;
        RECT  3.170 1.560 3.450 1.950 ;
        RECT  2.230 2.720 3.380 2.880 ;
        RECT  2.070 1.760 2.230 2.880 ;
        RECT  1.490 1.760 2.070 1.920 ;
        RECT  1.330 1.470 1.490 1.920 ;
        RECT  1.090 1.470 1.330 1.750 ;
        END
        ANTENNAGATEAREA 1.1328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 -0.280 10.400 0.280 ;
        RECT  9.550 -0.280 9.830 1.300 ;
        RECT  7.290 -0.280 9.550 0.280 ;
        RECT  7.010 -0.280 7.290 0.400 ;
        RECT  6.430 -0.280 7.010 0.280 ;
        RECT  6.210 -0.280 6.430 1.190 ;
        RECT  4.210 -0.280 6.210 0.280 ;
        RECT  3.930 -0.280 4.210 1.190 ;
        RECT  2.290 -0.280 3.930 0.280 ;
        RECT  2.010 -0.280 2.290 1.100 ;
        RECT  1.330 -0.280 2.010 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 3.320 10.400 3.880 ;
        RECT  9.610 2.930 9.830 3.880 ;
        RECT  7.190 3.260 9.610 3.880 ;
        RECT  6.910 3.170 7.190 3.880 ;
        RECT  6.370 3.320 6.910 3.880 ;
        RECT  6.090 2.960 6.370 3.880 ;
        RECT  4.230 3.320 6.090 3.880 ;
        RECT  3.950 2.920 4.230 3.880 ;
        RECT  3.190 3.320 3.950 3.880 ;
        RECT  2.910 3.170 3.190 3.880 ;
        RECT  1.910 3.260 2.910 3.880 ;
        RECT  1.690 2.080 1.910 3.880 ;
        RECT  0.370 3.320 1.690 3.880 ;
        RECT  0.090 2.230 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.720 1.470 10.000 1.680 ;
        RECT  9.450 1.520 9.720 1.680 ;
        RECT  9.290 1.520 9.450 3.100 ;
        RECT  9.130 1.030 9.310 1.310 ;
        RECT  8.190 2.940 9.290 3.100 ;
        RECT  8.970 1.030 9.130 2.190 ;
        RECT  8.850 1.510 8.970 2.190 ;
        RECT  8.770 1.510 8.850 1.790 ;
        RECT  8.610 0.920 8.770 1.200 ;
        RECT  8.610 1.950 8.670 2.780 ;
        RECT  8.450 0.600 8.610 2.780 ;
        RECT  7.370 0.600 8.450 0.760 ;
        RECT  8.190 0.920 8.290 1.200 ;
        RECT  8.030 0.920 8.190 3.100 ;
        RECT  8.010 0.920 8.030 1.200 ;
        RECT  7.910 2.180 8.030 2.890 ;
        RECT  7.750 0.920 7.810 1.200 ;
        RECT  7.590 0.920 7.750 3.100 ;
        RECT  7.530 0.920 7.590 1.200 ;
        RECT  7.430 2.180 7.590 3.100 ;
        RECT  7.370 1.360 7.430 1.640 ;
        RECT  7.270 0.600 7.370 1.640 ;
        RECT  7.210 0.600 7.270 2.800 ;
        RECT  7.110 1.360 7.210 2.800 ;
        RECT  5.030 2.580 7.110 2.800 ;
        RECT  6.890 0.910 6.990 1.190 ;
        RECT  6.610 0.910 6.890 2.420 ;
        RECT  5.410 2.260 6.610 2.420 ;
        RECT  6.050 1.350 6.170 1.630 ;
        RECT  5.890 0.440 6.050 1.630 ;
        RECT  4.710 0.440 5.890 0.600 ;
        RECT  5.730 1.820 5.850 2.100 ;
        RECT  5.570 0.910 5.730 2.100 ;
        RECT  5.450 0.910 5.570 1.190 ;
        RECT  5.190 1.500 5.410 2.420 ;
        RECT  5.030 0.910 5.210 1.190 ;
        RECT  4.870 0.910 5.030 2.800 ;
        RECT  4.550 0.440 4.710 2.890 ;
        RECT  4.430 0.440 4.550 1.190 ;
        RECT  4.490 1.850 4.550 2.890 ;
    END
END AFCSIHCONX4TR

MACRO AFCSIHCONX2TR
    CLASS CORE ;
    FOREIGN AFCSIHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 0.440 8.720 3.160 ;
        RECT  8.430 0.440 8.480 1.310 ;
        RECT  8.430 1.910 8.480 3.160 ;
        END
        ANTENNADIFFAREA 3.552 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.560 0.480 7.640 0.760 ;
        RECT  7.240 0.440 7.560 0.760 ;
        END
        ANTENNAGATEAREA 0.2976 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.800 1.170 3.160 ;
        RECT  0.240 1.800 0.880 1.960 ;
        RECT  0.570 0.750 0.850 1.030 ;
        RECT  0.240 0.870 0.570 1.030 ;
        RECT  0.080 0.870 0.240 1.960 ;
        END
        ANTENNADIFFAREA 3.376 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 2.030 2.320 2.950 ;
        RECT  1.490 2.030 1.870 2.190 ;
        RECT  1.490 1.090 1.670 1.310 ;
        RECT  1.330 1.090 1.490 2.190 ;
        END
        ANTENNADIFFAREA 2.832 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.270 2.310 1.550 ;
        RECT  1.990 1.270 2.030 1.430 ;
        RECT  1.830 0.770 1.990 1.430 ;
        RECT  1.170 0.770 1.830 0.930 ;
        RECT  1.010 0.770 1.170 1.350 ;
        RECT  0.760 1.190 1.010 1.350 ;
        RECT  0.480 1.190 0.760 1.560 ;
        RECT  0.400 1.190 0.480 1.470 ;
        END
        ANTENNAGATEAREA 0.7176 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.520 2.750 1.870 ;
        RECT  2.480 1.520 2.720 2.360 ;
        RECT  2.470 1.520 2.480 1.870 ;
        RECT  1.870 1.710 2.470 1.870 ;
        RECT  1.650 1.590 1.870 1.870 ;
        END
        ANTENNAGATEAREA 0.6768 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.230 -0.280 8.800 0.280 ;
        RECT  7.950 -0.280 8.230 1.310 ;
        RECT  5.710 -0.280 7.950 0.280 ;
        RECT  5.430 -0.280 5.710 0.400 ;
        RECT  4.850 -0.280 5.430 0.280 ;
        RECT  4.630 -0.280 4.850 1.190 ;
        RECT  2.510 -0.280 4.630 0.280 ;
        RECT  2.230 -0.280 2.510 1.110 ;
        RECT  1.330 -0.280 2.230 0.280 ;
        RECT  1.050 -0.280 1.330 0.610 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.230 3.320 8.800 3.880 ;
        RECT  8.010 1.910 8.230 3.880 ;
        RECT  5.590 3.260 8.010 3.880 ;
        RECT  5.310 3.170 5.590 3.880 ;
        RECT  4.790 3.320 5.310 3.880 ;
        RECT  4.510 2.960 4.790 3.880 ;
        RECT  2.700 3.320 4.510 3.880 ;
        RECT  2.480 2.610 2.700 3.880 ;
        RECT  1.670 3.260 2.480 3.880 ;
        RECT  1.390 2.350 1.670 3.880 ;
        RECT  0.370 3.320 1.390 3.880 ;
        RECT  0.090 2.120 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.160 1.470 8.320 1.750 ;
        RECT  7.850 1.590 8.160 1.750 ;
        RECT  7.690 1.590 7.850 3.100 ;
        RECT  7.530 1.030 7.710 1.310 ;
        RECT  6.590 2.940 7.690 3.100 ;
        RECT  7.370 1.030 7.530 2.190 ;
        RECT  7.250 1.510 7.370 2.190 ;
        RECT  7.130 1.510 7.250 1.790 ;
        RECT  6.970 0.920 7.190 1.200 ;
        RECT  6.970 1.950 7.070 2.780 ;
        RECT  6.810 0.600 6.970 2.780 ;
        RECT  5.790 0.600 6.810 0.760 ;
        RECT  6.590 0.920 6.650 1.200 ;
        RECT  6.430 0.920 6.590 3.100 ;
        RECT  6.310 2.180 6.430 2.890 ;
        RECT  6.150 0.920 6.230 1.200 ;
        RECT  5.990 0.920 6.150 3.100 ;
        RECT  5.950 0.920 5.990 1.200 ;
        RECT  5.830 2.180 5.990 3.100 ;
        RECT  5.790 1.360 5.830 1.640 ;
        RECT  5.670 0.600 5.790 1.640 ;
        RECT  5.630 0.600 5.670 2.800 ;
        RECT  5.510 1.360 5.630 2.800 ;
        RECT  3.450 2.580 5.510 2.800 ;
        RECT  5.290 0.910 5.410 1.190 ;
        RECT  5.010 0.910 5.290 2.420 ;
        RECT  3.830 2.260 5.010 2.420 ;
        RECT  4.470 1.350 4.590 1.630 ;
        RECT  4.310 0.440 4.470 1.630 ;
        RECT  3.130 0.440 4.310 0.600 ;
        RECT  4.150 1.820 4.270 2.100 ;
        RECT  3.990 0.910 4.150 2.100 ;
        RECT  3.870 0.910 3.990 1.190 ;
        RECT  3.610 1.500 3.830 2.420 ;
        RECT  3.450 0.910 3.630 1.190 ;
        RECT  3.290 0.910 3.450 2.800 ;
        RECT  2.970 0.440 3.130 2.890 ;
        RECT  2.850 0.440 2.970 1.190 ;
        RECT  2.910 1.850 2.970 2.890 ;
    END
END AFCSIHCONX2TR

MACRO AFCSHCONX4TR
    CLASS CORE ;
    FOREIGN AFCSHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  24.940 0.440 25.120 3.160 ;
        RECT  24.830 0.440 24.940 1.360 ;
        RECT  24.830 2.060 24.940 3.160 ;
        RECT  24.480 0.640 24.830 1.360 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  24.040 1.000 24.320 1.660 ;
        RECT  23.990 1.490 24.040 1.660 ;
        END
        ANTENNAGATEAREA 0.2928 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.760 1.480 16.910 1.700 ;
        RECT  16.150 2.380 16.440 2.660 ;
        RECT  15.490 2.380 16.150 2.540 ;
        RECT  14.760 2.380 15.490 2.660 ;
        RECT  14.440 1.480 14.760 2.660 ;
        END
        ANTENNADIFFAREA 6.599 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.640 2.980 14.480 3.140 ;
        RECT  12.480 2.280 12.640 3.140 ;
        RECT  12.360 2.280 12.480 2.440 ;
        RECT  12.040 1.400 12.360 2.440 ;
        RECT  11.900 2.280 12.040 2.440 ;
        RECT  11.680 2.280 11.900 2.560 ;
        END
        ANTENNADIFFAREA 7.18 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  19.230 1.580 20.360 1.960 ;
        END
        ANTENNAGATEAREA 0.8832 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.560 1.800 8.300 2.020 ;
        RECT  7.000 1.800 7.560 2.360 ;
        END
        ANTENNAGATEAREA 0.9576 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.240 4.720 1.560 ;
        RECT  4.010 1.280 4.440 1.560 ;
        END
        ANTENNAGATEAREA 0.7272 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.470 1.060 1.750 ;
        RECT  0.480 1.470 0.760 1.960 ;
        RECT  0.420 1.470 0.480 1.750 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  24.540 -0.280 25.200 0.280 ;
        RECT  24.260 -0.280 24.540 0.400 ;
        RECT  23.790 -0.280 24.260 0.280 ;
        RECT  23.510 -0.280 23.790 0.340 ;
        RECT  23.230 -0.280 23.510 0.280 ;
        RECT  22.950 -0.280 23.230 0.610 ;
        RECT  21.130 -0.280 22.950 0.280 ;
        RECT  20.850 -0.280 21.130 0.290 ;
        RECT  20.090 -0.280 20.850 0.280 ;
        RECT  19.810 -0.280 20.090 0.290 ;
        RECT  19.050 -0.280 19.810 0.280 ;
        RECT  18.770 -0.280 19.050 0.290 ;
        RECT  9.300 -0.280 18.770 0.280 ;
        RECT  9.020 -0.280 9.300 0.620 ;
        RECT  8.220 -0.280 9.020 0.280 ;
        RECT  7.940 -0.280 8.220 0.580 ;
        RECT  3.920 -0.280 7.940 0.340 ;
        RECT  1.740 -0.280 3.920 0.280 ;
        RECT  1.460 -0.280 1.740 0.360 ;
        RECT  0.860 -0.280 1.460 0.280 ;
        RECT  0.580 -0.280 0.860 1.310 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  24.590 3.320 25.200 3.880 ;
        RECT  24.310 2.800 24.590 3.880 ;
        RECT  24.030 3.320 24.310 3.880 ;
        RECT  23.750 2.670 24.030 3.880 ;
        RECT  21.150 3.320 23.750 3.880 ;
        RECT  20.870 1.990 21.150 3.880 ;
        RECT  20.210 3.320 20.870 3.880 ;
        RECT  19.930 2.870 20.210 3.880 ;
        RECT  19.190 3.320 19.930 3.880 ;
        RECT  18.910 3.200 19.190 3.880 ;
        RECT  9.700 3.320 18.910 3.880 ;
        RECT  9.420 3.050 9.700 3.880 ;
        RECT  8.460 3.260 9.420 3.880 ;
        RECT  7.700 3.320 8.460 3.880 ;
        RECT  7.420 3.260 7.700 3.880 ;
        RECT  6.580 3.320 7.420 3.880 ;
        RECT  5.100 3.260 6.580 3.880 ;
        RECT  4.380 3.320 5.100 3.880 ;
        RECT  1.850 3.260 4.380 3.880 ;
        RECT  1.570 3.180 1.850 3.880 ;
        RECT  0.860 3.320 1.570 3.880 ;
        RECT  0.580 2.960 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  24.660 1.520 24.720 1.800 ;
        RECT  24.500 1.520 24.660 2.510 ;
        RECT  23.590 2.350 24.500 2.510 ;
        RECT  23.760 1.910 24.070 2.190 ;
        RECT  23.760 1.000 23.880 1.280 ;
        RECT  23.600 1.000 23.760 2.190 ;
        RECT  23.270 2.030 23.600 2.190 ;
        RECT  23.430 2.350 23.590 3.060 ;
        RECT  22.070 2.900 23.430 3.060 ;
        RECT  23.270 1.380 23.390 1.660 ;
        RECT  23.110 0.770 23.270 1.660 ;
        RECT  23.110 2.030 23.270 2.740 ;
        RECT  22.550 0.770 23.110 0.930 ;
        RECT  22.510 2.580 23.110 2.740 ;
        RECT  22.670 1.090 22.950 2.420 ;
        RECT  22.430 1.090 22.670 1.310 ;
        RECT  22.390 0.450 22.550 0.930 ;
        RECT  22.230 1.470 22.510 2.740 ;
        RECT  17.150 0.450 22.390 0.610 ;
        RECT  22.070 0.880 22.230 1.160 ;
        RECT  21.850 0.880 22.070 3.060 ;
        RECT  21.530 0.880 21.690 3.000 ;
        RECT  21.410 0.880 21.530 1.160 ;
        RECT  21.370 1.990 21.530 3.000 ;
        RECT  21.250 1.360 21.370 1.640 ;
        RECT  21.090 0.770 21.250 1.640 ;
        RECT  18.150 0.770 21.090 0.930 ;
        RECT  20.530 1.090 20.690 3.090 ;
        RECT  20.330 1.090 20.530 1.310 ;
        RECT  20.410 2.120 20.530 3.090 ;
        RECT  19.390 2.540 20.410 2.700 ;
        RECT  19.070 2.120 19.730 2.380 ;
        RECT  19.070 1.090 19.570 1.310 ;
        RECT  19.230 2.540 19.390 2.950 ;
        RECT  17.230 2.790 19.230 2.950 ;
        RECT  18.910 1.090 19.070 2.630 ;
        RECT  18.750 1.540 18.910 1.820 ;
        RECT  17.790 2.470 18.910 2.630 ;
        RECT  18.590 2.030 18.750 2.310 ;
        RECT  18.430 1.090 18.590 2.310 ;
        RECT  18.310 1.090 18.430 1.310 ;
        RECT  18.150 2.030 18.270 2.310 ;
        RECT  17.990 0.770 18.150 2.310 ;
        RECT  17.790 0.770 17.990 1.050 ;
        RECT  17.630 2.350 17.790 2.630 ;
        RECT  17.470 1.000 17.630 2.630 ;
        RECT  17.310 1.000 17.470 1.280 ;
        RECT  17.070 1.940 17.230 2.950 ;
        RECT  16.990 0.450 17.150 1.320 ;
        RECT  16.520 1.940 17.070 2.140 ;
        RECT  14.280 1.160 16.990 1.320 ;
        RECT  16.610 0.440 16.830 0.770 ;
        RECT  14.090 0.440 16.610 0.600 ;
        RECT  16.150 1.900 16.520 2.140 ;
        RECT  13.630 0.840 16.430 1.000 ;
        RECT  15.340 1.900 16.150 2.060 ;
        RECT  15.020 1.900 15.340 2.180 ;
        RECT  14.120 1.160 14.280 2.820 ;
        RECT  12.960 2.660 14.120 2.820 ;
        RECT  13.840 0.440 14.090 0.660 ;
        RECT  13.280 2.280 13.960 2.500 ;
        RECT  13.470 0.440 13.630 1.000 ;
        RECT  9.620 0.440 13.470 0.600 ;
        RECT  13.120 0.760 13.280 2.500 ;
        RECT  9.940 0.760 13.120 0.920 ;
        RECT  12.800 1.080 12.960 2.820 ;
        RECT  10.780 1.080 12.800 1.240 ;
        RECT  12.100 2.610 12.320 3.160 ;
        RECT  11.520 3.000 12.100 3.160 ;
        RECT  11.700 1.400 11.840 1.620 ;
        RECT  11.540 1.400 11.700 1.940 ;
        RECT  11.520 1.780 11.540 1.940 ;
        RECT  11.360 1.780 11.520 3.160 ;
        RECT  11.140 1.400 11.380 1.620 ;
        RECT  10.020 3.000 11.360 3.160 ;
        RECT  11.140 2.560 11.200 2.840 ;
        RECT  10.980 1.400 11.140 2.840 ;
        RECT  10.340 2.680 10.980 2.840 ;
        RECT  10.580 1.080 10.780 2.520 ;
        RECT  10.500 2.300 10.580 2.520 ;
        RECT  10.260 1.080 10.380 1.300 ;
        RECT  10.180 2.400 10.340 2.840 ;
        RECT  10.100 1.080 10.260 2.180 ;
        RECT  9.780 2.400 10.180 2.570 ;
        RECT  9.940 1.900 10.100 2.180 ;
        RECT  9.860 2.730 10.020 3.160 ;
        RECT  9.780 0.760 9.940 1.260 ;
        RECT  9.780 1.460 9.940 1.740 ;
        RECT  9.260 2.730 9.860 2.890 ;
        RECT  9.460 1.100 9.780 1.260 ;
        RECT  9.620 1.460 9.780 2.570 ;
        RECT  9.460 0.440 9.620 0.940 ;
        RECT  8.940 2.410 9.620 2.570 ;
        RECT  7.600 0.780 9.460 0.940 ;
        RECT  9.300 1.100 9.460 2.250 ;
        RECT  7.540 1.100 9.300 1.320 ;
        RECT  8.620 2.090 9.300 2.250 ;
        RECT  9.100 2.730 9.260 3.100 ;
        RECT  8.860 1.480 9.140 1.930 ;
        RECT  2.170 2.940 9.100 3.100 ;
        RECT  8.780 2.410 8.940 2.780 ;
        RECT  7.280 1.480 8.860 1.640 ;
        RECT  6.840 2.620 8.780 2.780 ;
        RECT  8.460 2.090 8.620 2.460 ;
        RECT  7.940 2.240 8.460 2.460 ;
        RECT  7.440 0.540 7.600 0.940 ;
        RECT  5.040 0.540 7.440 0.700 ;
        RECT  7.120 0.860 7.280 1.640 ;
        RECT  5.520 0.860 7.120 1.020 ;
        RECT  6.840 1.180 6.960 1.390 ;
        RECT  6.680 1.180 6.840 2.780 ;
        RECT  5.690 1.180 6.680 1.340 ;
        RECT  5.970 1.500 6.130 2.380 ;
        RECT  5.520 1.500 5.970 1.660 ;
        RECT  5.930 2.220 5.970 2.380 ;
        RECT  5.640 2.220 5.930 2.500 ;
        RECT  5.360 1.840 5.700 2.060 ;
        RECT  5.360 0.860 5.520 1.660 ;
        RECT  5.240 0.860 5.360 1.210 ;
        RECT  5.200 1.840 5.360 2.700 ;
        RECT  2.850 2.540 5.200 2.700 ;
        RECT  4.880 0.540 5.040 2.290 ;
        RECT  4.320 0.800 4.880 1.080 ;
        RECT  4.620 2.010 4.880 2.290 ;
        RECT  3.720 2.060 3.860 2.340 ;
        RECT  3.680 1.230 3.720 2.340 ;
        RECT  3.560 0.440 3.680 2.340 ;
        RECT  3.400 0.440 3.560 1.750 ;
        RECT  3.330 1.470 3.400 1.750 ;
        RECT  3.170 2.150 3.370 2.380 ;
        RECT  3.170 0.520 3.220 1.210 ;
        RECT  3.010 0.520 3.170 2.380 ;
        RECT  3.000 0.520 3.010 1.220 ;
        RECT  1.380 0.520 3.000 0.680 ;
        RECT  2.740 2.130 2.850 2.780 ;
        RECT  2.550 0.840 2.740 2.780 ;
        RECT  2.520 0.840 2.550 1.130 ;
        RECT  2.140 0.840 2.310 2.370 ;
        RECT  2.010 2.630 2.170 3.100 ;
        RECT  1.980 0.840 2.140 1.120 ;
        RECT  2.090 2.060 2.140 2.370 ;
        RECT  0.380 2.630 2.010 2.790 ;
        RECT  1.490 1.280 1.940 1.560 ;
        RECT  1.380 1.280 1.490 2.330 ;
        RECT  1.220 0.520 1.380 2.330 ;
        RECT  1.060 1.030 1.220 1.310 ;
        RECT  1.060 2.050 1.220 2.330 ;
        RECT  0.260 0.470 0.380 1.310 ;
        RECT  0.320 2.630 0.380 3.160 ;
        RECT  0.260 1.910 0.320 3.160 ;
        RECT  0.100 0.470 0.260 3.160 ;
    END
END AFCSHCONX4TR

MACRO AFCSHCONX2TR
    CLASS CORE ;
    FOREIGN AFCSHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  22.940 0.440 23.120 3.160 ;
        RECT  22.830 0.440 22.940 1.310 ;
        RECT  22.830 1.940 22.940 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  22.270 0.840 22.360 1.160 ;
        RECT  22.040 0.840 22.270 1.760 ;
        RECT  21.990 1.480 22.040 1.760 ;
        END
        ANTENNAGATEAREA 0.2976 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.520 1.580 15.590 1.860 ;
        RECT  13.710 2.540 14.070 2.860 ;
        RECT  13.520 2.540 13.710 2.700 ;
        RECT  13.280 1.580 13.520 2.700 ;
        END
        ANTENNADIFFAREA 7.314 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.000 2.950 13.290 3.160 ;
        RECT  11.720 2.290 12.000 3.160 ;
        RECT  11.520 2.290 11.720 2.450 ;
        RECT  11.520 1.410 11.600 1.630 ;
        RECT  11.320 1.410 11.520 2.450 ;
        RECT  11.280 1.640 11.320 2.450 ;
        RECT  11.040 2.290 11.280 2.450 ;
        RECT  10.760 2.290 11.040 2.570 ;
        END
        ANTENNADIFFAREA 4.564 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  17.910 1.640 18.530 1.960 ;
        END
        ANTENNAGATEAREA 0.4896 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 1.760 7.560 2.360 ;
        RECT  7.070 1.760 7.240 2.100 ;
        END
        ANTENNAGATEAREA 0.528 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 1.230 5.120 1.650 ;
        END
        ANTENNAGATEAREA 0.7944 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.440 1.020 1.660 ;
        RECT  0.480 1.440 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  22.590 -0.280 23.200 0.280 ;
        RECT  22.310 -0.280 22.590 0.400 ;
        RECT  21.290 -0.280 22.310 0.340 ;
        RECT  21.010 -0.280 21.290 0.580 ;
        RECT  19.250 -0.280 21.010 0.280 ;
        RECT  18.970 -0.280 19.250 0.360 ;
        RECT  17.750 -0.280 18.970 0.280 ;
        RECT  17.470 -0.280 17.750 0.360 ;
        RECT  8.560 -0.280 17.470 0.280 ;
        RECT  8.280 -0.280 8.560 0.580 ;
        RECT  6.900 -0.280 8.280 0.280 ;
        RECT  6.120 -0.280 6.900 0.580 ;
        RECT  4.280 -0.280 6.120 0.340 ;
        RECT  1.680 -0.280 4.280 0.280 ;
        RECT  1.400 -0.280 1.680 0.340 ;
        RECT  0.860 -0.280 1.400 0.280 ;
        RECT  0.580 -0.280 0.860 1.220 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  22.590 3.320 23.200 3.880 ;
        RECT  22.310 2.800 22.590 3.880 ;
        RECT  22.030 3.320 22.310 3.880 ;
        RECT  21.750 2.700 22.030 3.880 ;
        RECT  19.290 3.320 21.750 3.880 ;
        RECT  19.010 2.040 19.290 3.880 ;
        RECT  17.830 3.320 19.010 3.880 ;
        RECT  17.550 3.200 17.830 3.880 ;
        RECT  8.760 3.320 17.550 3.880 ;
        RECT  8.480 3.020 8.760 3.880 ;
        RECT  7.620 3.320 8.480 3.880 ;
        RECT  7.340 3.260 7.620 3.880 ;
        RECT  6.820 3.320 7.340 3.880 ;
        RECT  5.500 3.260 6.820 3.880 ;
        RECT  4.500 3.320 5.500 3.880 ;
        RECT  4.220 3.260 4.500 3.880 ;
        RECT  1.900 3.320 4.220 3.880 ;
        RECT  1.590 2.800 1.900 3.880 ;
        RECT  0.860 3.320 1.590 3.880 ;
        RECT  0.580 2.800 0.860 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  22.660 1.500 22.780 1.780 ;
        RECT  22.500 1.500 22.660 2.540 ;
        RECT  21.590 2.380 22.500 2.540 ;
        RECT  21.760 1.940 22.070 2.220 ;
        RECT  21.760 1.010 21.880 1.290 ;
        RECT  21.600 1.010 21.760 2.220 ;
        RECT  21.270 2.060 21.600 2.220 ;
        RECT  21.430 2.380 21.590 3.090 ;
        RECT  20.190 2.930 21.430 3.090 ;
        RECT  21.270 1.450 21.390 1.730 ;
        RECT  21.110 0.790 21.270 1.730 ;
        RECT  21.110 2.060 21.270 2.770 ;
        RECT  20.610 0.790 21.110 0.950 ;
        RECT  20.570 2.610 21.110 2.770 ;
        RECT  20.730 1.110 20.950 2.450 ;
        RECT  20.480 1.110 20.730 1.330 ;
        RECT  20.450 0.520 20.610 0.950 ;
        RECT  20.350 1.500 20.570 2.770 ;
        RECT  16.330 0.520 20.450 0.680 ;
        RECT  20.190 0.910 20.290 1.190 ;
        RECT  19.970 0.910 20.190 3.090 ;
        RECT  19.650 0.910 19.810 3.060 ;
        RECT  19.530 0.910 19.650 1.190 ;
        RECT  19.490 2.040 19.650 3.060 ;
        RECT  19.370 1.490 19.490 1.770 ;
        RECT  19.210 0.840 19.370 1.770 ;
        RECT  16.830 0.840 19.210 1.000 ;
        RECT  18.690 1.160 18.850 3.160 ;
        RECT  18.450 1.160 18.690 1.440 ;
        RECT  18.530 2.120 18.690 3.160 ;
        RECT  15.590 2.860 18.530 3.020 ;
        RECT  18.070 2.420 18.350 2.700 ;
        RECT  17.750 1.160 18.270 1.440 ;
        RECT  17.750 2.540 18.070 2.700 ;
        RECT  17.590 1.160 17.750 2.700 ;
        RECT  17.450 1.490 17.590 1.770 ;
        RECT  16.470 2.540 17.590 2.700 ;
        RECT  17.290 2.100 17.430 2.380 ;
        RECT  17.130 1.160 17.290 2.380 ;
        RECT  17.010 1.160 17.130 1.440 ;
        RECT  16.830 2.100 16.950 2.380 ;
        RECT  16.670 0.840 16.830 2.380 ;
        RECT  16.490 0.840 16.670 1.120 ;
        RECT  16.330 2.420 16.470 2.700 ;
        RECT  16.170 0.520 16.330 0.980 ;
        RECT  16.170 1.140 16.330 2.700 ;
        RECT  15.850 0.820 16.170 0.980 ;
        RECT  16.010 1.140 16.170 1.420 ;
        RECT  13.600 0.440 16.010 0.660 ;
        RECT  15.690 0.820 15.850 1.420 ;
        RECT  13.090 1.260 15.690 1.420 ;
        RECT  15.430 2.020 15.590 3.020 ;
        RECT  13.080 0.880 15.530 1.100 ;
        RECT  14.760 2.020 15.430 2.380 ;
        RECT  13.770 2.100 14.760 2.380 ;
        RECT  13.310 0.440 13.600 0.720 ;
        RECT  12.930 1.260 13.090 2.790 ;
        RECT  12.920 0.440 13.080 1.100 ;
        RECT  12.320 2.630 12.930 2.790 ;
        RECT  8.880 0.440 12.920 0.600 ;
        RECT  12.660 2.190 12.770 2.470 ;
        RECT  12.490 0.760 12.660 2.470 ;
        RECT  11.800 0.760 12.490 0.930 ;
        RECT  12.160 1.090 12.320 2.790 ;
        RECT  10.120 1.090 12.160 1.250 ;
        RECT  9.200 0.760 11.800 0.920 ;
        RECT  11.240 2.610 11.520 2.980 ;
        RECT  10.600 2.820 11.240 2.980 ;
        RECT  10.960 1.410 11.120 1.630 ;
        RECT  10.800 1.410 10.960 2.010 ;
        RECT  10.600 1.850 10.800 2.010 ;
        RECT  10.280 1.410 10.640 1.690 ;
        RECT  10.440 1.850 10.600 2.980 ;
        RECT  9.080 2.820 10.440 2.980 ;
        RECT  10.120 1.410 10.280 2.660 ;
        RECT  9.960 1.080 10.120 1.250 ;
        RECT  10.000 2.380 10.120 2.660 ;
        RECT  8.840 2.380 10.000 2.540 ;
        RECT  9.800 1.080 9.960 2.220 ;
        RECT  9.480 2.000 9.800 2.220 ;
        RECT  9.520 1.080 9.640 1.300 ;
        RECT  9.360 1.080 9.520 1.540 ;
        RECT  9.320 1.380 9.360 1.540 ;
        RECT  9.160 1.380 9.320 2.220 ;
        RECT  9.040 0.760 9.200 1.220 ;
        RECT  9.000 2.000 9.160 2.220 ;
        RECT  8.920 2.700 9.080 2.980 ;
        RECT  8.520 1.060 9.040 1.220 ;
        RECT  8.200 2.700 8.920 2.860 ;
        RECT  8.720 0.440 8.880 0.900 ;
        RECT  8.680 1.670 8.840 2.540 ;
        RECT  8.120 0.740 8.720 0.900 ;
        RECT  7.880 2.380 8.680 2.540 ;
        RECT  8.360 1.060 8.520 2.220 ;
        RECT  7.800 1.060 8.360 1.280 ;
        RECT  7.900 2.060 8.360 2.220 ;
        RECT  7.980 1.440 8.200 1.860 ;
        RECT  8.040 2.700 8.200 3.100 ;
        RECT  7.960 0.440 8.120 0.900 ;
        RECT  2.390 2.940 8.040 3.100 ;
        RECT  7.220 1.440 7.980 1.600 ;
        RECT  7.320 0.440 7.960 0.600 ;
        RECT  7.720 2.380 7.880 2.680 ;
        RECT  7.640 0.910 7.800 1.280 ;
        RECT  6.780 2.520 7.720 2.680 ;
        RECT  7.140 0.440 7.320 0.900 ;
        RECT  7.060 1.060 7.220 1.600 ;
        RECT  6.140 0.740 7.140 0.900 ;
        RECT  6.460 1.060 7.060 1.220 ;
        RECT  6.780 1.380 6.900 1.660 ;
        RECT  6.620 1.380 6.780 2.680 ;
        RECT  6.300 1.060 6.460 2.470 ;
        RECT  6.020 2.300 6.300 2.580 ;
        RECT  5.980 0.740 6.140 2.130 ;
        RECT  4.440 2.300 6.020 2.460 ;
        RECT  5.440 1.970 5.980 2.130 ;
        RECT  5.600 0.530 5.820 1.000 ;
        RECT  4.440 0.530 5.600 0.690 ;
        RECT  5.280 0.850 5.440 2.130 ;
        RECT  3.580 2.620 5.370 2.780 ;
        RECT  4.620 0.850 5.280 1.070 ;
        RECT  4.700 1.970 5.280 2.130 ;
        RECT  4.280 0.530 4.440 2.460 ;
        RECT  3.760 0.440 3.920 2.210 ;
        RECT  3.160 0.500 3.760 0.660 ;
        RECT  3.420 0.950 3.580 2.780 ;
        RECT  2.780 2.620 3.420 2.780 ;
        RECT  3.100 0.890 3.260 2.330 ;
        RECT  3.000 0.890 3.100 1.160 ;
        RECT  2.840 0.500 3.000 1.160 ;
        RECT  1.380 0.500 2.840 0.660 ;
        RECT  2.620 1.380 2.780 2.780 ;
        RECT  2.460 0.900 2.620 1.570 ;
        RECT  2.230 2.480 2.390 3.100 ;
        RECT  2.240 1.910 2.300 2.190 ;
        RECT  2.080 0.820 2.240 2.190 ;
        RECT  0.380 2.480 2.230 2.640 ;
        RECT  1.920 0.820 2.080 1.100 ;
        RECT  1.380 1.340 1.920 1.620 ;
        RECT  1.220 0.500 1.380 2.130 ;
        RECT  1.060 0.940 1.220 1.220 ;
        RECT  1.060 1.970 1.220 2.130 ;
        RECT  0.260 0.480 0.380 1.220 ;
        RECT  0.320 2.480 0.380 3.080 ;
        RECT  0.260 1.910 0.320 3.080 ;
        RECT  0.100 0.480 0.260 3.080 ;
    END
END AFCSHCONX2TR

MACRO AFCSHCINX4TR
    CLASS CORE ;
    FOREIGN AFCSHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  24.040 0.550 24.300 3.160 ;
        RECT  23.660 0.640 24.040 1.370 ;
        END
        ANTENNADIFFAREA 3.499 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  23.260 1.510 23.520 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.990 0.760 17.150 2.390 ;
        RECT  16.830 0.760 16.990 1.040 ;
        RECT  16.090 0.760 16.830 0.920 ;
        RECT  15.820 0.760 16.090 2.830 ;
        RECT  15.810 1.440 15.820 2.830 ;
        RECT  15.680 1.440 15.810 2.160 ;
        RECT  15.190 1.440 15.680 1.720 ;
        RECT  15.160 1.440 15.190 2.560 ;
        RECT  14.900 1.200 15.160 2.560 ;
        END
        ANTENNADIFFAREA 8.221 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.320 2.670 13.600 2.830 ;
        RECT  12.320 1.080 13.140 1.240 ;
        RECT  12.080 1.080 12.320 2.830 ;
        RECT  10.840 1.080 12.080 1.240 ;
        RECT  11.070 2.280 12.080 2.440 ;
        END
        ANTENNADIFFAREA 10.1655 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  19.250 1.640 19.650 1.960 ;
        END
        ANTENNAGATEAREA 0.588 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.920 1.620 7.930 1.780 ;
        RECT  7.550 1.620 7.920 1.960 ;
        END
        ANTENNAGATEAREA 0.6456 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.290 1.630 ;
        END
        ANTENNAGATEAREA 0.7104 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.540 0.570 1.800 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2544 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  23.800 -0.280 24.400 0.280 ;
        RECT  23.440 -0.280 23.800 0.470 ;
        RECT  23.100 -0.280 23.440 0.280 ;
        RECT  22.940 -0.280 23.100 0.850 ;
        RECT  19.630 -0.280 22.940 0.280 ;
        RECT  18.940 -0.280 19.630 0.340 ;
        RECT  8.740 -0.280 18.940 0.280 ;
        RECT  8.060 -0.280 8.740 0.610 ;
        RECT  7.300 -0.280 8.060 0.280 ;
        RECT  7.020 -0.280 7.300 0.610 ;
        RECT  1.750 -0.280 7.020 0.280 ;
        RECT  1.470 -0.280 1.750 0.460 ;
        RECT  0.900 -0.280 1.470 0.280 ;
        RECT  0.610 -0.280 0.900 0.460 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  23.840 3.320 24.400 3.880 ;
        RECT  23.530 2.940 23.840 3.880 ;
        RECT  22.980 3.320 23.530 3.880 ;
        RECT  22.700 2.940 22.980 3.880 ;
        RECT  20.960 3.320 22.700 3.880 ;
        RECT  20.660 2.440 20.960 3.880 ;
        RECT  19.960 3.320 20.660 3.880 ;
        RECT  18.890 3.140 19.960 3.880 ;
        RECT  8.810 3.320 18.890 3.880 ;
        RECT  8.530 2.930 8.810 3.880 ;
        RECT  7.610 3.320 8.530 3.880 ;
        RECT  7.330 2.930 7.610 3.880 ;
        RECT  5.670 3.320 7.330 3.880 ;
        RECT  5.390 3.260 5.670 3.880 ;
        RECT  2.070 3.320 5.390 3.880 ;
        RECT  1.610 3.260 2.070 3.880 ;
        RECT  0.860 3.320 1.610 3.880 ;
        RECT  0.560 2.910 0.860 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  23.700 1.580 23.860 2.780 ;
        RECT  21.980 2.620 23.700 2.780 ;
        RECT  23.100 2.200 23.330 2.450 ;
        RECT  23.100 1.030 23.160 1.310 ;
        RECT  22.940 1.030 23.100 2.450 ;
        RECT  22.020 2.290 22.940 2.450 ;
        RECT  22.620 0.500 22.780 1.660 ;
        RECT  17.470 0.500 22.620 0.660 ;
        RECT  22.300 1.090 22.460 2.130 ;
        RECT  22.120 1.090 22.300 1.250 ;
        RECT  22.180 1.970 22.300 2.130 ;
        RECT  22.020 1.540 22.060 1.820 ;
        RECT  21.860 1.540 22.020 2.450 ;
        RECT  21.700 2.620 21.980 2.890 ;
        RECT  21.700 1.010 21.920 1.170 ;
        RECT  21.540 1.010 21.700 2.890 ;
        RECT  21.220 0.950 21.380 3.120 ;
        RECT  20.900 0.870 21.060 1.750 ;
        RECT  18.050 0.870 20.900 1.030 ;
        RECT  20.260 1.200 20.420 2.890 ;
        RECT  20.120 1.200 20.260 1.360 ;
        RECT  17.630 2.730 20.260 2.890 ;
        RECT  19.090 2.210 19.570 2.370 ;
        RECT  19.090 1.200 19.520 1.360 ;
        RECT  18.930 1.200 19.090 2.370 ;
        RECT  18.570 1.540 18.930 1.700 ;
        RECT  18.430 1.860 18.590 2.430 ;
        RECT  18.400 1.190 18.530 1.350 ;
        RECT  18.400 1.860 18.430 2.020 ;
        RECT  18.240 1.190 18.400 2.020 ;
        RECT  18.050 2.210 18.170 2.370 ;
        RECT  17.890 0.870 18.050 2.370 ;
        RECT  17.790 0.870 17.890 1.150 ;
        RECT  17.470 0.890 17.630 2.890 ;
        RECT  17.310 0.440 17.470 0.660 ;
        RECT  17.310 0.890 17.470 1.170 ;
        RECT  16.740 2.730 17.470 2.890 ;
        RECT  14.100 0.440 17.310 0.600 ;
        RECT  16.450 2.170 16.740 2.890 ;
        RECT  16.450 1.080 16.570 1.240 ;
        RECT  16.290 1.080 16.450 2.380 ;
        RECT  14.740 0.880 15.630 1.040 ;
        RECT  15.450 2.490 15.610 2.920 ;
        RECT  14.740 2.730 15.450 2.920 ;
        RECT  14.630 0.880 14.740 2.920 ;
        RECT  14.580 0.880 14.630 3.150 ;
        RECT  14.380 0.880 14.580 1.200 ;
        RECT  14.340 2.670 14.580 3.150 ;
        RECT  14.260 1.700 14.420 2.510 ;
        RECT  9.130 2.990 14.340 3.150 ;
        RECT  14.100 1.700 14.260 1.860 ;
        RECT  12.640 2.350 14.260 2.510 ;
        RECT  13.940 0.440 14.100 1.860 ;
        RECT  13.780 2.030 14.090 2.190 ;
        RECT  13.620 0.440 13.780 2.190 ;
        RECT  9.060 0.440 13.620 0.600 ;
        RECT  12.800 2.030 13.620 2.190 ;
        RECT  13.300 0.760 13.460 1.560 ;
        RECT  10.120 0.760 13.300 0.920 ;
        RECT  12.640 1.400 13.300 1.560 ;
        RECT  12.480 1.400 12.640 2.510 ;
        RECT  10.810 2.670 11.860 2.830 ;
        RECT  10.810 1.400 11.640 1.560 ;
        RECT  10.650 1.400 10.810 2.830 ;
        RECT  10.560 1.400 10.650 1.560 ;
        RECT  9.450 2.670 10.650 2.830 ;
        RECT  10.400 1.090 10.560 1.560 ;
        RECT  10.280 1.090 10.400 1.250 ;
        RECT  10.120 2.280 10.390 2.440 ;
        RECT  9.960 0.760 10.120 2.440 ;
        RECT  9.800 0.860 9.960 1.020 ;
        RECT  9.610 1.180 9.770 2.510 ;
        RECT  9.600 1.180 9.610 1.340 ;
        RECT  9.320 0.980 9.600 1.340 ;
        RECT  9.290 2.290 9.450 2.830 ;
        RECT  9.190 1.780 9.350 2.130 ;
        RECT  8.250 2.290 9.290 2.450 ;
        RECT  8.740 1.970 9.190 2.130 ;
        RECT  8.970 2.610 9.130 3.150 ;
        RECT  8.900 0.440 9.060 0.930 ;
        RECT  6.660 2.610 8.970 2.770 ;
        RECT  6.230 0.770 8.900 0.930 ;
        RECT  8.580 1.090 8.740 2.130 ;
        RECT  8.460 1.090 8.580 1.250 ;
        RECT  8.090 1.090 8.250 2.450 ;
        RECT  6.660 1.090 8.090 1.250 ;
        RECT  6.660 2.290 8.090 2.450 ;
        RECT  3.950 0.440 6.660 0.600 ;
        RECT  6.500 1.090 6.660 2.450 ;
        RECT  6.500 2.610 6.660 3.100 ;
        RECT  5.230 2.940 6.500 3.100 ;
        RECT  6.180 2.500 6.340 2.780 ;
        RECT  6.070 0.770 6.230 2.190 ;
        RECT  4.910 2.500 6.180 2.660 ;
        RECT  5.830 0.940 6.070 1.100 ;
        RECT  5.610 1.320 5.910 1.480 ;
        RECT  5.450 0.770 5.610 1.950 ;
        RECT  4.790 0.770 5.450 0.930 ;
        RECT  5.150 1.790 5.450 1.950 ;
        RECT  5.070 2.940 5.230 3.160 ;
        RECT  4.870 1.790 5.150 2.130 ;
        RECT  2.390 3.000 5.070 3.160 ;
        RECT  4.750 2.500 4.910 2.840 ;
        RECT  4.710 1.790 4.870 1.950 ;
        RECT  2.830 2.680 4.750 2.840 ;
        RECT  4.550 1.390 4.710 1.950 ;
        RECT  4.390 2.240 4.590 2.520 ;
        RECT  4.390 0.950 4.430 1.230 ;
        RECT  4.230 0.950 4.390 2.520 ;
        RECT  3.150 2.360 4.230 2.520 ;
        RECT  3.950 2.040 4.070 2.200 ;
        RECT  3.790 0.440 3.950 2.200 ;
        RECT  3.470 2.040 3.590 2.200 ;
        RECT  3.310 0.440 3.470 2.200 ;
        RECT  2.070 0.440 3.310 0.600 ;
        RECT  2.990 0.760 3.150 2.520 ;
        RECT  2.390 0.760 2.990 0.920 ;
        RECT  2.550 1.080 2.830 2.840 ;
        RECT  2.350 0.760 2.390 1.160 ;
        RECT  2.230 2.780 2.390 3.160 ;
        RECT  2.230 0.760 2.350 2.600 ;
        RECT  2.190 1.030 2.230 2.600 ;
        RECT  1.330 2.780 2.230 2.950 ;
        RECT  2.030 1.030 2.190 1.200 ;
        RECT  1.910 0.440 2.070 0.870 ;
        RECT  1.730 0.710 1.910 0.870 ;
        RECT  1.570 0.710 1.730 1.580 ;
        RECT  0.890 0.710 1.570 0.870 ;
        RECT  1.450 1.420 1.570 1.580 ;
        RECT  1.210 1.090 1.410 1.250 ;
        RECT  1.210 1.910 1.330 2.950 ;
        RECT  1.050 1.090 1.210 2.950 ;
        RECT  0.730 0.710 0.890 2.680 ;
        RECT  0.150 0.710 0.730 1.000 ;
        RECT  0.310 2.520 0.730 2.680 ;
        RECT  0.150 2.520 0.310 3.160 ;
    END
END AFCSHCINX4TR

MACRO AFCSHCINX2TR
    CLASS CORE ;
    FOREIGN AFCSHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.280 0.440 19.520 3.160 ;
        RECT  19.270 1.310 19.280 3.160 ;
        RECT  19.190 1.950 19.270 3.160 ;
        END
        ANTENNADIFFAREA 3.686 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  18.880 0.840 19.120 1.160 ;
        RECT  18.710 1.000 18.880 1.160 ;
        RECT  18.550 1.000 18.710 1.770 ;
        RECT  18.510 1.490 18.550 1.770 ;
        END
        ANTENNAGATEAREA 0.2904 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.570 0.910 12.730 2.360 ;
        RECT  12.500 1.850 12.570 2.360 ;
        RECT  12.250 1.850 12.500 2.700 ;
        END
        ANTENNADIFFAREA 3.72 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 1.080 10.720 2.840 ;
        RECT  10.370 1.080 10.470 1.570 ;
        END
        ANTENNADIFFAREA 5.499 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.120 1.720 15.510 1.960 ;
        RECT  14.710 1.640 15.120 1.960 ;
        END
        ANTENNAGATEAREA 0.3024 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.120 1.410 7.370 1.690 ;
        RECT  6.880 1.240 7.120 1.690 ;
        RECT  6.750 1.410 6.880 1.690 ;
        END
        ANTENNAGATEAREA 0.336 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.240 5.210 1.640 ;
        END
        ANTENNAGATEAREA 0.7416 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.370 0.630 1.630 ;
        RECT  0.320 0.840 0.350 1.630 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.970 -0.280 19.600 0.280 ;
        RECT  18.690 -0.280 18.970 0.650 ;
        RECT  18.350 -0.280 18.690 0.280 ;
        RECT  18.190 -0.280 18.350 0.870 ;
        RECT  8.610 -0.280 18.190 0.280 ;
        RECT  8.330 -0.280 8.610 0.610 ;
        RECT  5.510 -0.280 8.330 0.280 ;
        RECT  5.230 -0.280 5.510 0.300 ;
        RECT  1.770 -0.280 5.230 0.280 ;
        RECT  1.490 -0.280 1.770 0.340 ;
        RECT  0.910 -0.280 1.490 0.280 ;
        RECT  0.630 -0.280 0.910 0.340 ;
        RECT  0.000 -0.280 0.630 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.950 3.320 19.600 3.880 ;
        RECT  18.650 2.950 18.950 3.880 ;
        RECT  18.260 3.320 18.650 3.880 ;
        RECT  17.980 3.020 18.260 3.880 ;
        RECT  16.150 3.320 17.980 3.880 ;
        RECT  15.990 2.240 16.150 3.880 ;
        RECT  14.750 3.320 15.990 3.880 ;
        RECT  14.470 3.240 14.750 3.880 ;
        RECT  5.590 3.320 14.470 3.880 ;
        RECT  5.310 3.260 5.590 3.880 ;
        RECT  1.810 3.320 5.310 3.880 ;
        RECT  1.530 3.260 1.810 3.880 ;
        RECT  0.880 3.320 1.530 3.880 ;
        RECT  0.580 2.560 0.880 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  19.030 1.510 19.110 1.790 ;
        RECT  18.870 1.510 19.030 2.770 ;
        RECT  18.360 2.610 18.870 2.770 ;
        RECT  18.350 2.090 18.530 2.250 ;
        RECT  18.350 1.050 18.390 1.330 ;
        RECT  18.200 2.610 18.360 2.850 ;
        RECT  18.190 1.050 18.350 2.250 ;
        RECT  17.190 2.690 18.200 2.850 ;
        RECT  18.030 2.090 18.190 2.250 ;
        RECT  17.870 0.580 18.030 1.710 ;
        RECT  17.870 2.090 18.030 2.530 ;
        RECT  11.760 0.580 17.870 0.740 ;
        RECT  17.270 2.370 17.870 2.530 ;
        RECT  17.550 1.110 17.710 2.210 ;
        RECT  17.350 1.110 17.550 1.270 ;
        RECT  17.430 2.050 17.550 2.210 ;
        RECT  17.270 1.570 17.290 1.850 ;
        RECT  17.110 1.570 17.270 2.530 ;
        RECT  16.950 2.690 17.190 2.910 ;
        RECT  16.950 1.040 17.150 1.200 ;
        RECT  16.910 1.040 16.950 2.910 ;
        RECT  16.790 1.040 16.910 2.850 ;
        RECT  16.610 2.240 16.630 3.160 ;
        RECT  16.450 0.980 16.610 3.160 ;
        RECT  16.130 0.900 16.290 1.780 ;
        RECT  13.690 0.900 16.130 1.060 ;
        RECT  15.670 1.220 15.830 3.160 ;
        RECT  15.450 1.220 15.670 1.380 ;
        RECT  15.510 2.120 15.670 3.160 ;
        RECT  13.210 2.770 15.510 2.930 ;
        RECT  14.550 2.120 15.270 2.280 ;
        RECT  14.550 1.220 15.260 1.380 ;
        RECT  14.390 1.220 14.550 2.280 ;
        RECT  14.290 1.840 14.390 2.120 ;
        RECT  14.110 1.220 14.230 1.380 ;
        RECT  14.110 2.450 14.230 2.610 ;
        RECT  13.950 1.220 14.110 2.610 ;
        RECT  13.690 2.450 13.770 2.610 ;
        RECT  13.530 0.900 13.690 2.610 ;
        RECT  13.460 2.450 13.530 2.610 ;
        RECT  13.050 0.910 13.210 2.930 ;
        RECT  12.900 2.210 13.050 2.930 ;
        RECT  12.090 1.030 12.250 1.310 ;
        RECT  11.930 1.150 12.090 2.830 ;
        RECT  11.880 2.670 11.930 2.830 ;
        RECT  11.690 2.670 11.880 3.160 ;
        RECT  11.600 0.580 11.760 2.510 ;
        RECT  7.330 3.000 11.690 3.160 ;
        RECT  11.060 2.350 11.600 2.510 ;
        RECT  11.220 0.440 11.380 2.190 ;
        RECT  8.930 0.440 11.220 0.600 ;
        RECT  10.900 0.760 11.060 2.510 ;
        RECT  9.550 0.760 10.900 0.920 ;
        RECT  10.090 2.100 10.210 2.780 ;
        RECT  9.930 1.080 10.090 2.780 ;
        RECT  9.810 1.080 9.930 1.240 ;
        RECT  8.790 2.620 9.930 2.780 ;
        RECT  9.550 2.300 9.730 2.460 ;
        RECT  9.390 0.760 9.550 2.460 ;
        RECT  8.950 1.090 9.130 2.410 ;
        RECT  8.850 1.090 8.950 1.250 ;
        RECT  8.770 0.440 8.930 0.930 ;
        RECT  7.870 1.420 8.790 1.580 ;
        RECT  8.630 2.290 8.790 2.780 ;
        RECT  6.150 0.770 8.770 0.930 ;
        RECT  6.560 2.290 8.630 2.450 ;
        RECT  4.830 2.620 8.410 2.780 ;
        RECT  5.830 0.440 8.160 0.600 ;
        RECT  7.710 1.090 7.870 2.130 ;
        RECT  7.590 1.090 7.710 1.250 ;
        RECT  7.370 1.970 7.710 2.130 ;
        RECT  7.110 2.940 7.330 3.160 ;
        RECT  5.150 2.940 7.110 3.100 ;
        RECT  6.560 1.090 6.670 1.250 ;
        RECT  6.390 1.090 6.560 2.450 ;
        RECT  5.990 0.770 6.150 2.190 ;
        RECT  5.750 0.780 5.990 0.940 ;
        RECT  5.890 1.910 5.990 2.190 ;
        RECT  5.670 0.440 5.830 0.620 ;
        RECT  5.530 1.420 5.830 1.580 ;
        RECT  3.870 0.460 5.670 0.620 ;
        RECT  5.370 0.920 5.530 1.960 ;
        RECT  4.710 0.920 5.370 1.080 ;
        RECT  5.010 1.800 5.370 1.960 ;
        RECT  4.990 2.940 5.150 3.160 ;
        RECT  4.850 1.800 5.010 2.190 ;
        RECT  2.130 3.000 4.990 3.160 ;
        RECT  4.630 1.800 4.850 1.960 ;
        RECT  4.670 2.620 4.830 2.840 ;
        RECT  2.750 2.680 4.670 2.840 ;
        RECT  4.470 1.500 4.630 1.960 ;
        RECT  4.310 2.260 4.510 2.520 ;
        RECT  4.310 0.960 4.410 1.240 ;
        RECT  4.150 0.960 4.310 2.520 ;
        RECT  3.070 2.360 4.150 2.520 ;
        RECT  3.870 2.040 3.990 2.200 ;
        RECT  3.710 0.460 3.870 2.200 ;
        RECT  3.390 2.040 3.510 2.200 ;
        RECT  3.230 0.440 3.390 2.200 ;
        RECT  2.090 0.440 3.230 0.600 ;
        RECT  2.910 0.780 3.070 2.520 ;
        RECT  2.410 0.780 2.910 0.940 ;
        RECT  2.590 1.100 2.750 2.840 ;
        RECT  2.310 0.780 2.410 0.980 ;
        RECT  2.250 0.780 2.310 2.580 ;
        RECT  2.150 0.820 2.250 2.580 ;
        RECT  2.010 0.820 2.150 0.980 ;
        RECT  2.110 2.300 2.150 2.580 ;
        RECT  1.970 2.940 2.130 3.160 ;
        RECT  1.930 0.440 2.090 0.660 ;
        RECT  1.750 1.500 1.990 1.780 ;
        RECT  1.290 2.940 1.970 3.100 ;
        RECT  1.750 0.500 1.930 0.660 ;
        RECT  1.590 0.500 1.750 1.780 ;
        RECT  0.950 0.500 1.590 0.660 ;
        RECT  1.430 1.500 1.590 1.780 ;
        RECT  1.270 1.090 1.430 1.250 ;
        RECT  1.270 2.000 1.290 3.160 ;
        RECT  1.110 1.090 1.270 3.160 ;
        RECT  0.790 0.500 0.950 2.400 ;
        RECT  0.110 0.500 0.790 0.680 ;
        RECT  0.330 2.240 0.790 2.400 ;
        RECT  0.170 2.240 0.330 3.160 ;
    END
END AFCSHCINX2TR

MACRO ADDHXLTR
    CLASS CORE ;
    FOREIGN ADDHXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.990 0.500 3.120 1.160 ;
        RECT  2.990 1.720 3.050 2.660 ;
        RECT  2.890 0.500 2.990 2.660 ;
        RECT  2.830 0.500 2.890 1.880 ;
        RECT  2.310 2.500 2.890 2.660 ;
        RECT  1.770 0.500 2.830 0.720 ;
        RECT  2.050 2.340 2.310 2.660 ;
        END
        ANTENNADIFFAREA 2.478 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.440 4.720 1.560 ;
        RECT  4.640 2.060 4.700 2.340 ;
        RECT  4.480 0.440 4.640 2.340 ;
        RECT  4.430 2.060 4.480 2.340 ;
        END
        ANTENNADIFFAREA 1.188 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.660 1.640 3.920 1.960 ;
        RECT  3.370 1.800 3.660 1.960 ;
        RECT  3.210 1.800 3.370 2.980 ;
        RECT  2.070 2.820 3.210 2.980 ;
        RECT  2.150 1.260 2.350 2.180 ;
        RECT  1.890 2.020 2.150 2.180 ;
        RECT  1.890 2.820 2.070 3.100 ;
        RECT  1.730 2.020 1.890 3.100 ;
        END
        ANTENNAGATEAREA 0.228 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.190 3.520 1.560 ;
        RECT  3.150 1.340 3.280 1.560 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 -0.280 4.800 0.280 ;
        RECT  3.860 -0.280 4.140 0.700 ;
        RECT  3.530 -0.280 3.860 0.280 ;
        RECT  3.250 -0.280 3.530 0.400 ;
        RECT  0.460 -0.280 3.250 0.280 ;
        RECT  0.180 -0.280 0.460 0.340 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 3.320 4.800 3.880 ;
        RECT  4.030 3.200 4.310 3.880 ;
        RECT  3.190 3.260 4.030 3.880 ;
        RECT  2.910 3.200 3.190 3.880 ;
        RECT  0.980 3.260 2.910 3.880 ;
        RECT  0.700 3.200 0.980 3.880 ;
        RECT  0.000 3.320 0.700 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.240 1.000 4.320 1.560 ;
        RECT  4.080 1.000 4.240 2.280 ;
        RECT  4.070 1.000 4.080 1.160 ;
        RECT  3.750 2.120 4.080 2.280 ;
        RECT  3.790 0.880 4.070 1.160 ;
        RECT  3.530 2.120 3.750 2.400 ;
        RECT  2.670 2.060 2.730 2.340 ;
        RECT  2.510 0.880 2.670 2.340 ;
        RECT  1.990 0.880 2.510 1.100 ;
        RECT  1.830 0.880 1.990 1.860 ;
        RECT  1.010 1.700 1.830 1.860 ;
        RECT  1.450 0.910 1.670 1.540 ;
        RECT  1.290 2.690 1.570 2.990 ;
        RECT  1.240 0.450 1.530 0.730 ;
        RECT  0.630 0.910 1.450 1.190 ;
        RECT  1.140 2.020 1.420 2.530 ;
        RECT  0.310 2.690 1.290 2.850 ;
        RECT  0.310 0.570 1.240 0.730 ;
        RECT  0.630 2.020 1.140 2.180 ;
        RECT  0.790 1.580 1.010 1.860 ;
        RECT  0.470 0.910 0.630 2.180 ;
        RECT  0.090 0.570 0.310 2.850 ;
    END
END ADDHXLTR

MACRO ADDHX4TR
    CLASS CORE ;
    FOREIGN ADDHX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.720 0.500 7.960 0.780 ;
        RECT  7.280 1.840 7.520 2.720 ;
        RECT  7.160 1.960 7.280 2.720 ;
        RECT  6.480 1.960 7.160 2.120 ;
        RECT  6.040 0.500 6.720 0.660 ;
        RECT  6.210 1.960 6.480 2.840 ;
        RECT  6.160 1.960 6.210 2.280 ;
        RECT  5.520 2.120 6.160 2.280 ;
        RECT  5.760 0.500 6.040 1.480 ;
        RECT  5.080 1.320 5.760 1.480 ;
        RECT  5.240 2.120 5.520 2.400 ;
        RECT  4.560 2.120 5.240 2.280 ;
        RECT  4.800 1.030 5.080 1.480 ;
        RECT  4.120 1.320 4.800 1.480 ;
        RECT  4.280 2.120 4.560 2.400 ;
        RECT  3.600 2.120 4.280 2.280 ;
        RECT  3.840 1.000 4.120 1.480 ;
        RECT  3.060 1.320 3.840 1.480 ;
        RECT  3.320 2.120 3.600 2.400 ;
        RECT  3.060 2.120 3.320 2.280 ;
        RECT  2.900 1.320 3.060 2.280 ;
        END
        ANTENNADIFFAREA 18.168 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.880 0.830 13.120 2.430 ;
        RECT  12.340 0.830 12.880 1.070 ;
        RECT  12.340 2.190 12.880 2.430 ;
        RECT  12.060 0.580 12.340 1.070 ;
        RECT  12.060 2.190 12.340 3.000 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 1.380 7.560 1.600 ;
        RECT  6.830 1.380 7.040 1.800 ;
        RECT  3.560 1.640 6.830 1.800 ;
        RECT  3.240 1.640 3.560 1.960 ;
        RECT  3.220 1.640 3.240 1.920 ;
        END
        ANTENNAGATEAREA 1.6656 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.160 1.490 10.760 1.770 ;
        RECT  8.640 1.240 9.160 1.770 ;
        END
        ANTENNAGATEAREA 1.6344 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.820 -0.280 13.200 0.280 ;
        RECT  12.540 -0.280 12.820 0.630 ;
        RECT  11.860 -0.280 12.540 0.280 ;
        RECT  11.580 -0.280 11.860 0.690 ;
        RECT  11.040 -0.280 11.580 0.280 ;
        RECT  10.760 -0.280 11.040 1.010 ;
        RECT  10.080 -0.280 10.760 0.280 ;
        RECT  9.800 -0.280 10.080 1.010 ;
        RECT  9.120 -0.280 9.800 0.280 ;
        RECT  8.840 -0.280 9.120 0.670 ;
        RECT  1.340 -0.280 8.840 0.280 ;
        RECT  1.060 -0.280 1.340 0.900 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 0.880 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.820 3.320 13.200 3.880 ;
        RECT  12.540 2.710 12.820 3.880 ;
        RECT  11.860 3.320 12.540 3.880 ;
        RECT  11.580 2.250 11.860 3.880 ;
        RECT  10.900 3.320 11.580 3.880 ;
        RECT  10.620 2.690 10.900 3.880 ;
        RECT  9.940 3.320 10.620 3.880 ;
        RECT  9.660 2.570 9.940 3.880 ;
        RECT  8.940 3.320 9.660 3.880 ;
        RECT  8.660 3.200 8.940 3.880 ;
        RECT  7.900 3.260 8.660 3.880 ;
        RECT  7.620 3.200 7.900 3.880 ;
        RECT  3.140 3.320 7.620 3.880 ;
        RECT  2.860 3.200 3.140 3.880 ;
        RECT  2.340 3.260 2.860 3.880 ;
        RECT  2.060 3.200 2.340 3.880 ;
        RECT  1.340 3.320 2.060 3.880 ;
        RECT  1.060 2.250 1.340 3.880 ;
        RECT  0.380 3.320 1.060 3.880 ;
        RECT  0.100 2.250 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.560 1.230 12.720 2.030 ;
        RECT  11.520 1.230 12.560 1.390 ;
        RECT  11.400 1.870 12.560 2.030 ;
        RECT  11.080 1.550 12.400 1.710 ;
        RECT  11.240 1.050 11.520 1.390 ;
        RECT  11.240 1.870 11.400 3.050 ;
        RECT  11.230 1.170 11.240 1.390 ;
        RECT  11.100 2.250 11.240 3.050 ;
        RECT  10.560 1.170 11.230 1.330 ;
        RECT  10.420 2.250 11.100 2.410 ;
        RECT  10.920 1.550 11.080 2.090 ;
        RECT  8.420 1.930 10.920 2.090 ;
        RECT  10.280 0.440 10.560 1.330 ;
        RECT  10.140 2.250 10.420 3.090 ;
        RECT  9.600 1.170 10.280 1.330 ;
        RECT  9.460 2.250 10.140 2.410 ;
        RECT  9.330 1.030 9.600 1.330 ;
        RECT  9.180 2.250 9.460 3.040 ;
        RECT  9.320 1.030 9.330 1.310 ;
        RECT  7.880 2.880 9.180 3.040 ;
        RECT  8.320 1.930 8.420 2.720 ;
        RECT  8.140 1.030 8.320 2.720 ;
        RECT  8.040 1.030 8.140 2.090 ;
        RECT  7.720 1.060 7.880 3.040 ;
        RECT  7.480 1.060 7.720 1.220 ;
        RECT  6.960 2.880 7.720 3.040 ;
        RECT  7.200 0.940 7.480 1.220 ;
        RECT  6.520 1.060 7.200 1.220 ;
        RECT  6.680 2.280 6.960 3.160 ;
        RECT  6.000 3.000 6.680 3.160 ;
        RECT  6.240 0.940 6.520 1.220 ;
        RECT  5.720 2.560 6.000 3.160 ;
        RECT  2.140 2.560 5.720 2.720 ;
        RECT  5.280 0.500 5.560 1.160 ;
        RECT  4.600 0.500 5.280 0.660 ;
        RECT  4.760 2.880 5.040 3.160 ;
        RECT  4.080 2.880 4.760 3.040 ;
        RECT  4.320 0.500 4.600 1.160 ;
        RECT  1.820 0.500 4.320 0.660 ;
        RECT  3.800 2.880 4.080 3.160 ;
        RECT  1.820 2.880 3.800 3.040 ;
        RECT  2.740 0.880 3.680 1.160 ;
        RECT  2.580 0.880 2.740 2.190 ;
        RECT  2.460 1.910 2.580 2.190 ;
        RECT  2.020 1.610 2.140 2.720 ;
        RECT  1.980 1.490 2.020 2.720 ;
        RECT  0.400 1.490 1.980 1.770 ;
        RECT  1.540 0.500 1.820 1.330 ;
        RECT  1.540 1.930 1.820 3.040 ;
        RECT  0.860 1.170 1.540 1.330 ;
        RECT  0.860 1.930 1.540 2.090 ;
        RECT  0.580 0.440 0.860 1.330 ;
        RECT  0.580 1.930 0.860 3.160 ;
        RECT  0.240 1.170 0.580 1.330 ;
        RECT  0.240 1.930 0.580 2.090 ;
        RECT  0.080 1.170 0.240 2.090 ;
    END
END ADDHX4TR

MACRO ADDHX2TR
    CLASS CORE ;
    FOREIGN ADDHX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 0.800 4.420 1.080 ;
        RECT  4.120 1.800 4.400 2.720 ;
        RECT  3.520 0.920 4.200 1.080 ;
        RECT  3.520 1.800 4.120 1.960 ;
        RECT  3.240 0.440 3.520 1.080 ;
        RECT  3.320 1.640 3.520 1.960 ;
        RECT  3.040 1.640 3.320 2.720 ;
        RECT  2.560 0.920 3.240 1.080 ;
        RECT  2.440 2.060 3.040 2.220 ;
        RECT  2.440 0.800 2.560 1.080 ;
        RECT  2.280 0.800 2.440 2.220 ;
        RECT  2.040 1.940 2.280 2.220 ;
        END
        ANTENNADIFFAREA 11.744 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.150 0.440 8.320 3.160 ;
        RECT  8.030 0.440 8.150 1.270 ;
        RECT  8.030 1.950 8.150 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.240 4.400 1.630 ;
        RECT  2.880 1.240 3.680 1.400 ;
        RECT  2.600 1.240 2.880 1.890 ;
        END
        ANTENNAGATEAREA 0.8448 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.560 1.580 7.040 1.860 ;
        RECT  5.280 1.240 5.560 1.860 ;
        END
        ANTENNAGATEAREA 0.8592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.830 -0.280 8.400 0.280 ;
        RECT  7.550 -0.280 7.830 1.180 ;
        RECT  6.840 -0.280 7.550 0.280 ;
        RECT  6.560 -0.280 6.840 1.100 ;
        RECT  5.840 -0.280 6.560 0.280 ;
        RECT  5.560 -0.280 5.840 0.340 ;
        RECT  1.340 -0.280 5.560 0.280 ;
        RECT  1.060 -0.280 1.340 1.100 ;
        RECT  0.380 -0.280 1.060 0.280 ;
        RECT  0.100 -0.280 0.380 1.280 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.830 3.320 8.400 3.880 ;
        RECT  7.550 1.910 7.830 3.880 ;
        RECT  6.840 3.320 7.550 3.880 ;
        RECT  6.560 2.820 6.840 3.880 ;
        RECT  5.840 3.320 6.560 3.880 ;
        RECT  5.560 3.200 5.840 3.880 ;
        RECT  4.980 3.260 5.560 3.880 ;
        RECT  4.700 3.200 4.980 3.880 ;
        RECT  1.380 3.320 4.700 3.880 ;
        RECT  1.100 3.200 1.380 3.880 ;
        RECT  0.380 3.320 1.100 3.880 ;
        RECT  0.100 2.910 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.710 1.470 7.920 1.750 ;
        RECT  7.360 1.590 7.710 1.750 ;
        RECT  7.200 1.590 7.360 2.180 ;
        RECT  7.040 0.530 7.320 1.420 ;
        RECT  7.040 2.340 7.320 3.100 ;
        RECT  5.380 2.020 7.200 2.180 ;
        RECT  6.360 1.260 7.040 1.420 ;
        RECT  6.360 2.340 7.040 2.500 ;
        RECT  6.080 0.500 6.360 1.420 ;
        RECT  6.080 2.340 6.360 3.040 ;
        RECT  4.740 0.500 6.080 0.660 ;
        RECT  4.740 2.880 6.080 3.040 ;
        RECT  5.120 2.020 5.380 2.300 ;
        RECT  5.100 1.000 5.120 2.300 ;
        RECT  4.900 1.000 5.100 2.180 ;
        RECT  4.580 0.480 4.740 3.040 ;
        RECT  4.000 0.480 4.580 0.640 ;
        RECT  3.800 2.880 4.580 3.040 ;
        RECT  3.720 0.480 4.000 0.760 ;
        RECT  3.520 2.270 3.800 3.040 ;
        RECT  0.700 2.880 3.520 3.040 ;
        RECT  2.760 0.480 3.040 0.760 ;
        RECT  1.340 2.380 2.800 2.660 ;
        RECT  1.660 0.480 2.760 0.640 ;
        RECT  1.820 0.810 2.100 1.740 ;
        RECT  1.780 1.580 1.820 1.740 ;
        RECT  1.620 1.580 1.780 2.160 ;
        RECT  1.500 0.480 1.660 1.420 ;
        RECT  1.500 1.880 1.620 2.160 ;
        RECT  1.340 1.260 1.500 1.420 ;
        RECT  1.180 1.260 1.340 2.660 ;
        RECT  0.860 1.260 1.180 1.420 ;
        RECT  0.580 2.020 1.180 2.300 ;
        RECT  0.420 1.580 1.020 1.860 ;
        RECT  0.580 0.440 0.860 1.420 ;
        RECT  0.540 2.460 0.700 3.040 ;
        RECT  0.420 2.460 0.540 2.620 ;
        RECT  0.260 1.580 0.420 2.620 ;
    END
END ADDHX2TR

MACRO ADDHX1TR
    CLASS CORE ;
    FOREIGN ADDHX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.140 1.000 3.300 2.010 ;
        RECT  2.720 1.000 3.140 1.160 ;
        RECT  2.380 1.850 3.140 2.010 ;
        RECT  2.400 0.840 2.720 1.160 ;
        RECT  2.100 1.850 2.380 2.250 ;
        END
        ANTENNADIFFAREA 3.888 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.030 4.720 2.190 ;
        RECT  4.430 1.030 4.440 1.310 ;
        RECT  4.430 1.910 4.440 2.190 ;
        END
        ANTENNADIFFAREA 1.688 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 2.550 4.470 2.770 ;
        RECT  3.020 2.550 3.180 3.100 ;
        RECT  2.220 2.940 3.020 3.100 ;
        RECT  2.700 1.360 2.980 1.690 ;
        RECT  1.920 1.530 2.700 1.690 ;
        RECT  2.060 2.410 2.220 3.100 ;
        RECT  1.920 2.410 2.060 2.570 ;
        RECT  1.760 1.530 1.920 2.570 ;
        RECT  1.640 1.530 1.760 1.960 ;
        RECT  1.320 1.620 1.640 1.900 ;
        END
        ANTENNAGATEAREA 0.4248 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.860 1.640 3.920 1.960 ;
        RECT  3.640 1.520 3.860 1.960 ;
        RECT  3.580 1.520 3.640 1.800 ;
        END
        ANTENNAGATEAREA 0.4296 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 -0.280 5.200 0.280 ;
        RECT  4.830 -0.280 5.110 0.400 ;
        RECT  3.620 -0.280 4.830 0.280 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  0.920 -0.280 3.340 0.280 ;
        RECT  0.640 -0.280 0.920 0.400 ;
        RECT  0.000 -0.280 0.640 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.950 3.320 5.200 3.880 ;
        RECT  4.600 3.260 4.950 3.880 ;
        RECT  3.620 3.320 4.600 3.880 ;
        RECT  3.340 3.200 3.620 3.880 ;
        RECT  0.920 3.260 3.340 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.040 1.580 5.100 1.860 ;
        RECT  4.880 0.560 5.040 3.090 ;
        RECT  4.650 0.560 4.880 0.720 ;
        RECT  4.230 2.930 4.880 3.090 ;
        RECT  4.370 0.450 4.650 0.720 ;
        RECT  4.080 0.960 4.240 2.390 ;
        RECT  3.950 2.930 4.230 3.150 ;
        RECT  4.020 0.960 4.080 1.240 ;
        RECT  2.860 2.170 4.080 2.390 ;
        RECT  3.860 0.640 4.020 1.240 ;
        RECT  3.100 0.640 3.860 0.800 ;
        RECT  2.880 0.520 3.100 0.800 ;
        RECT  2.240 0.520 2.880 0.680 ;
        RECT  2.580 2.170 2.860 2.780 ;
        RECT  2.080 0.520 2.240 1.370 ;
        RECT  1.160 1.210 2.080 1.370 ;
        RECT  1.700 0.440 1.920 0.720 ;
        RECT  0.720 0.890 1.920 1.050 ;
        RECT  1.620 2.820 1.900 3.100 ;
        RECT  0.400 0.560 1.700 0.720 ;
        RECT  0.400 2.820 1.620 3.040 ;
        RECT  1.130 2.250 1.430 2.530 ;
        RECT  0.880 1.210 1.160 1.860 ;
        RECT  0.720 2.250 1.130 2.410 ;
        RECT  0.560 0.890 0.720 2.410 ;
        RECT  0.120 0.560 0.400 3.040 ;
    END
END ADDHX1TR

MACRO ADDFHXLTR
    CLASS CORE ;
    FOREIGN ADDFHXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.630 0.840 9.920 2.190 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.920 1.640 9.150 1.960 ;
        RECT  8.760 1.030 8.920 2.190 ;
        RECT  8.680 1.030 8.760 1.310 ;
        END
        ANTENNADIFFAREA 1.16 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 1.240 8.320 1.830 ;
        END
        ANTENNAGATEAREA 0.0576 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.580 4.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2688 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.330 0.580 1.610 ;
        RECT  0.360 0.840 0.380 1.610 ;
        RECT  0.080 0.840 0.360 1.960 ;
        END
        ANTENNAGATEAREA 0.1152 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.340 -0.280 10.000 0.280 ;
        RECT  9.060 -0.280 9.340 0.760 ;
        RECT  8.100 -0.280 9.060 0.280 ;
        RECT  7.820 -0.280 8.100 0.340 ;
        RECT  5.080 -0.280 7.820 0.280 ;
        RECT  4.800 -0.280 5.080 0.290 ;
        RECT  1.850 -0.280 4.800 0.280 ;
        RECT  0.680 -0.280 1.850 0.340 ;
        RECT  0.000 -0.280 0.680 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.500 3.320 10.000 3.880 ;
        RECT  9.220 3.260 9.500 3.880 ;
        RECT  8.020 3.320 9.220 3.880 ;
        RECT  7.670 3.260 8.020 3.880 ;
        RECT  4.460 3.320 7.670 3.880 ;
        RECT  4.300 2.740 4.460 3.880 ;
        RECT  1.450 3.320 4.300 3.880 ;
        RECT  0.750 2.700 1.450 3.880 ;
        RECT  0.000 3.320 0.750 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.490 2.380 9.650 2.680 ;
        RECT  7.000 2.520 9.490 2.680 ;
        RECT  6.100 2.840 9.170 3.000 ;
        RECT  8.480 0.520 8.760 0.800 ;
        RECT  7.920 2.200 8.520 2.360 ;
        RECT  7.920 0.520 8.480 0.680 ;
        RECT  7.760 0.520 7.920 2.360 ;
        RECT  6.640 0.520 7.760 0.680 ;
        RECT  7.680 1.600 7.760 2.360 ;
        RECT  7.440 0.880 7.600 1.440 ;
        RECT  7.280 1.280 7.440 2.360 ;
        RECT  7.160 2.200 7.280 2.360 ;
        RECT  7.000 0.840 7.120 1.120 ;
        RECT  6.960 0.840 7.000 2.680 ;
        RECT  6.840 0.960 6.960 2.680 ;
        RECT  6.680 2.200 6.840 2.360 ;
        RECT  6.480 0.520 6.640 1.120 ;
        RECT  6.320 0.960 6.480 2.420 ;
        RECT  6.160 0.440 6.320 0.720 ;
        RECT  6.260 2.140 6.320 2.420 ;
        RECT  5.360 0.450 6.160 0.720 ;
        RECT  6.100 0.880 6.160 1.160 ;
        RECT  5.940 0.880 6.100 3.000 ;
        RECT  5.500 2.740 5.940 3.000 ;
        RECT  5.620 0.880 5.780 2.580 ;
        RECT  5.520 0.880 5.620 1.160 ;
        RECT  5.250 2.420 5.620 2.580 ;
        RECT  5.360 1.320 5.460 2.260 ;
        RECT  5.300 0.450 5.360 2.260 ;
        RECT  5.200 0.450 5.300 1.480 ;
        RECT  5.180 2.100 5.300 2.260 ;
        RECT  4.980 2.420 5.250 2.700 ;
        RECT  3.680 0.450 5.200 0.610 ;
        RECT  5.040 1.640 5.140 1.920 ;
        RECT  4.880 0.770 5.040 1.920 ;
        RECT  4.320 2.420 4.980 2.580 ;
        RECT  4.000 0.770 4.880 0.930 ;
        RECT  4.320 1.090 4.440 1.250 ;
        RECT  4.160 1.090 4.320 2.120 ;
        RECT  4.160 2.280 4.320 2.580 ;
        RECT  4.000 1.960 4.160 2.120 ;
        RECT  3.840 0.770 4.000 1.800 ;
        RECT  3.840 1.960 4.000 3.160 ;
        RECT  3.680 1.640 3.840 1.800 ;
        RECT  2.080 3.000 3.840 3.160 ;
        RECT  3.520 0.450 3.680 1.480 ;
        RECT  3.520 1.640 3.680 2.840 ;
        RECT  3.360 1.320 3.520 1.480 ;
        RECT  2.560 2.680 3.520 2.840 ;
        RECT  3.200 1.320 3.360 2.520 ;
        RECT  3.040 1.000 3.260 1.160 ;
        RECT  2.880 0.660 3.040 1.900 ;
        RECT  0.960 0.660 2.880 0.820 ;
        RECT  2.720 1.740 2.880 2.520 ;
        RECT  2.560 0.980 2.720 1.580 ;
        RECT  2.400 1.420 2.560 2.840 ;
        RECT  2.240 2.520 2.400 2.840 ;
        RECT  2.080 0.980 2.240 1.260 ;
        RECT  1.920 1.100 2.080 3.160 ;
        RECT  1.700 2.380 1.920 2.690 ;
        RECT  1.340 1.450 1.660 1.610 ;
        RECT  1.180 0.990 1.340 2.420 ;
        RECT  0.800 0.520 0.960 2.280 ;
        RECT  0.400 0.520 0.800 0.680 ;
        RECT  0.340 2.120 0.800 2.280 ;
        RECT  0.120 0.460 0.400 0.680 ;
        RECT  0.180 2.120 0.340 2.340 ;
    END
END ADDFHXLTR

MACRO ADDFHX4TR
    CLASS CORE ;
    FOREIGN ADDFHX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  22.640 1.440 22.720 2.160 ;
        RECT  22.560 1.440 22.640 3.160 ;
        RECT  22.320 0.440 22.560 3.160 ;
        RECT  22.280 0.440 22.320 1.320 ;
        END
        ANTENNADIFFAREA 4.38 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  21.280 0.440 21.600 2.200 ;
        END
        ANTENNADIFFAREA 3.942 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  19.680 1.240 20.040 1.760 ;
        END
        ANTENNAGATEAREA 0.5304 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.590 1.580 11.390 1.960 ;
        END
        ANTENNAGATEAREA 2.2032 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.240 1.530 1.630 ;
        END
        ANTENNAGATEAREA 0.9216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  23.080 -0.280 23.200 0.280 ;
        RECT  22.800 -0.280 23.080 1.080 ;
        RECT  22.080 -0.280 22.800 0.280 ;
        RECT  21.800 -0.280 22.080 1.320 ;
        RECT  21.120 -0.280 21.800 0.280 ;
        RECT  20.840 -0.280 21.120 1.320 ;
        RECT  20.080 -0.280 20.840 0.280 ;
        RECT  19.800 -0.280 20.080 0.670 ;
        RECT  18.620 -0.280 19.800 0.280 ;
        RECT  18.340 -0.280 18.620 0.320 ;
        RECT  12.510 -0.280 18.340 0.280 ;
        RECT  12.230 -0.280 12.510 0.340 ;
        RECT  11.550 -0.280 12.230 0.280 ;
        RECT  11.270 -0.280 11.550 0.340 ;
        RECT  0.850 -0.280 11.270 0.280 ;
        RECT  0.570 -0.280 0.850 1.080 ;
        RECT  0.000 -0.280 0.570 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  23.080 3.320 23.200 3.880 ;
        RECT  22.800 2.440 23.080 3.880 ;
        RECT  22.080 3.320 22.800 3.880 ;
        RECT  21.800 2.920 22.080 3.880 ;
        RECT  21.120 3.320 21.800 3.880 ;
        RECT  20.900 2.920 21.120 3.880 ;
        RECT  19.980 3.320 20.900 3.880 ;
        RECT  19.700 3.260 19.980 3.880 ;
        RECT  18.480 3.320 19.700 3.880 ;
        RECT  11.990 3.260 18.480 3.880 ;
        RECT  11.710 2.440 11.990 3.880 ;
        RECT  11.030 3.320 11.710 3.880 ;
        RECT  10.750 2.440 11.030 3.880 ;
        RECT  3.590 3.320 10.750 3.880 ;
        RECT  3.310 2.180 3.590 3.880 ;
        RECT  2.630 3.260 3.310 3.880 ;
        RECT  2.350 2.670 2.630 3.880 ;
        RECT  1.810 3.320 2.350 3.880 ;
        RECT  1.530 2.270 1.810 3.880 ;
        RECT  0.850 3.320 1.530 3.880 ;
        RECT  0.570 2.320 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  22.100 1.480 22.160 1.880 ;
        RECT  21.920 1.480 22.100 2.720 ;
        RECT  16.600 2.500 21.920 2.720 ;
        RECT  14.830 2.880 20.680 3.100 ;
        RECT  20.280 0.440 20.560 1.320 ;
        RECT  20.220 1.920 20.500 2.200 ;
        RECT  19.600 0.830 20.280 0.990 ;
        RECT  19.460 1.920 20.220 2.080 ;
        RECT  19.570 0.480 19.600 0.990 ;
        RECT  19.460 0.480 19.570 1.080 ;
        RECT  19.300 0.480 19.460 2.200 ;
        RECT  15.740 0.480 19.300 0.700 ;
        RECT  19.180 1.620 19.300 2.200 ;
        RECT  18.720 1.620 19.180 1.780 ;
        RECT  18.860 1.010 19.140 1.290 ;
        RECT  17.000 2.060 19.000 2.340 ;
        RECT  18.100 1.010 18.860 1.170 ;
        RECT  17.960 1.620 18.720 1.900 ;
        RECT  17.980 1.010 18.100 1.290 ;
        RECT  17.820 1.010 17.980 1.460 ;
        RECT  17.000 1.240 17.820 1.460 ;
        RECT  16.600 0.860 17.620 1.080 ;
        RECT  16.780 1.240 17.000 2.340 ;
        RECT  16.440 0.860 16.600 2.720 ;
        RECT  16.280 0.860 16.440 1.020 ;
        RECT  15.510 2.500 16.440 2.720 ;
        RECT  16.000 0.860 16.280 1.140 ;
        RECT  16.030 2.060 16.250 2.340 ;
        RECT  15.680 2.180 16.030 2.340 ;
        RECT  15.680 0.480 15.740 1.200 ;
        RECT  15.520 0.480 15.680 2.340 ;
        RECT  14.880 0.480 15.520 0.640 ;
        RECT  15.310 2.180 15.520 2.340 ;
        RECT  15.040 1.010 15.320 1.360 ;
        RECT  15.030 2.180 15.310 2.550 ;
        RECT  13.830 1.200 15.040 1.360 ;
        RECT  14.350 2.270 15.030 2.430 ;
        RECT  14.720 0.480 14.880 1.040 ;
        RECT  14.550 2.610 14.830 3.100 ;
        RECT  14.560 0.820 14.720 1.040 ;
        RECT  12.870 0.440 14.560 0.660 ;
        RECT  13.830 2.940 14.550 3.100 ;
        RECT  13.390 0.820 14.350 1.040 ;
        RECT  14.070 2.270 14.350 2.550 ;
        RECT  13.670 1.200 13.830 3.100 ;
        RECT  13.550 1.200 13.670 1.420 ;
        RECT  13.550 2.610 13.670 3.100 ;
        RECT  12.950 2.660 13.550 2.820 ;
        RECT  13.390 2.130 13.510 2.410 ;
        RECT  13.230 0.820 13.390 2.410 ;
        RECT  13.030 0.820 13.230 1.040 ;
        RECT  12.470 2.220 13.230 2.380 ;
        RECT  12.870 1.200 13.070 2.060 ;
        RECT  12.670 2.540 12.950 2.820 ;
        RECT  12.790 0.440 12.870 2.060 ;
        RECT  12.710 0.440 12.790 1.360 ;
        RECT  9.950 0.500 12.710 0.660 ;
        RECT  12.510 1.520 12.630 1.740 ;
        RECT  12.350 0.820 12.510 1.740 ;
        RECT  12.350 2.220 12.470 3.030 ;
        RECT  8.990 0.820 12.350 0.980 ;
        RECT  12.190 2.120 12.350 3.030 ;
        RECT  11.950 2.120 12.190 2.280 ;
        RECT  11.710 1.140 11.950 2.280 ;
        RECT  10.750 1.140 11.710 1.420 ;
        RECT  11.510 2.120 11.710 2.280 ;
        RECT  11.230 2.120 11.510 3.160 ;
        RECT  10.550 2.120 11.230 2.280 ;
        RECT  10.430 2.120 10.550 3.160 ;
        RECT  10.010 1.140 10.470 1.400 ;
        RECT  10.270 1.560 10.430 3.160 ;
        RECT  10.170 1.560 10.270 1.810 ;
        RECT  9.850 1.140 10.010 3.160 ;
        RECT  8.670 0.440 9.950 0.660 ;
        RECT  9.150 1.140 9.850 1.420 ;
        RECT  5.030 2.940 9.850 3.160 ;
        RECT  9.530 1.580 9.690 2.780 ;
        RECT  8.990 1.580 9.530 1.740 ;
        RECT  6.470 2.620 9.530 2.780 ;
        RECT  9.150 2.180 9.370 2.460 ;
        RECT  8.670 2.300 9.150 2.460 ;
        RECT  8.830 0.820 8.990 1.740 ;
        RECT  8.390 0.440 8.670 2.460 ;
        RECT  7.710 0.440 8.390 0.600 ;
        RECT  8.190 2.180 8.390 2.460 ;
        RECT  7.950 0.880 8.190 1.160 ;
        RECT  7.150 2.240 8.190 2.460 ;
        RECT  7.790 0.880 7.950 2.080 ;
        RECT  7.230 0.880 7.790 1.040 ;
        RECT  6.990 1.860 7.790 2.080 ;
        RECT  7.430 0.440 7.710 0.720 ;
        RECT  7.230 1.220 7.510 1.500 ;
        RECT  7.110 0.760 7.230 1.040 ;
        RECT  6.670 1.340 7.230 1.500 ;
        RECT  6.950 0.440 7.110 1.040 ;
        RECT  6.830 1.860 6.990 2.460 ;
        RECT  6.270 0.440 6.950 0.600 ;
        RECT  6.670 2.180 6.830 2.460 ;
        RECT  6.470 0.780 6.750 1.060 ;
        RECT  6.510 1.340 6.670 2.020 ;
        RECT  5.990 2.180 6.670 2.340 ;
        RECT  6.390 1.740 6.510 2.020 ;
        RECT  5.790 0.900 6.470 1.060 ;
        RECT  6.190 2.500 6.470 2.780 ;
        RECT  5.990 0.440 6.270 0.720 ;
        RECT  5.510 2.620 6.190 2.780 ;
        RECT  5.950 1.220 6.070 1.500 ;
        RECT  1.330 0.440 5.990 0.600 ;
        RECT  5.710 2.180 5.990 2.460 ;
        RECT  5.790 1.220 5.950 1.910 ;
        RECT  5.630 0.780 5.790 1.060 ;
        RECT  5.230 1.750 5.790 1.910 ;
        RECT  5.470 0.780 5.630 1.300 ;
        RECT  5.350 2.190 5.510 2.780 ;
        RECT  4.670 1.080 5.470 1.300 ;
        RECT  5.230 2.190 5.350 2.470 ;
        RECT  4.270 0.760 5.310 0.920 ;
        RECT  4.950 1.750 5.230 2.030 ;
        RECT  4.670 2.190 5.230 2.350 ;
        RECT  4.750 2.510 5.030 3.160 ;
        RECT  4.110 3.000 4.750 3.160 ;
        RECT  4.550 1.080 4.670 2.350 ;
        RECT  4.510 1.080 4.550 2.840 ;
        RECT  4.270 2.100 4.510 2.840 ;
        RECT  4.110 0.760 4.270 1.040 ;
        RECT  3.990 0.760 4.110 3.160 ;
        RECT  3.950 0.880 3.990 3.160 ;
        RECT  3.230 0.880 3.950 1.040 ;
        RECT  3.790 1.800 3.950 2.890 ;
        RECT  2.370 1.360 3.790 1.640 ;
        RECT  3.110 1.800 3.790 2.020 ;
        RECT  2.950 0.760 3.230 1.040 ;
        RECT  2.830 1.800 3.110 2.950 ;
        RECT  2.210 0.870 2.370 2.330 ;
        RECT  2.090 0.870 2.210 1.300 ;
        RECT  2.010 1.910 2.210 2.330 ;
        RECT  1.690 0.920 1.850 2.110 ;
        RECT  1.330 0.920 1.690 1.080 ;
        RECT  1.330 1.950 1.690 2.110 ;
        RECT  1.050 0.440 1.330 1.080 ;
        RECT  1.050 1.950 1.330 2.990 ;
        RECT  0.370 1.950 1.050 2.110 ;
        RECT  0.310 0.440 0.370 1.080 ;
        RECT  0.310 1.910 0.370 2.990 ;
        RECT  0.150 0.440 0.310 2.990 ;
        RECT  0.090 0.440 0.150 1.080 ;
        RECT  0.100 1.910 0.150 2.990 ;
    END
END ADDFHX4TR

MACRO ADDFHX2TR
    CLASS CORE ;
    FOREIGN ADDFHX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.480 0.440 14.720 3.160 ;
        END
        ANTENNADIFFAREA 3.74 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.760 2.040 13.920 2.360 ;
        RECT  13.600 0.440 13.760 2.360 ;
        RECT  13.440 0.440 13.600 1.140 ;
        RECT  13.440 1.910 13.600 2.360 ;
        END
        ANTENNADIFFAREA 3.499 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.740 1.580 13.120 1.960 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.410 1.620 9.030 2.010 ;
        END
        ANTENNAGATEAREA 1.0944 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.240 0.940 1.630 ;
        END
        ANTENNAGATEAREA 0.4752 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.200 -0.280 14.800 0.280 ;
        RECT  13.920 -0.280 14.200 1.270 ;
        RECT  12.720 -0.280 13.920 0.280 ;
        RECT  12.440 -0.280 12.720 0.360 ;
        RECT  0.380 -0.280 12.440 0.280 ;
        RECT  0.090 -0.280 0.380 0.910 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.200 3.320 14.800 3.880 ;
        RECT  13.920 2.910 14.200 3.880 ;
        RECT  12.640 3.320 13.920 3.880 ;
        RECT  12.360 3.260 12.640 3.880 ;
        RECT  8.950 3.320 12.360 3.880 ;
        RECT  8.670 2.490 8.950 3.880 ;
        RECT  2.610 3.320 8.670 3.880 ;
        RECT  2.330 2.780 2.610 3.880 ;
        RECT  1.370 3.320 2.330 3.880 ;
        RECT  1.090 2.880 1.370 3.880 ;
        RECT  0.370 3.320 1.090 3.880 ;
        RECT  0.090 1.920 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  14.100 1.580 14.320 2.720 ;
        RECT  11.600 2.560 14.100 2.720 ;
        RECT  10.680 2.880 13.400 3.100 ;
        RECT  12.960 0.570 13.240 1.320 ;
        RECT  12.880 2.120 13.160 2.400 ;
        RECT  12.490 0.760 12.960 0.920 ;
        RECT  12.490 2.120 12.880 2.280 ;
        RECT  12.330 0.760 12.490 2.280 ;
        RECT  11.240 0.760 12.330 0.920 ;
        RECT  12.180 1.760 12.330 2.040 ;
        RECT  12.080 1.090 12.170 1.320 ;
        RECT  11.980 1.090 12.080 1.600 ;
        RECT  11.920 1.090 11.980 2.370 ;
        RECT  11.820 1.440 11.920 2.370 ;
        RECT  11.600 1.080 11.720 1.300 ;
        RECT  11.440 1.080 11.600 2.720 ;
        RECT  11.280 2.440 11.440 2.720 ;
        RECT  11.080 0.760 11.240 1.540 ;
        RECT  11.020 0.960 11.080 1.540 ;
        RECT  10.960 0.960 11.020 2.570 ;
        RECT  10.700 0.440 10.980 0.610 ;
        RECT  10.860 1.380 10.960 2.570 ;
        RECT  9.800 0.450 10.700 0.610 ;
        RECT  10.520 0.940 10.680 3.100 ;
        RECT  10.120 2.740 10.520 3.100 ;
        RECT  10.200 0.850 10.360 2.490 ;
        RECT  9.960 0.850 10.200 1.130 ;
        RECT  9.770 2.330 10.200 2.490 ;
        RECT  9.880 1.290 10.040 2.150 ;
        RECT  9.800 1.290 9.880 1.450 ;
        RECT  9.820 1.990 9.880 2.150 ;
        RECT  9.640 0.450 9.800 1.450 ;
        RECT  9.570 2.330 9.770 3.150 ;
        RECT  7.110 0.450 9.640 0.610 ;
        RECT  9.410 1.610 9.640 1.890 ;
        RECT  9.400 2.170 9.570 3.150 ;
        RECT  9.250 0.770 9.410 1.890 ;
        RECT  8.350 2.170 9.400 2.330 ;
        RECT  7.430 0.770 9.250 0.930 ;
        RECT  8.250 1.090 9.000 1.310 ;
        RECT  8.250 2.170 8.350 3.150 ;
        RECT  8.030 1.090 8.250 3.150 ;
        RECT  7.710 1.090 7.870 3.160 ;
        RECT  7.590 1.090 7.710 1.310 ;
        RECT  4.050 3.000 7.710 3.160 ;
        RECT  7.430 1.470 7.550 2.840 ;
        RECT  7.390 0.770 7.430 2.840 ;
        RECT  7.270 0.770 7.390 1.630 ;
        RECT  4.990 2.680 7.390 2.840 ;
        RECT  7.110 2.240 7.230 2.520 ;
        RECT  6.950 0.450 7.110 2.520 ;
        RECT  6.310 0.450 6.950 0.610 ;
        RECT  5.670 2.300 6.950 2.520 ;
        RECT  6.510 0.980 6.790 1.760 ;
        RECT  6.470 1.600 6.510 1.760 ;
        RECT  6.190 1.600 6.470 2.140 ;
        RECT  6.150 0.450 6.310 0.990 ;
        RECT  5.670 1.600 6.190 1.760 ;
        RECT  6.030 0.710 6.150 0.990 ;
        RECT  5.670 0.710 5.830 0.990 ;
        RECT  5.510 0.440 5.670 1.760 ;
        RECT  4.870 0.440 5.510 0.600 ;
        RECT  5.470 1.600 5.510 1.760 ;
        RECT  5.190 1.600 5.470 2.200 ;
        RECT  5.230 0.980 5.350 1.260 ;
        RECT  5.070 0.980 5.230 1.360 ;
        RECT  4.510 1.600 5.190 1.760 ;
        RECT  3.890 1.200 5.070 1.360 ;
        RECT  4.710 1.920 4.990 2.840 ;
        RECT  4.590 0.440 4.870 0.990 ;
        RECT  3.770 2.360 4.710 2.520 ;
        RECT  0.850 0.440 4.590 0.600 ;
        RECT  4.350 1.600 4.510 2.200 ;
        RECT  4.130 0.760 4.410 1.040 ;
        RECT  4.230 1.920 4.350 2.200 ;
        RECT  3.370 0.760 4.130 0.920 ;
        RECT  3.770 2.780 4.050 3.160 ;
        RECT  3.770 1.080 3.890 1.360 ;
        RECT  3.610 1.080 3.770 2.520 ;
        RECT  3.130 3.000 3.770 3.160 ;
        RECT  3.290 2.240 3.610 2.520 ;
        RECT  3.130 0.760 3.370 1.040 ;
        RECT  2.970 0.760 3.130 3.160 ;
        RECT  2.330 0.760 2.970 0.920 ;
        RECT  2.810 2.240 2.970 3.160 ;
        RECT  2.130 1.220 2.810 1.500 ;
        RECT  2.130 2.360 2.810 2.520 ;
        RECT  2.050 0.760 2.330 1.040 ;
        RECT  1.770 1.220 2.130 1.380 ;
        RECT  1.970 2.360 2.130 3.060 ;
        RECT  1.850 2.780 1.970 3.060 ;
        RECT  1.610 0.820 1.770 2.190 ;
        RECT  1.490 0.820 1.610 1.150 ;
        RECT  1.490 1.910 1.610 2.190 ;
        RECT  1.170 0.920 1.330 2.110 ;
        RECT  0.850 0.920 1.170 1.080 ;
        RECT  0.850 1.950 1.170 2.110 ;
        RECT  0.570 0.440 0.850 1.080 ;
        RECT  0.570 1.950 0.850 2.690 ;
    END
END ADDFHX2TR

MACRO ADDFHX1TR
    CLASS CORE ;
    FOREIGN ADDFHX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.630 1.030 9.920 2.360 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.910 1.240 9.120 1.560 ;
        RECT  8.750 1.030 8.910 2.190 ;
        END
        ANTENNADIFFAREA 1.652 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.020 1.240 8.230 1.940 ;
        RECT  7.680 1.240 8.020 1.560 ;
        END
        ANTENNAGATEAREA 0.1488 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 1.080 4.720 1.560 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.540 2.360 ;
        END
        ANTENNAGATEAREA 0.2328 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.370 -0.280 10.000 0.280 ;
        RECT  9.090 -0.280 9.370 0.340 ;
        RECT  8.080 -0.280 9.090 0.280 ;
        RECT  7.800 -0.280 8.080 0.340 ;
        RECT  1.650 -0.280 7.800 0.280 ;
        RECT  0.610 -0.280 1.650 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.490 3.320 10.000 3.880 ;
        RECT  9.210 3.260 9.490 3.880 ;
        RECT  7.910 3.320 9.210 3.880 ;
        RECT  7.630 3.260 7.910 3.880 ;
        RECT  4.450 3.320 7.630 3.880 ;
        RECT  4.180 2.820 4.450 3.880 ;
        RECT  1.370 3.320 4.180 3.880 ;
        RECT  1.110 2.690 1.370 3.880 ;
        RECT  0.000 3.320 1.110 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.480 2.570 9.640 2.880 ;
        RECT  7.030 2.570 9.480 2.730 ;
        RECT  6.020 2.890 9.160 3.050 ;
        RECT  8.550 0.570 8.630 0.840 ;
        RECT  8.390 0.570 8.550 2.410 ;
        RECT  6.660 0.570 8.390 0.730 ;
        RECT  7.790 2.250 8.390 2.410 ;
        RECT  7.630 1.880 7.790 2.410 ;
        RECT  7.460 0.890 7.690 1.080 ;
        RECT  7.510 1.880 7.630 2.080 ;
        RECT  7.350 2.250 7.470 2.410 ;
        RECT  7.350 0.890 7.460 1.530 ;
        RECT  7.300 0.890 7.350 2.410 ;
        RECT  7.190 1.370 7.300 2.410 ;
        RECT  7.030 0.930 7.140 1.210 ;
        RECT  6.980 0.930 7.030 2.730 ;
        RECT  6.870 1.050 6.980 2.730 ;
        RECT  6.660 2.190 6.870 2.460 ;
        RECT  6.500 0.570 6.660 1.580 ;
        RECT  6.440 1.420 6.500 1.580 ;
        RECT  6.280 1.420 6.440 2.480 ;
        RECT  5.380 0.440 6.340 0.720 ;
        RECT  6.180 2.190 6.280 2.480 ;
        RECT  6.020 0.930 6.180 1.210 ;
        RECT  5.860 1.050 6.020 3.050 ;
        RECT  5.180 2.700 5.860 3.050 ;
        RECT  5.540 0.930 5.700 2.540 ;
        RECT  4.880 2.380 5.540 2.540 ;
        RECT  5.220 0.440 5.380 2.220 ;
        RECT  3.550 0.440 5.220 0.600 ;
        RECT  5.000 2.060 5.220 2.220 ;
        RECT  4.900 0.760 5.060 1.900 ;
        RECT  3.870 0.760 4.900 0.920 ;
        RECT  4.880 1.690 4.900 1.900 ;
        RECT  4.720 2.380 4.880 2.700 ;
        RECT  4.190 2.380 4.720 2.540 ;
        RECT  4.030 1.080 4.190 1.930 ;
        RECT  4.030 2.090 4.190 2.540 ;
        RECT  3.870 1.770 4.030 1.930 ;
        RECT  3.710 0.760 3.870 1.610 ;
        RECT  3.710 1.770 3.870 3.160 ;
        RECT  3.550 1.450 3.710 1.610 ;
        RECT  1.950 3.000 3.710 3.160 ;
        RECT  3.390 0.440 3.550 1.290 ;
        RECT  3.390 1.450 3.550 2.840 ;
        RECT  3.230 1.130 3.390 1.290 ;
        RECT  2.270 2.680 3.390 2.840 ;
        RECT  3.070 1.130 3.230 2.500 ;
        RECT  2.910 0.710 3.130 0.970 ;
        RECT  2.750 0.590 2.910 1.830 ;
        RECT  0.910 0.590 2.750 0.750 ;
        RECT  2.590 1.670 2.750 2.500 ;
        RECT  2.430 0.910 2.590 1.510 ;
        RECT  2.270 1.350 2.430 1.510 ;
        RECT  2.110 1.350 2.270 2.840 ;
        RECT  1.950 0.910 2.110 1.190 ;
        RECT  1.790 1.030 1.950 3.160 ;
        RECT  1.570 2.470 1.790 2.750 ;
        RECT  1.350 1.430 1.510 1.710 ;
        RECT  1.330 1.030 1.350 1.710 ;
        RECT  1.170 1.030 1.330 2.230 ;
        RECT  1.110 1.030 1.170 1.310 ;
        RECT  1.110 2.000 1.170 2.230 ;
        RECT  0.750 0.590 0.910 2.680 ;
        RECT  0.090 0.790 0.750 0.950 ;
        RECT  0.350 2.520 0.750 2.680 ;
        RECT  0.190 2.520 0.350 2.740 ;
    END
END ADDFHX1TR

MACRO ADDFXLTR
    CLASS CORE ;
    FOREIGN ADDFXLTR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.870 0.840 9.090 2.190 ;
        RECT  8.480 0.840 8.870 1.310 ;
        END
        ANTENNADIFFAREA 1.244 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.120 1.640 8.320 1.960 ;
        RECT  8.030 1.640 8.120 2.190 ;
        RECT  7.810 1.030 8.030 2.190 ;
        END
        ANTENNADIFFAREA 1.174 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 2.440 6.320 2.840 ;
        RECT  5.890 1.210 6.050 2.840 ;
        END
        ANTENNAGATEAREA 0.1632 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.580 0.510 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.1056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.410 3.120 1.960 ;
        RECT  2.510 1.410 2.870 1.690 ;
        END
        ANTENNAGATEAREA 0.1056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.550 -0.280 9.200 0.280 ;
        RECT  8.250 -0.280 8.550 0.670 ;
        RECT  6.270 -0.280 8.250 0.280 ;
        RECT  5.990 -0.280 6.270 0.330 ;
        RECT  2.970 -0.280 5.990 0.280 ;
        RECT  2.690 -0.280 2.970 0.610 ;
        RECT  0.890 -0.280 2.690 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 3.320 9.200 3.880 ;
        RECT  8.250 3.260 8.530 3.880 ;
        RECT  2.990 3.320 8.250 3.880 ;
        RECT  2.710 3.260 2.990 3.880 ;
        RECT  0.890 3.320 2.710 3.880 ;
        RECT  0.610 3.260 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.550 1.580 8.710 2.720 ;
        RECT  7.030 2.560 8.550 2.720 ;
        RECT  7.500 2.920 7.800 3.160 ;
        RECT  7.490 0.820 7.510 1.100 ;
        RECT  5.250 3.000 7.500 3.160 ;
        RECT  7.330 0.490 7.490 2.400 ;
        RECT  5.690 0.490 7.330 0.650 ;
        RECT  6.870 0.860 7.030 2.720 ;
        RECT  6.810 2.120 6.870 2.400 ;
        RECT  6.490 0.820 6.550 1.100 ;
        RECT  6.420 0.820 6.490 2.190 ;
        RECT  6.330 0.810 6.420 2.190 ;
        RECT  5.430 0.810 6.330 0.970 ;
        RECT  5.550 1.130 5.710 2.420 ;
        RECT  5.560 0.440 5.690 0.650 ;
        RECT  3.990 0.440 5.560 0.600 ;
        RECT  5.430 1.130 5.550 1.290 ;
        RECT  5.410 2.140 5.550 2.420 ;
        RECT  5.300 0.760 5.430 0.970 ;
        RECT  4.310 0.760 5.300 0.920 ;
        RECT  5.090 1.130 5.250 3.160 ;
        RECT  4.950 1.130 5.090 1.290 ;
        RECT  4.790 2.440 5.090 2.600 ;
        RECT  4.770 1.450 4.930 2.280 ;
        RECT  4.750 1.450 4.770 1.610 ;
        RECT  4.630 2.120 4.770 2.280 ;
        RECT  4.470 1.130 4.750 1.610 ;
        RECT  4.470 2.120 4.630 2.480 ;
        RECT  4.310 1.800 4.610 1.960 ;
        RECT  4.310 2.320 4.470 2.480 ;
        RECT  4.150 0.760 4.310 2.160 ;
        RECT  4.150 2.320 4.310 2.920 ;
        RECT  3.790 2.000 4.150 2.160 ;
        RECT  2.450 2.760 4.150 2.920 ;
        RECT  3.830 0.440 3.990 1.290 ;
        RECT  3.830 1.560 3.990 1.840 ;
        RECT  3.810 0.440 3.830 0.930 ;
        RECT  3.450 1.680 3.830 1.840 ;
        RECT  2.170 0.770 3.810 0.930 ;
        RECT  3.630 2.000 3.790 2.600 ;
        RECT  2.450 2.440 3.630 2.600 ;
        RECT  3.440 1.090 3.450 1.840 ;
        RECT  3.280 1.090 3.440 2.280 ;
        RECT  2.350 1.090 3.280 1.250 ;
        RECT  3.090 2.120 3.280 2.280 ;
        RECT  2.350 1.970 2.470 2.130 ;
        RECT  2.290 2.290 2.450 2.600 ;
        RECT  2.290 2.760 2.450 3.090 ;
        RECT  2.190 1.090 2.350 2.130 ;
        RECT  2.030 2.290 2.290 2.450 ;
        RECT  0.830 2.930 2.290 3.090 ;
        RECT  2.130 1.090 2.190 1.250 ;
        RECT  2.030 0.710 2.170 0.930 ;
        RECT  1.230 2.610 2.130 2.770 ;
        RECT  1.550 0.710 2.030 0.870 ;
        RECT  1.870 1.410 2.030 2.450 ;
        RECT  1.710 1.030 1.870 1.570 ;
        RECT  1.550 1.730 1.710 2.190 ;
        RECT  1.390 0.710 1.550 1.890 ;
        RECT  1.070 1.030 1.230 2.770 ;
        RECT  0.830 1.360 0.910 1.640 ;
        RECT  0.670 0.500 0.830 3.090 ;
        RECT  0.090 0.500 0.670 0.680 ;
        RECT  0.090 2.120 0.670 2.280 ;
    END
END ADDFXLTR

MACRO ADDFX4TR
    CLASS CORE ;
    FOREIGN ADDFX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.730 0.640 9.920 1.360 ;
        RECT  9.470 0.440 9.730 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.480 0.440 8.780 2.190 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.320 2.570 6.600 2.730 ;
        RECT  6.220 2.040 6.320 2.730 ;
        RECT  6.060 1.170 6.220 2.730 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.230 0.620 1.660 ;
        RECT  0.080 1.230 0.360 2.360 ;
        END
        ANTENNAGATEAREA 0.2616 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.450 3.120 1.960 ;
        RECT  2.540 1.450 2.880 1.610 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.310 -0.280 10.400 0.280 ;
        RECT  10.090 -0.280 10.310 1.310 ;
        RECT  9.250 -0.280 10.090 0.280 ;
        RECT  8.970 -0.280 9.250 1.310 ;
        RECT  8.160 -0.280 8.970 0.280 ;
        RECT  7.890 -0.280 8.160 1.180 ;
        RECT  6.360 -0.280 7.890 0.280 ;
        RECT  6.080 -0.280 6.360 0.340 ;
        RECT  3.160 -0.280 6.080 0.280 ;
        RECT  2.880 -0.280 3.160 0.580 ;
        RECT  0.000 -0.280 2.880 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.210 3.320 10.400 3.880 ;
        RECT  9.930 1.910 10.210 3.880 ;
        RECT  9.260 3.320 9.930 3.880 ;
        RECT  8.940 2.910 9.260 3.880 ;
        RECT  8.250 3.320 8.940 3.880 ;
        RECT  7.970 3.220 8.250 3.880 ;
        RECT  6.180 3.320 7.970 3.880 ;
        RECT  5.790 3.260 6.180 3.880 ;
        RECT  3.100 3.320 5.790 3.880 ;
        RECT  2.820 3.260 3.100 3.880 ;
        RECT  1.000 3.320 2.820 3.880 ;
        RECT  0.720 3.260 1.000 3.880 ;
        RECT  0.000 3.320 0.720 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.150 1.510 9.310 2.560 ;
        RECT  7.120 2.400 9.150 2.560 ;
        RECT  7.680 2.720 7.940 3.050 ;
        RECT  5.320 2.890 7.680 3.050 ;
        RECT  7.600 1.960 7.640 2.240 ;
        RECT  7.440 0.500 7.600 2.240 ;
        RECT  5.800 0.500 7.440 0.660 ;
        RECT  6.960 0.820 7.120 2.560 ;
        RECT  6.480 0.820 6.640 2.190 ;
        RECT  5.520 0.820 6.480 0.980 ;
        RECT  5.740 1.170 5.900 2.530 ;
        RECT  5.660 0.440 5.800 0.660 ;
        RECT  5.520 1.170 5.740 1.330 ;
        RECT  5.480 2.250 5.740 2.530 ;
        RECT  3.880 0.440 5.660 0.600 ;
        RECT  5.380 0.760 5.520 0.980 ;
        RECT  4.400 0.760 5.380 0.920 ;
        RECT  5.160 1.170 5.320 3.050 ;
        RECT  5.040 1.170 5.160 1.330 ;
        RECT  5.140 2.530 5.160 3.050 ;
        RECT  4.880 2.530 5.140 2.770 ;
        RECT  4.840 1.490 4.950 2.370 ;
        RECT  4.790 1.170 4.840 2.370 ;
        RECT  4.560 1.170 4.790 1.650 ;
        RECT  4.720 2.210 4.790 2.370 ;
        RECT  4.560 2.210 4.720 2.470 ;
        RECT  4.400 1.890 4.630 2.050 ;
        RECT  4.360 2.310 4.560 2.470 ;
        RECT  4.240 0.760 4.400 2.150 ;
        RECT  4.200 2.310 4.360 2.920 ;
        RECT  3.880 1.990 4.240 2.150 ;
        RECT  2.650 2.760 4.200 2.920 ;
        RECT  3.460 1.520 4.080 1.800 ;
        RECT  3.720 0.440 3.880 1.230 ;
        RECT  3.720 1.990 3.880 2.600 ;
        RECT  2.720 0.740 3.720 0.900 ;
        RECT  2.400 2.440 3.720 2.600 ;
        RECT  3.300 1.090 3.460 2.280 ;
        RECT  2.460 1.090 3.300 1.290 ;
        RECT  2.720 2.120 3.300 2.280 ;
        RECT  2.590 0.690 2.720 0.900 ;
        RECT  2.560 2.040 2.720 2.280 ;
        RECT  2.490 2.760 2.650 3.160 ;
        RECT  1.660 0.690 2.590 0.850 ;
        RECT  2.300 2.040 2.560 2.200 ;
        RECT  1.320 3.000 2.490 3.160 ;
        RECT  2.300 1.010 2.460 1.290 ;
        RECT  2.240 2.360 2.400 2.600 ;
        RECT  2.140 2.360 2.240 2.520 ;
        RECT  1.980 1.130 2.140 2.520 ;
        RECT  1.640 2.680 2.080 2.840 ;
        RECT  1.820 1.010 1.980 1.290 ;
        RECT  1.660 1.450 1.820 2.210 ;
        RECT  1.500 0.690 1.660 1.610 ;
        RECT  1.480 2.470 1.640 2.840 ;
        RECT  1.340 2.470 1.480 2.630 ;
        RECT  1.180 1.010 1.340 2.630 ;
        RECT  1.160 2.940 1.320 3.160 ;
        RECT  0.420 2.940 1.160 3.100 ;
        RECT  0.940 1.340 1.020 1.620 ;
        RECT  0.780 0.560 0.940 2.680 ;
        RECT  0.420 0.560 0.780 0.720 ;
        RECT  0.420 2.520 0.780 2.680 ;
        RECT  0.260 0.440 0.420 0.720 ;
        RECT  0.260 2.520 0.420 3.100 ;
    END
END ADDFX4TR

MACRO ADDFX2TR
    CLASS CORE ;
    FOREIGN ADDFX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.030 0.440 9.120 1.560 ;
        RECT  8.790 0.440 9.030 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.820 0.440 7.990 2.190 ;
        RECT  7.680 1.610 7.820 1.960 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.010 2.560 6.370 2.730 ;
        RECT  5.840 1.140 6.010 2.730 ;
        RECT  5.680 2.040 5.840 2.360 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.840 0.510 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.440 3.120 1.960 ;
        RECT  2.510 1.440 2.880 1.600 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 -0.280 9.200 0.280 ;
        RECT  8.250 -0.280 8.530 1.310 ;
        RECT  6.230 -0.280 8.250 0.280 ;
        RECT  5.950 -0.280 6.230 0.340 ;
        RECT  2.930 -0.280 5.950 0.280 ;
        RECT  2.650 -0.280 2.930 0.580 ;
        RECT  0.890 -0.280 2.650 0.280 ;
        RECT  0.610 -0.280 0.890 0.300 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 3.320 9.200 3.880 ;
        RECT  8.240 2.910 8.530 3.880 ;
        RECT  5.830 3.320 8.240 3.880 ;
        RECT  5.420 3.260 5.830 3.880 ;
        RECT  3.030 3.320 5.420 3.880 ;
        RECT  2.750 3.260 3.030 3.880 ;
        RECT  0.890 3.320 2.750 3.880 ;
        RECT  0.610 3.260 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.470 1.580 8.630 2.720 ;
        RECT  6.990 2.560 8.470 2.720 ;
        RECT  7.490 2.880 7.650 3.160 ;
        RECT  5.190 2.890 7.490 3.050 ;
        RECT  7.410 0.790 7.470 1.070 ;
        RECT  7.410 2.240 7.470 2.400 ;
        RECT  7.250 0.500 7.410 2.400 ;
        RECT  5.670 0.500 7.250 0.660 ;
        RECT  7.190 2.240 7.250 2.400 ;
        RECT  6.830 0.870 6.990 2.720 ;
        RECT  6.670 2.190 6.830 2.350 ;
        RECT  6.410 0.820 6.510 1.100 ;
        RECT  6.250 0.820 6.410 2.190 ;
        RECT  5.390 0.820 6.250 0.980 ;
        RECT  5.530 0.440 5.670 0.660 ;
        RECT  5.510 1.170 5.670 1.330 ;
        RECT  3.760 0.440 5.530 0.600 ;
        RECT  5.350 1.170 5.510 2.730 ;
        RECT  5.250 0.760 5.390 0.980 ;
        RECT  4.270 0.760 5.250 0.920 ;
        RECT  5.030 1.170 5.190 3.050 ;
        RECT  4.910 1.170 5.030 1.330 ;
        RECT  4.490 2.730 5.030 3.050 ;
        RECT  4.710 1.490 4.830 2.570 ;
        RECT  4.670 1.170 4.710 2.570 ;
        RECT  4.430 1.170 4.670 1.650 ;
        RECT  4.240 2.410 4.670 2.570 ;
        RECT  4.270 2.090 4.510 2.250 ;
        RECT  4.110 0.760 4.270 2.250 ;
        RECT  4.080 2.410 4.240 3.090 ;
        RECT  3.760 2.090 4.110 2.250 ;
        RECT  0.310 2.930 4.080 3.090 ;
        RECT  3.440 1.460 3.950 1.740 ;
        RECT  3.600 0.440 3.760 1.230 ;
        RECT  3.600 2.090 3.760 2.770 ;
        RECT  3.590 0.440 3.600 0.900 ;
        RECT  2.450 2.610 3.600 2.770 ;
        RECT  2.140 0.740 3.590 0.900 ;
        RECT  3.280 1.090 3.440 2.280 ;
        RECT  2.350 1.090 3.280 1.250 ;
        RECT  3.050 2.120 3.280 2.280 ;
        RECT  2.350 1.970 2.470 2.130 ;
        RECT  2.290 2.290 2.450 2.770 ;
        RECT  2.190 1.090 2.350 2.130 ;
        RECT  2.030 2.290 2.290 2.450 ;
        RECT  2.130 1.090 2.190 1.250 ;
        RECT  2.030 0.710 2.140 0.900 ;
        RECT  1.230 2.610 2.130 2.770 ;
        RECT  1.550 0.710 2.030 0.870 ;
        RECT  1.870 1.410 2.030 2.450 ;
        RECT  1.710 1.030 1.870 1.570 ;
        RECT  1.550 1.730 1.710 2.190 ;
        RECT  1.390 0.710 1.550 1.890 ;
        RECT  1.070 1.030 1.230 2.770 ;
        RECT  0.830 1.360 0.910 1.640 ;
        RECT  0.670 0.500 0.830 2.280 ;
        RECT  0.090 0.500 0.670 0.660 ;
        RECT  0.310 2.120 0.670 2.280 ;
        RECT  0.150 2.120 0.310 3.160 ;
    END
END ADDFX2TR

MACRO ADDFX1TR
    CLASS CORE ;
    FOREIGN ADDFX1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.800 1.030 9.120 2.550 ;
        RECT  8.740 1.030 8.800 1.310 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.830 1.030 8.040 2.190 ;
        RECT  7.780 1.030 7.830 1.960 ;
        RECT  7.680 1.610 7.780 1.960 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 2.370 6.390 2.760 ;
        RECT  6.020 2.370 6.080 2.550 ;
        RECT  5.860 1.140 6.020 2.550 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.240 0.520 1.670 ;
        RECT  0.080 1.240 0.330 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 1.440 3.120 1.960 ;
        RECT  2.590 1.440 2.800 1.770 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.540 -0.280 9.200 0.280 ;
        RECT  8.260 -0.280 8.540 1.130 ;
        RECT  6.240 -0.280 8.260 0.280 ;
        RECT  5.960 -0.280 6.240 0.340 ;
        RECT  2.940 -0.280 5.960 0.280 ;
        RECT  2.660 -0.280 2.940 0.580 ;
        RECT  0.900 -0.280 2.660 0.280 ;
        RECT  0.620 -0.280 0.900 0.300 ;
        RECT  0.000 -0.280 0.620 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.500 3.320 9.200 3.880 ;
        RECT  8.220 3.260 8.500 3.880 ;
        RECT  5.750 3.320 8.220 3.880 ;
        RECT  5.460 3.260 5.750 3.880 ;
        RECT  3.040 3.320 5.460 3.880 ;
        RECT  2.760 3.260 3.040 3.880 ;
        RECT  0.900 3.320 2.760 3.880 ;
        RECT  0.620 3.260 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.480 1.580 8.640 2.680 ;
        RECT  7.000 2.520 8.480 2.680 ;
        RECT  7.480 2.900 7.870 3.080 ;
        RECT  7.440 0.740 7.480 1.020 ;
        RECT  5.200 2.920 7.480 3.080 ;
        RECT  7.280 0.500 7.440 2.360 ;
        RECT  5.680 0.500 7.280 0.660 ;
        RECT  6.840 0.820 7.000 2.680 ;
        RECT  6.700 2.140 6.840 2.300 ;
        RECT  6.440 0.820 6.520 1.100 ;
        RECT  6.280 0.820 6.440 2.190 ;
        RECT  5.400 0.820 6.280 0.980 ;
        RECT  5.540 0.440 5.680 0.660 ;
        RECT  5.520 1.170 5.680 2.680 ;
        RECT  3.760 0.440 5.540 0.600 ;
        RECT  5.400 1.170 5.520 1.330 ;
        RECT  5.360 2.400 5.520 2.680 ;
        RECT  5.260 0.760 5.400 0.980 ;
        RECT  4.280 0.760 5.260 0.920 ;
        RECT  5.040 1.170 5.200 3.080 ;
        RECT  4.920 1.170 5.040 1.330 ;
        RECT  4.950 2.680 5.040 3.080 ;
        RECT  4.500 2.680 4.950 2.840 ;
        RECT  4.720 1.490 4.830 2.520 ;
        RECT  4.670 1.170 4.720 2.520 ;
        RECT  4.440 1.170 4.670 1.650 ;
        RECT  4.240 2.360 4.670 2.520 ;
        RECT  4.280 2.040 4.510 2.200 ;
        RECT  4.120 0.760 4.280 2.200 ;
        RECT  4.080 2.360 4.240 2.920 ;
        RECT  3.760 2.040 4.120 2.200 ;
        RECT  2.460 2.760 4.080 2.920 ;
        RECT  3.440 1.390 3.960 1.670 ;
        RECT  3.600 0.440 3.760 1.230 ;
        RECT  3.600 2.040 3.760 2.600 ;
        RECT  2.150 0.740 3.600 0.900 ;
        RECT  2.460 2.440 3.600 2.600 ;
        RECT  3.280 1.090 3.440 2.280 ;
        RECT  2.360 1.090 3.280 1.250 ;
        RECT  3.060 2.120 3.280 2.280 ;
        RECT  2.360 1.970 2.480 2.130 ;
        RECT  2.300 2.290 2.460 2.600 ;
        RECT  2.300 2.760 2.460 3.090 ;
        RECT  2.200 1.090 2.360 2.130 ;
        RECT  2.040 2.290 2.300 2.450 ;
        RECT  0.840 2.930 2.300 3.090 ;
        RECT  2.140 1.090 2.200 1.250 ;
        RECT  2.040 0.710 2.150 0.900 ;
        RECT  1.540 2.610 2.140 2.770 ;
        RECT  1.560 0.710 2.040 0.870 ;
        RECT  1.880 1.390 2.040 2.450 ;
        RECT  1.720 1.030 1.880 1.550 ;
        RECT  1.560 1.710 1.720 2.190 ;
        RECT  1.400 0.710 1.560 1.870 ;
        RECT  1.380 2.510 1.540 2.770 ;
        RECT  1.240 2.510 1.380 2.670 ;
        RECT  1.080 1.030 1.240 2.670 ;
        RECT  0.840 1.360 0.920 1.640 ;
        RECT  0.680 0.920 0.840 3.090 ;
        RECT  0.320 0.920 0.680 1.080 ;
        RECT  0.390 2.930 0.680 3.090 ;
        RECT  0.320 2.540 0.390 3.090 ;
        RECT  0.160 0.440 0.320 1.080 ;
        RECT  0.160 2.540 0.320 3.160 ;
    END
END ADDFX1TR

MACRO CMPR42X4TR
    CLASS CORE ;
    FOREIGN CMPR42X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  24.080 1.050 24.320 2.150 ;
        RECT  23.820 1.050 24.080 1.310 ;
        RECT  23.920 1.910 24.080 2.150 ;
        RECT  23.820 1.910 23.920 2.960 ;
        RECT  23.540 0.440 23.820 1.310 ;
        RECT  23.540 1.910 23.820 3.160 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.440 0.850 1.320 ;
        RECT  0.770 1.920 0.850 3.160 ;
        RECT  0.570 0.440 0.770 3.160 ;
        RECT  0.530 1.160 0.570 2.960 ;
        RECT  0.480 2.240 0.530 2.960 ;
        END
        ANTENNADIFFAREA 4.142 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  19.680 1.640 20.080 1.960 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.520 1.310 14.320 1.620 ;
        RECT  13.230 1.240 13.520 1.620 ;
        RECT  13.160 1.460 13.230 1.620 ;
        RECT  13.000 1.460 13.160 1.870 ;
        RECT  12.790 1.710 13.000 1.870 ;
        RECT  12.570 1.710 12.790 1.990 ;
        END
        ANTENNAGATEAREA 0.4848 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  18.120 1.030 18.380 1.760 ;
        RECT  17.800 1.030 18.120 2.210 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.470 2.940 13.680 3.160 ;
        RECT  12.310 2.880 12.470 3.160 ;
        RECT  11.030 2.880 12.310 3.040 ;
        RECT  10.870 2.880 11.030 3.160 ;
        RECT  10.030 3.000 10.870 3.160 ;
        RECT  9.870 2.840 10.030 3.160 ;
        RECT  8.360 2.840 9.870 3.000 ;
        RECT  8.040 2.840 8.360 3.160 ;
        RECT  3.610 2.840 8.040 3.000 ;
        RECT  3.450 2.840 3.610 3.160 ;
        RECT  3.330 2.940 3.450 3.160 ;
        END
        ANTENNAGATEAREA 0.6336 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.790 1.700 9.070 1.980 ;
        RECT  7.910 1.820 8.790 1.980 ;
        RECT  7.750 1.820 7.910 2.680 ;
        RECT  6.510 2.520 7.750 2.680 ;
        RECT  6.350 1.820 6.510 2.680 ;
        RECT  1.960 1.820 6.350 1.980 ;
        RECT  1.680 1.570 1.960 1.980 ;
        RECT  1.670 1.570 1.680 1.850 ;
        END
        ANTENNAGATEAREA 1.1712 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.990 1.500 7.270 1.920 ;
        RECT  4.760 1.500 6.990 1.660 ;
        RECT  4.480 1.240 4.760 1.660 ;
        RECT  2.750 1.500 4.480 1.660 ;
        RECT  2.590 1.250 2.750 1.660 ;
        RECT  2.470 1.250 2.590 1.530 ;
        RECT  1.490 1.250 2.470 1.410 ;
        RECT  1.330 1.250 1.490 1.640 ;
        END
        ANTENNAGATEAREA 1.0704 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  24.300 -0.280 24.400 0.280 ;
        RECT  24.020 -0.280 24.300 0.670 ;
        RECT  23.340 -0.280 24.020 0.280 ;
        RECT  23.120 -0.280 23.340 1.130 ;
        RECT  21.680 -0.280 23.120 0.280 ;
        RECT  21.400 -0.280 21.680 0.340 ;
        RECT  19.900 -0.280 21.400 0.280 ;
        RECT  19.680 -0.280 19.900 0.800 ;
        RECT  19.580 -0.280 19.680 0.400 ;
        RECT  18.960 -0.280 19.580 0.280 ;
        RECT  18.680 -0.280 18.960 0.400 ;
        RECT  17.920 -0.280 18.680 0.280 ;
        RECT  17.640 -0.280 17.920 0.400 ;
        RECT  14.240 -0.280 17.640 0.280 ;
        RECT  13.960 -0.280 14.240 0.380 ;
        RECT  9.450 -0.280 13.960 0.280 ;
        RECT  9.170 -0.280 9.450 0.550 ;
        RECT  7.450 -0.280 9.170 0.280 ;
        RECT  7.170 -0.280 7.450 0.880 ;
        RECT  6.670 -0.280 7.170 0.280 ;
        RECT  6.390 -0.280 6.670 1.340 ;
        RECT  5.670 -0.280 6.390 0.340 ;
        RECT  5.390 -0.280 5.670 0.760 ;
        RECT  4.630 -0.280 5.390 0.280 ;
        RECT  4.350 -0.280 4.630 0.400 ;
        RECT  2.990 -0.280 4.350 0.340 ;
        RECT  2.710 -0.280 2.990 0.400 ;
        RECT  1.350 -0.280 2.710 0.280 ;
        RECT  1.070 -0.280 1.350 0.680 ;
        RECT  0.370 -0.280 1.070 0.280 ;
        RECT  0.090 -0.280 0.370 1.320 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  24.300 3.320 24.400 3.880 ;
        RECT  24.080 2.360 24.300 3.880 ;
        RECT  23.260 3.320 24.080 3.880 ;
        RECT  22.980 2.930 23.260 3.880 ;
        RECT  21.620 3.320 22.980 3.880 ;
        RECT  21.340 3.200 21.620 3.880 ;
        RECT  19.760 3.320 21.340 3.880 ;
        RECT  19.480 3.200 19.760 3.880 ;
        RECT  18.600 3.320 19.480 3.880 ;
        RECT  18.320 3.200 18.600 3.880 ;
        RECT  17.560 3.320 18.320 3.880 ;
        RECT  17.280 3.200 17.560 3.880 ;
        RECT  14.370 3.320 17.280 3.880 ;
        RECT  14.090 2.160 14.370 3.880 ;
        RECT  12.150 3.320 14.090 3.880 ;
        RECT  11.870 3.200 12.150 3.880 ;
        RECT  9.710 3.320 11.870 3.880 ;
        RECT  9.430 3.200 9.710 3.880 ;
        RECT  7.830 3.320 9.430 3.880 ;
        RECT  7.550 3.200 7.830 3.880 ;
        RECT  7.030 3.260 7.550 3.880 ;
        RECT  6.750 3.200 7.030 3.880 ;
        RECT  5.670 3.320 6.750 3.880 ;
        RECT  5.390 3.200 5.670 3.880 ;
        RECT  4.630 3.320 5.390 3.880 ;
        RECT  4.350 3.200 4.630 3.880 ;
        RECT  2.990 3.320 4.350 3.880 ;
        RECT  2.710 3.200 2.990 3.880 ;
        RECT  1.350 3.260 2.710 3.880 ;
        RECT  1.070 2.670 1.350 3.880 ;
        RECT  0.320 3.320 1.070 3.880 ;
        RECT  0.090 1.800 0.320 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  23.380 1.470 23.860 1.750 ;
        RECT  23.220 1.290 23.380 2.680 ;
        RECT  22.960 1.290 23.220 1.450 ;
        RECT  22.460 2.520 23.220 2.680 ;
        RECT  22.640 1.640 23.060 1.920 ;
        RECT  22.800 0.500 22.960 1.450 ;
        RECT  20.580 0.500 22.800 0.720 ;
        RECT  22.480 0.880 22.640 2.360 ;
        RECT  20.100 0.880 22.480 1.160 ;
        RECT  21.860 2.200 22.480 2.360 ;
        RECT  22.340 2.520 22.460 2.800 ;
        RECT  22.180 2.520 22.340 3.040 ;
        RECT  22.040 1.320 22.320 1.600 ;
        RECT  22.020 1.760 22.300 2.040 ;
        RECT  20.480 2.820 22.180 3.040 ;
        RECT  20.560 1.320 22.040 1.480 ;
        RECT  21.000 1.760 22.020 1.920 ;
        RECT  21.580 2.080 21.860 2.360 ;
        RECT  21.240 2.200 21.580 2.360 ;
        RECT  21.080 2.200 21.240 2.660 ;
        RECT  20.280 2.440 21.080 2.660 ;
        RECT  20.880 1.640 21.000 1.920 ;
        RECT  20.720 1.640 20.880 2.280 ;
        RECT  19.240 2.120 20.720 2.280 ;
        RECT  20.280 1.320 20.560 1.960 ;
        RECT  19.520 1.320 20.280 1.480 ;
        RECT  20.000 2.440 20.280 3.160 ;
        RECT  17.110 2.880 20.000 3.040 ;
        RECT  19.360 0.560 19.520 1.730 ;
        RECT  17.480 0.560 19.360 0.720 ;
        RECT  19.240 1.450 19.360 1.730 ;
        RECT  19.080 1.970 19.240 2.720 ;
        RECT  19.080 1.010 19.200 1.290 ;
        RECT  18.980 1.010 19.080 2.720 ;
        RECT  18.920 1.130 18.980 2.720 ;
        RECT  17.430 2.560 18.920 2.720 ;
        RECT  17.260 0.440 17.480 0.720 ;
        RECT  17.270 1.920 17.430 2.720 ;
        RECT  17.100 0.880 17.300 1.100 ;
        RECT  17.110 1.920 17.270 2.200 ;
        RECT  15.020 0.440 17.260 0.600 ;
        RECT  16.950 2.450 17.110 3.040 ;
        RECT  16.940 0.760 17.100 1.100 ;
        RECT  16.790 1.260 16.950 3.160 ;
        RECT  16.340 0.760 16.940 0.920 ;
        RECT  16.780 1.260 16.790 1.420 ;
        RECT  15.870 2.940 16.790 3.160 ;
        RECT  16.620 1.080 16.780 1.420 ;
        RECT  16.510 1.580 16.630 1.800 ;
        RECT  16.510 2.190 16.630 2.470 ;
        RECT  16.500 1.080 16.620 1.360 ;
        RECT  16.350 1.580 16.510 2.780 ;
        RECT  16.340 1.580 16.350 1.740 ;
        RECT  15.330 2.620 16.350 2.780 ;
        RECT  16.180 0.760 16.340 1.740 ;
        RECT  15.400 0.760 16.180 0.980 ;
        RECT  15.690 1.160 15.920 1.440 ;
        RECT  15.690 2.180 15.810 2.460 ;
        RECT  15.640 1.160 15.690 2.460 ;
        RECT  15.530 1.280 15.640 2.460 ;
        RECT  14.850 2.180 15.530 2.340 ;
        RECT  15.180 0.760 15.400 1.040 ;
        RECT  15.050 2.500 15.330 3.160 ;
        RECT  15.020 1.740 15.140 2.020 ;
        RECT  14.860 0.440 15.020 2.020 ;
        RECT  14.560 0.440 14.860 0.600 ;
        RECT  14.700 2.180 14.850 3.160 ;
        RECT  14.540 0.980 14.700 3.160 ;
        RECT  14.400 0.440 14.560 0.700 ;
        RECT  14.480 0.980 14.540 2.000 ;
        RECT  13.600 1.840 14.480 2.000 ;
        RECT  13.070 0.540 14.400 0.700 ;
        RECT  13.190 2.160 13.890 2.440 ;
        RECT  13.070 0.860 13.710 1.080 ;
        RECT  13.320 1.780 13.600 2.000 ;
        RECT  12.410 2.160 13.190 2.320 ;
        RECT  12.910 0.440 13.070 0.700 ;
        RECT  12.910 0.860 13.070 1.300 ;
        RECT  12.710 2.480 12.990 2.760 ;
        RECT  11.720 0.440 12.910 0.600 ;
        RECT  12.410 1.140 12.910 1.300 ;
        RECT  12.040 0.760 12.750 0.920 ;
        RECT  11.850 2.480 12.710 2.640 ;
        RECT  12.250 1.140 12.410 2.320 ;
        RECT  12.110 1.710 12.250 1.990 ;
        RECT  11.880 0.760 12.040 1.360 ;
        RECT  11.850 1.200 11.880 1.360 ;
        RECT  11.690 1.200 11.850 2.640 ;
        RECT  11.560 0.440 11.720 1.040 ;
        RECT  11.030 1.200 11.690 1.420 ;
        RECT  11.630 2.040 11.690 2.320 ;
        RECT  10.710 0.880 11.560 1.040 ;
        RECT  11.450 1.620 11.470 1.900 ;
        RECT  11.290 1.620 11.450 2.680 ;
        RECT  11.120 0.440 11.400 0.720 ;
        RECT  11.190 1.620 11.290 1.900 ;
        RECT  10.710 2.520 11.290 2.680 ;
        RECT  10.910 2.080 11.130 2.360 ;
        RECT  10.270 0.480 11.120 0.720 ;
        RECT  10.870 1.200 11.030 1.920 ;
        RECT  10.590 2.080 10.910 2.240 ;
        RECT  10.750 1.640 10.870 1.920 ;
        RECT  10.590 0.880 10.710 1.160 ;
        RECT  10.430 2.520 10.710 2.840 ;
        RECT  10.430 0.880 10.590 2.240 ;
        RECT  9.830 2.520 10.430 2.680 ;
        RECT  10.110 0.480 10.270 2.330 ;
        RECT  9.950 0.480 10.110 0.640 ;
        RECT  9.990 2.040 10.110 2.330 ;
        RECT  9.830 1.300 9.950 1.580 ;
        RECT  9.670 0.800 9.830 2.680 ;
        RECT  8.450 0.800 9.670 0.960 ;
        RECT  8.870 2.520 9.670 2.680 ;
        RECT  9.390 1.320 9.510 1.600 ;
        RECT  9.230 1.120 9.390 2.300 ;
        RECT  7.970 1.120 9.230 1.280 ;
        RECT  8.350 2.140 9.230 2.300 ;
        RECT  8.590 2.460 8.870 2.680 ;
        RECT  7.590 1.440 8.630 1.660 ;
        RECT  8.170 0.680 8.450 0.960 ;
        RECT  8.070 2.140 8.350 2.420 ;
        RECT  7.810 0.740 7.970 1.280 ;
        RECT  7.690 0.740 7.810 1.020 ;
        RECT  7.430 1.180 7.590 2.360 ;
        RECT  7.150 1.180 7.430 1.340 ;
        RECT  6.790 2.080 7.430 2.360 ;
        RECT  6.870 1.060 7.150 1.340 ;
        RECT  5.910 0.650 6.190 1.340 ;
        RECT  5.910 2.140 6.190 2.460 ;
        RECT  5.150 0.920 5.910 1.080 ;
        RECT  5.150 2.140 5.910 2.300 ;
        RECT  4.870 0.660 5.150 1.080 ;
        RECT  4.870 2.140 5.150 2.460 ;
        RECT  3.530 0.660 4.870 0.940 ;
        RECT  3.530 2.140 4.870 2.360 ;
        RECT  3.330 1.100 4.290 1.320 ;
        RECT  3.330 2.520 4.290 2.680 ;
        RECT  3.050 0.930 3.330 1.320 ;
        RECT  3.050 2.370 3.330 2.680 ;
        RECT  2.150 0.930 3.050 1.090 ;
        RECT  2.150 2.520 3.050 2.680 ;
        RECT  1.870 0.440 2.150 1.090 ;
        RECT  1.870 2.140 2.150 2.860 ;
        RECT  1.170 0.930 1.870 1.090 ;
        RECT  1.170 2.140 1.870 2.300 ;
        RECT  1.010 0.930 1.170 2.300 ;
        RECT  0.930 1.480 1.010 1.760 ;
    END
END CMPR42X4TR

MACRO CMPR42X2TR
    CLASS CORE ;
    FOREIGN CMPR42X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.880 0.450 17.120 2.760 ;
        RECT  16.780 0.450 16.880 1.250 ;
        RECT  16.780 1.910 16.880 2.760 ;
        RECT  16.620 1.910 16.780 3.160 ;
        END
        ANTENNADIFFAREA 3.488 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 1.640 0.320 3.160 ;
        RECT  0.080 0.440 0.310 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.370 1.610 14.720 1.960 ;
        END
        ANTENNAGATEAREA 0.252 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.720 1.420 10.950 1.580 ;
        RECT  10.540 1.240 10.720 1.580 ;
        RECT  10.480 1.240 10.540 1.560 ;
        RECT  10.020 1.400 10.480 1.560 ;
        RECT  9.860 1.280 10.020 1.560 ;
        RECT  9.260 1.400 9.860 1.560 ;
        RECT  9.100 1.400 9.260 1.900 ;
        END
        ANTENNAGATEAREA 0.5016 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.440 2.040 13.520 2.360 ;
        RECT  13.280 0.820 13.440 2.360 ;
        RECT  12.790 0.820 13.280 0.980 ;
        RECT  12.910 2.100 13.280 2.360 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 2.880 10.630 3.160 ;
        RECT  8.960 3.000 10.470 3.160 ;
        RECT  8.820 2.940 8.960 3.160 ;
        RECT  7.450 2.940 8.820 3.100 ;
        RECT  7.290 2.940 7.450 3.160 ;
        RECT  6.720 3.000 7.290 3.160 ;
        RECT  6.480 2.840 6.720 3.160 ;
        RECT  2.010 2.940 6.480 3.100 ;
        RECT  1.850 2.940 2.010 3.160 ;
        RECT  1.730 3.000 1.850 3.160 ;
        END
        ANTENNAGATEAREA 0.4608 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 1.710 5.610 2.020 ;
        RECT  4.610 1.860 5.450 2.020 ;
        RECT  4.450 1.860 4.610 2.680 ;
        RECT  3.470 2.520 4.450 2.680 ;
        RECT  3.470 1.760 3.630 1.920 ;
        RECT  3.310 1.760 3.470 2.680 ;
        RECT  1.530 1.760 3.310 1.920 ;
        RECT  1.520 1.600 1.530 1.920 ;
        RECT  1.250 1.600 1.520 1.960 ;
        END
        ANTENNAGATEAREA 0.7512 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.810 1.440 3.970 1.980 ;
        RECT  2.490 1.440 3.810 1.600 ;
        RECT  2.080 1.240 2.490 1.600 ;
        RECT  1.070 1.280 2.080 1.440 ;
        RECT  0.910 1.280 1.070 1.640 ;
        END
        ANTENNAGATEAREA 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.540 -0.280 17.200 0.280 ;
        RECT  16.260 -0.280 16.540 0.340 ;
        RECT  14.590 -0.280 16.260 0.280 ;
        RECT  14.310 -0.280 14.590 0.340 ;
        RECT  13.790 -0.280 14.310 0.280 ;
        RECT  13.510 -0.280 13.790 0.340 ;
        RECT  10.810 -0.280 13.510 0.280 ;
        RECT  10.530 -0.280 10.810 0.340 ;
        RECT  6.110 -0.280 10.530 0.280 ;
        RECT  5.830 -0.280 6.110 0.740 ;
        RECT  4.180 -0.280 5.830 0.280 ;
        RECT  3.910 -0.280 4.180 0.960 ;
        RECT  2.730 -0.280 3.910 0.280 ;
        RECT  2.450 -0.280 2.730 0.760 ;
        RECT  0.890 -0.280 2.450 0.280 ;
        RECT  0.610 -0.280 0.890 0.800 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.320 3.320 17.200 3.880 ;
        RECT  16.040 3.260 16.320 3.880 ;
        RECT  14.150 3.320 16.040 3.880 ;
        RECT  13.430 3.260 14.150 3.880 ;
        RECT  10.950 3.320 13.430 3.880 ;
        RECT  10.790 2.160 10.950 3.880 ;
        RECT  10.200 2.160 10.790 2.320 ;
        RECT  8.680 3.320 10.790 3.880 ;
        RECT  8.400 3.260 8.680 3.880 ;
        RECT  6.310 3.320 8.400 3.880 ;
        RECT  6.030 3.260 6.310 3.880 ;
        RECT  4.470 3.320 6.030 3.880 ;
        RECT  3.330 3.260 4.470 3.880 ;
        RECT  2.510 3.320 3.330 3.880 ;
        RECT  2.230 3.260 2.510 3.880 ;
        RECT  0.890 3.320 2.230 3.880 ;
        RECT  0.610 2.650 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  16.460 1.440 16.640 1.600 ;
        RECT  16.300 0.610 16.460 2.940 ;
        RECT  15.640 0.610 16.300 0.770 ;
        RECT  15.090 2.760 16.300 2.940 ;
        RECT  16.020 0.930 16.140 1.770 ;
        RECT  15.980 0.930 16.020 2.600 ;
        RECT  15.230 0.930 15.980 1.090 ;
        RECT  15.860 1.610 15.980 2.600 ;
        RECT  14.890 2.440 15.860 2.600 ;
        RECT  15.040 1.270 15.820 1.430 ;
        RECT  15.480 0.490 15.640 0.770 ;
        RECT  15.280 1.610 15.440 2.280 ;
        RECT  14.130 2.120 15.280 2.280 ;
        RECT  14.950 0.490 15.230 1.090 ;
        RECT  14.880 1.270 15.040 1.890 ;
        RECT  14.610 2.440 14.890 3.000 ;
        RECT  14.450 1.270 14.880 1.430 ;
        RECT  12.350 2.840 14.610 3.000 ;
        RECT  14.290 0.710 14.450 1.430 ;
        RECT  13.770 0.710 14.290 0.870 ;
        RECT  13.970 1.030 14.130 2.280 ;
        RECT  13.930 1.030 13.970 1.310 ;
        RECT  13.950 2.050 13.970 2.280 ;
        RECT  13.790 2.050 13.950 2.680 ;
        RECT  13.770 1.430 13.810 1.710 ;
        RECT  12.390 2.520 13.790 2.680 ;
        RECT  13.610 0.500 13.770 1.710 ;
        RECT  12.750 0.500 13.610 0.660 ;
        RECT  12.960 1.140 13.120 1.940 ;
        RECT  12.390 1.140 12.960 1.300 ;
        RECT  12.230 1.780 12.960 1.940 ;
        RECT  11.910 1.460 12.800 1.620 ;
        RECT  12.500 0.440 12.750 0.660 ;
        RECT  11.590 0.500 12.500 0.660 ;
        RECT  12.230 0.870 12.390 1.300 ;
        RECT  12.230 2.840 12.350 3.150 ;
        RECT  12.070 1.780 12.230 3.150 ;
        RECT  11.750 0.870 11.910 3.160 ;
        RECT  11.580 2.300 11.750 3.160 ;
        RECT  11.430 0.500 11.590 2.140 ;
        RECT  9.700 0.500 11.430 0.660 ;
        RECT  11.270 2.300 11.370 3.160 ;
        RECT  11.110 1.030 11.270 3.160 ;
        RECT  9.820 1.840 11.110 2.000 ;
        RECT  9.700 0.960 10.280 1.120 ;
        RECT  9.780 2.160 9.940 2.840 ;
        RECT  9.660 1.720 9.820 2.000 ;
        RECT  8.940 2.160 9.780 2.320 ;
        RECT  9.540 0.440 9.700 0.660 ;
        RECT  9.540 0.960 9.700 1.240 ;
        RECT  9.220 2.510 9.570 2.760 ;
        RECT  8.100 0.440 9.540 0.600 ;
        RECT  8.940 1.080 9.540 1.240 ;
        RECT  8.420 0.760 9.380 0.920 ;
        RECT  8.250 2.510 9.220 2.670 ;
        RECT  8.780 1.080 8.940 2.320 ;
        RECT  8.640 1.680 8.780 1.840 ;
        RECT  8.260 0.760 8.420 1.360 ;
        RECT  8.250 1.200 8.260 1.360 ;
        RECT  8.090 1.200 8.250 2.670 ;
        RECT  7.940 0.440 8.100 1.040 ;
        RECT  7.410 1.200 8.090 1.360 ;
        RECT  7.090 0.880 7.940 1.040 ;
        RECT  7.770 1.680 7.930 2.720 ;
        RECT  7.620 0.440 7.780 0.720 ;
        RECT  7.730 1.680 7.770 1.960 ;
        RECT  7.130 2.560 7.770 2.720 ;
        RECT  6.770 0.560 7.620 0.720 ;
        RECT  7.450 2.120 7.610 2.400 ;
        RECT  7.090 2.120 7.450 2.280 ;
        RECT  7.250 1.200 7.410 1.960 ;
        RECT  7.090 2.560 7.130 2.840 ;
        RECT  6.930 0.880 7.090 2.280 ;
        RECT  6.970 2.520 7.090 2.840 ;
        RECT  6.330 2.520 6.970 2.680 ;
        RECT  6.610 0.560 6.770 2.360 ;
        RECT  6.390 0.560 6.610 0.720 ;
        RECT  6.540 1.990 6.610 2.360 ;
        RECT  6.330 1.320 6.440 1.630 ;
        RECT  6.170 0.900 6.330 2.680 ;
        RECT  5.130 0.900 6.170 1.060 ;
        RECT  5.190 2.520 6.170 2.680 ;
        RECT  5.930 1.330 6.010 1.730 ;
        RECT  5.770 1.330 5.930 2.340 ;
        RECT  5.590 1.330 5.770 1.550 ;
        RECT  4.930 2.180 5.770 2.340 ;
        RECT  5.430 1.220 5.590 1.550 ;
        RECT  4.670 1.220 5.430 1.380 ;
        RECT  4.290 1.540 5.270 1.700 ;
        RECT  4.890 0.450 5.130 1.060 ;
        RECT  4.770 2.180 4.930 2.460 ;
        RECT  4.510 0.800 4.670 1.380 ;
        RECT  4.390 0.800 4.510 0.960 ;
        RECT  4.130 1.120 4.290 2.360 ;
        RECT  3.610 1.120 4.130 1.280 ;
        RECT  3.630 2.200 4.130 2.360 ;
        RECT  3.450 1.000 3.610 1.280 ;
        RECT  3.030 0.530 3.190 1.080 ;
        RECT  2.210 0.920 3.030 1.080 ;
        RECT  2.730 2.200 3.010 2.780 ;
        RECT  2.210 2.200 2.730 2.360 ;
        RECT  1.930 0.590 2.210 1.080 ;
        RECT  1.990 2.080 2.210 2.700 ;
        RECT  1.450 0.590 1.730 1.120 ;
        RECT  1.690 2.120 1.710 2.710 ;
        RECT  1.450 2.120 1.690 2.840 ;
        RECT  0.750 0.960 1.450 1.120 ;
        RECT  0.750 2.120 1.450 2.280 ;
        RECT  0.590 0.960 0.750 2.280 ;
        RECT  0.480 1.470 0.590 1.750 ;
    END
END CMPR42X2TR

MACRO CMPR42X1TR
    CLASS CORE ;
    FOREIGN CMPR42X1TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.760 0.750 15.920 2.760 ;
        RECT  15.560 0.750 15.760 0.910 ;
        RECT  15.680 1.640 15.760 2.760 ;
        RECT  15.580 1.910 15.680 2.550 ;
        RECT  15.400 0.630 15.560 0.910 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.640 0.320 2.760 ;
        RECT  0.240 1.030 0.310 1.310 ;
        RECT  0.080 1.030 0.240 2.760 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.520 2.250 13.560 2.410 ;
        RECT  13.280 2.250 13.520 2.760 ;
        END
        ANTENNAGATEAREA 0.144 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.680 1.220 9.980 1.640 ;
        END
        ANTENNAGATEAREA 0.3336 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.240 0.840 12.320 1.200 ;
        RECT  12.080 0.840 12.240 2.320 ;
        RECT  11.980 0.840 12.080 1.200 ;
        RECT  12.040 2.040 12.080 2.320 ;
        END
        ANTENNADIFFAREA 1.76 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.340 2.760 9.500 3.040 ;
        RECT  7.520 2.760 9.340 2.920 ;
        RECT  7.360 2.760 7.520 3.130 ;
        RECT  6.240 2.970 7.360 3.130 ;
        RECT  6.080 2.940 6.240 3.130 ;
        RECT  1.790 2.940 6.080 3.100 ;
        RECT  1.630 2.590 1.790 3.100 ;
        RECT  1.520 2.840 1.630 3.100 ;
        RECT  1.280 2.840 1.520 3.160 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.980 1.740 5.140 2.020 ;
        RECT  4.220 1.860 4.980 2.020 ;
        RECT  4.060 1.860 4.220 2.780 ;
        RECT  3.010 2.620 4.060 2.780 ;
        RECT  2.850 1.830 3.010 2.780 ;
        RECT  2.670 1.830 2.850 2.250 ;
        RECT  1.920 1.830 2.670 1.990 ;
        RECT  1.170 1.640 1.920 1.990 ;
        END
        ANTENNAGATEAREA 0.4248 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.510 3.580 1.930 ;
        RECT  2.410 1.510 3.420 1.670 ;
        RECT  2.080 1.240 2.410 1.670 ;
        RECT  1.070 1.320 2.080 1.480 ;
        RECT  0.910 1.200 1.070 1.480 ;
        END
        ANTENNAGATEAREA 0.3672 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.100 -0.280 16.000 0.280 ;
        RECT  14.820 -0.280 15.100 0.340 ;
        RECT  13.220 -0.280 14.820 0.280 ;
        RECT  12.500 -0.280 13.220 0.340 ;
        RECT  9.980 -0.280 12.500 0.280 ;
        RECT  9.820 -0.280 9.980 0.720 ;
        RECT  8.080 -0.280 9.820 0.280 ;
        RECT  7.800 -0.280 8.080 0.340 ;
        RECT  3.750 -0.280 7.800 0.280 ;
        RECT  3.590 -0.280 3.750 1.030 ;
        RECT  2.730 -0.280 3.590 0.280 ;
        RECT  2.450 -0.280 2.730 0.340 ;
        RECT  0.890 -0.280 2.450 0.280 ;
        RECT  0.610 -0.280 0.890 0.340 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.300 3.320 16.000 3.880 ;
        RECT  15.020 3.260 15.300 3.880 ;
        RECT  13.190 3.320 15.020 3.880 ;
        RECT  12.500 3.260 13.190 3.880 ;
        RECT  9.820 3.320 12.500 3.880 ;
        RECT  9.660 2.410 9.820 3.880 ;
        RECT  8.080 3.320 9.660 3.880 ;
        RECT  7.800 3.260 8.080 3.880 ;
        RECT  5.920 3.320 7.800 3.880 ;
        RECT  5.640 3.260 5.920 3.880 ;
        RECT  4.080 3.320 5.640 3.880 ;
        RECT  3.800 3.260 4.080 3.880 ;
        RECT  3.210 3.320 3.800 3.880 ;
        RECT  2.930 3.260 3.210 3.880 ;
        RECT  2.130 3.320 2.930 3.880 ;
        RECT  1.850 3.260 2.130 3.880 ;
        RECT  0.770 3.320 1.850 3.880 ;
        RECT  0.490 3.260 0.770 3.880 ;
        RECT  0.000 3.320 0.490 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.240 1.070 15.420 1.230 ;
        RECT  15.080 0.610 15.240 3.040 ;
        RECT  13.940 0.610 15.080 0.770 ;
        RECT  14.400 2.880 15.080 3.040 ;
        RECT  14.760 0.930 14.920 2.720 ;
        RECT  13.680 0.930 14.760 1.090 ;
        RECT  13.880 2.560 14.760 2.720 ;
        RECT  14.440 1.250 14.600 2.400 ;
        RECT  13.160 1.250 14.440 1.410 ;
        RECT  13.120 1.930 14.440 2.090 ;
        RECT  14.240 2.880 14.400 3.160 ;
        RECT  12.840 1.610 14.280 1.770 ;
        RECT  13.720 2.560 13.880 3.080 ;
        RECT  11.270 2.920 13.720 3.080 ;
        RECT  13.520 0.630 13.680 1.090 ;
        RECT  13.000 1.160 13.160 1.440 ;
        RECT  12.960 1.930 13.120 2.640 ;
        RECT  11.590 2.480 12.960 2.640 ;
        RECT  12.680 0.500 12.840 1.770 ;
        RECT  12.140 0.500 12.680 0.660 ;
        RECT  11.980 0.440 12.140 0.660 ;
        RECT  10.940 0.440 11.980 0.600 ;
        RECT  11.660 0.850 11.820 2.320 ;
        RECT  11.520 0.850 11.660 1.010 ;
        RECT  11.270 2.160 11.660 2.320 ;
        RECT  11.430 2.480 11.590 2.760 ;
        RECT  11.260 1.460 11.500 1.740 ;
        RECT  11.110 2.160 11.270 3.080 ;
        RECT  11.100 0.790 11.260 2.000 ;
        RECT  11.100 2.160 11.110 2.440 ;
        RECT  10.940 1.840 11.100 2.000 ;
        RECT  10.780 0.440 10.940 1.680 ;
        RECT  10.780 1.840 10.940 2.400 ;
        RECT  10.300 0.440 10.780 0.600 ;
        RECT  10.620 1.520 10.780 1.680 ;
        RECT  10.560 2.240 10.780 2.400 ;
        RECT  10.460 1.030 10.620 1.360 ;
        RECT  10.460 1.520 10.620 2.080 ;
        RECT  10.300 1.200 10.460 1.360 ;
        RECT  10.140 0.440 10.300 1.040 ;
        RECT  10.140 1.200 10.300 2.520 ;
        RECT  9.660 0.880 10.140 1.040 ;
        RECT  9.120 1.800 10.140 1.960 ;
        RECT  9.500 0.590 9.660 1.040 ;
        RECT  6.920 0.590 9.500 0.750 ;
        RECT  9.180 0.910 9.340 1.450 ;
        RECT  9.180 2.120 9.340 2.400 ;
        RECT  8.680 1.290 9.180 1.450 ;
        RECT  8.680 2.120 9.180 2.280 ;
        RECT  8.840 1.640 9.120 1.960 ;
        RECT  7.520 0.970 8.920 1.130 ;
        RECT  7.680 2.440 8.920 2.600 ;
        RECT  8.520 1.290 8.680 2.280 ;
        RECT  8.040 1.880 8.520 2.040 ;
        RECT  7.520 2.030 7.680 2.600 ;
        RECT  7.360 0.970 7.520 2.600 ;
        RECT  7.240 0.970 7.360 1.310 ;
        RECT  6.860 1.760 7.360 1.920 ;
        RECT  7.040 2.080 7.200 2.810 ;
        RECT  6.700 2.080 7.040 2.240 ;
        RECT  6.760 0.590 6.920 1.310 ;
        RECT  6.700 1.150 6.760 1.310 ;
        RECT  6.560 2.530 6.720 2.810 ;
        RECT  6.540 1.150 6.700 2.240 ;
        RECT  6.060 2.530 6.560 2.690 ;
        RECT  6.380 0.830 6.500 0.990 ;
        RECT  6.220 0.560 6.380 2.350 ;
        RECT  5.840 0.560 6.220 0.720 ;
        RECT  5.900 0.880 6.060 2.690 ;
        RECT  4.710 0.880 5.900 1.040 ;
        RECT  4.800 2.530 5.900 2.690 ;
        RECT  5.680 0.440 5.840 0.720 ;
        RECT  5.460 1.280 5.540 1.560 ;
        RECT  5.300 1.200 5.460 2.360 ;
        RECT  4.230 1.200 5.300 1.360 ;
        RECT  4.540 2.200 5.300 2.360 ;
        RECT  3.900 1.520 4.800 1.680 ;
        RECT  4.550 0.750 4.710 1.040 ;
        RECT  4.380 2.200 4.540 2.480 ;
        RECT  4.070 0.750 4.230 1.360 ;
        RECT  3.740 1.190 3.900 2.460 ;
        RECT  3.430 1.190 3.740 1.350 ;
        RECT  3.370 2.300 3.740 2.460 ;
        RECT  3.270 0.560 3.430 1.350 ;
        RECT  3.190 0.560 3.270 0.720 ;
        RECT  3.030 0.440 3.190 0.720 ;
        RECT  2.950 0.910 3.110 1.190 ;
        RECT  2.150 0.910 2.950 1.070 ;
        RECT  2.110 2.410 2.690 2.570 ;
        RECT  1.990 0.790 2.150 1.070 ;
        RECT  2.070 2.270 2.110 2.570 ;
        RECT  1.950 2.150 2.070 2.570 ;
        RECT  1.910 2.150 1.950 2.430 ;
        RECT  1.510 0.790 1.670 1.070 ;
        RECT  1.430 2.150 1.590 2.430 ;
        RECT  0.750 0.880 1.510 1.040 ;
        RECT  0.750 2.150 1.430 2.310 ;
        RECT  0.590 0.880 0.750 2.310 ;
        RECT  0.480 1.520 0.590 1.800 ;
    END
END CMPR42X1TR

MACRO CMPR32X4TR
    CLASS CORE ;
    FOREIGN CMPR32X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.120 0.440 9.360 3.160 ;
        RECT  9.060 0.440 9.120 1.310 ;
        RECT  9.060 1.840 9.120 3.160 ;
        RECT  8.880 1.840 9.060 2.560 ;
        END
        ANTENNADIFFAREA 4.328 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.440 8.320 2.780 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 2.040 5.920 2.450 ;
        END
        ANTENNAGATEAREA 0.2064 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.350 0.510 1.720 ;
        RECT  0.380 1.350 0.400 1.960 ;
        RECT  0.080 0.840 0.380 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.440 3.120 1.960 ;
        RECT  2.570 1.440 2.880 1.600 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 -0.280 10.000 0.280 ;
        RECT  9.550 -0.280 9.830 1.310 ;
        RECT  8.790 -0.280 9.550 0.280 ;
        RECT  8.510 -0.280 8.790 1.280 ;
        RECT  7.830 -0.280 8.510 0.280 ;
        RECT  7.550 -0.280 7.830 1.310 ;
        RECT  6.070 -0.280 7.550 0.280 ;
        RECT  5.790 -0.280 6.070 0.340 ;
        RECT  2.930 -0.280 5.790 0.280 ;
        RECT  2.650 -0.280 2.930 0.600 ;
        RECT  0.890 -0.280 2.650 0.280 ;
        RECT  0.610 -0.280 0.890 0.300 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.830 3.320 10.000 3.880 ;
        RECT  9.550 1.910 9.830 3.880 ;
        RECT  8.830 3.320 9.550 3.880 ;
        RECT  8.550 3.260 8.830 3.880 ;
        RECT  7.790 3.320 8.550 3.880 ;
        RECT  7.570 3.260 7.790 3.880 ;
        RECT  5.870 3.320 7.570 3.880 ;
        RECT  5.590 3.260 5.870 3.880 ;
        RECT  2.930 3.320 5.590 3.880 ;
        RECT  2.650 3.260 2.930 3.880 ;
        RECT  0.890 3.320 2.650 3.880 ;
        RECT  0.610 3.260 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.660 1.520 8.960 1.680 ;
        RECT  8.500 1.520 8.660 3.100 ;
        RECT  7.760 2.940 8.500 3.100 ;
        RECT  7.600 2.680 7.760 3.100 ;
        RECT  6.730 2.680 7.600 2.840 ;
        RECT  6.190 3.000 7.390 3.160 ;
        RECT  7.210 0.830 7.370 0.990 ;
        RECT  7.050 0.500 7.210 2.390 ;
        RECT  5.530 0.500 7.050 0.660 ;
        RECT  6.730 0.910 6.890 1.070 ;
        RECT  6.570 0.910 6.730 2.840 ;
        RECT  6.250 0.820 6.410 2.270 ;
        RECT  6.190 0.820 6.250 1.100 ;
        RECT  6.090 2.110 6.250 2.390 ;
        RECT  5.250 0.820 6.190 0.980 ;
        RECT  6.030 2.940 6.190 3.160 ;
        RECT  5.930 1.520 6.090 1.800 ;
        RECT  4.970 2.940 6.030 3.100 ;
        RECT  5.290 1.520 5.930 1.680 ;
        RECT  5.390 0.440 5.530 0.660 ;
        RECT  5.290 1.140 5.510 1.300 ;
        RECT  3.760 0.440 5.390 0.600 ;
        RECT  5.130 1.140 5.290 2.780 ;
        RECT  5.110 0.760 5.250 0.980 ;
        RECT  4.170 0.760 5.110 0.920 ;
        RECT  4.810 1.080 4.970 3.100 ;
        RECT  4.390 2.780 4.810 2.940 ;
        RECT  4.490 1.200 4.650 2.620 ;
        RECT  4.330 1.080 4.490 1.360 ;
        RECT  4.130 2.460 4.490 2.620 ;
        RECT  4.170 1.700 4.330 1.980 ;
        RECT  4.010 0.760 4.170 2.300 ;
        RECT  3.970 2.460 4.130 2.920 ;
        RECT  3.650 2.140 4.010 2.300 ;
        RECT  2.450 2.760 3.970 2.920 ;
        RECT  3.690 1.700 3.850 1.980 ;
        RECT  3.600 0.440 3.760 1.260 ;
        RECT  3.440 1.700 3.690 1.920 ;
        RECT  3.490 2.140 3.650 2.600 ;
        RECT  3.590 0.440 3.600 0.920 ;
        RECT  2.160 0.760 3.590 0.920 ;
        RECT  2.400 2.440 3.490 2.600 ;
        RECT  3.280 1.090 3.440 1.920 ;
        RECT  2.350 1.090 3.280 1.250 ;
        RECT  2.720 2.120 3.230 2.280 ;
        RECT  2.560 2.040 2.720 2.280 ;
        RECT  2.350 2.040 2.560 2.200 ;
        RECT  2.290 2.760 2.450 3.160 ;
        RECT  2.240 2.360 2.400 2.600 ;
        RECT  2.190 1.090 2.350 2.200 ;
        RECT  1.210 3.000 2.290 3.160 ;
        RECT  2.030 2.360 2.240 2.520 ;
        RECT  2.130 1.090 2.190 1.250 ;
        RECT  2.030 0.710 2.160 0.920 ;
        RECT  1.530 2.680 2.070 2.840 ;
        RECT  1.550 0.710 2.030 0.870 ;
        RECT  1.870 1.410 2.030 2.520 ;
        RECT  1.710 1.030 1.870 1.570 ;
        RECT  1.550 1.730 1.710 2.200 ;
        RECT  1.390 0.710 1.550 1.890 ;
        RECT  1.370 2.410 1.530 2.840 ;
        RECT  1.230 2.410 1.370 2.570 ;
        RECT  1.070 1.030 1.230 2.570 ;
        RECT  1.050 2.940 1.210 3.160 ;
        RECT  0.310 2.940 1.050 3.100 ;
        RECT  0.830 1.360 0.910 1.640 ;
        RECT  0.670 0.520 0.830 2.480 ;
        RECT  0.090 0.520 0.670 0.680 ;
        RECT  0.310 2.320 0.670 2.480 ;
        RECT  0.150 2.320 0.310 3.160 ;
    END
END CMPR32X4TR

MACRO CMPR32X2TR
    CLASS CORE ;
    FOREIGN CMPR32X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.610 1.080 8.720 2.450 ;
        RECT  8.450 0.440 8.610 3.130 ;
        RECT  8.330 0.440 8.450 1.240 ;
        RECT  8.330 1.970 8.450 3.130 ;
        END
        ANTENNADIFFAREA 3.392 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 0.440 7.590 2.060 ;
        RECT  7.280 1.640 7.430 2.060 ;
        END
        ANTENNADIFFAREA 2.838 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.510 2.160 5.920 2.760 ;
        END
        ANTENNAGATEAREA 0.1992 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.430 0.530 1.720 ;
        RECT  0.320 1.430 0.340 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.440 3.120 2.050 ;
        RECT  2.570 1.440 2.880 1.600 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.130 -0.280 8.800 0.280 ;
        RECT  7.850 -0.280 8.130 1.240 ;
        RECT  6.050 -0.280 7.850 0.280 ;
        RECT  5.770 -0.280 6.050 0.340 ;
        RECT  2.930 -0.280 5.770 0.280 ;
        RECT  2.650 -0.280 2.930 0.600 ;
        RECT  0.890 -0.280 2.650 0.280 ;
        RECT  0.610 -0.280 0.890 0.300 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.130 3.320 8.800 3.880 ;
        RECT  7.850 2.570 8.130 3.880 ;
        RECT  5.910 3.320 7.850 3.880 ;
        RECT  5.630 3.260 5.910 3.880 ;
        RECT  2.930 3.320 5.630 3.880 ;
        RECT  2.650 3.260 2.930 3.880 ;
        RECT  0.890 3.320 2.650 3.880 ;
        RECT  0.610 3.260 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.130 1.530 8.270 1.810 ;
        RECT  7.970 1.530 8.130 2.380 ;
        RECT  7.630 2.220 7.970 2.380 ;
        RECT  7.470 2.220 7.630 2.840 ;
        RECT  6.770 2.680 7.470 2.840 ;
        RECT  6.230 3.000 7.440 3.160 ;
        RECT  7.090 2.360 7.310 2.520 ;
        RECT  7.090 1.020 7.210 1.180 ;
        RECT  6.930 0.500 7.090 2.520 ;
        RECT  5.490 0.500 6.930 0.660 ;
        RECT  6.610 0.900 6.770 2.840 ;
        RECT  6.510 0.900 6.610 1.180 ;
        RECT  6.260 1.330 6.420 2.590 ;
        RECT  6.190 1.330 6.260 1.490 ;
        RECT  6.130 2.300 6.260 2.590 ;
        RECT  6.070 2.940 6.230 3.160 ;
        RECT  6.030 0.820 6.190 1.490 ;
        RECT  5.940 1.650 6.100 1.930 ;
        RECT  5.010 2.940 6.070 3.100 ;
        RECT  5.210 0.820 6.030 0.980 ;
        RECT  5.330 1.650 5.940 1.810 ;
        RECT  5.350 0.440 5.490 0.660 ;
        RECT  5.330 1.140 5.490 1.300 ;
        RECT  3.790 0.440 5.350 0.600 ;
        RECT  5.170 1.140 5.330 2.780 ;
        RECT  5.060 0.760 5.210 0.980 ;
        RECT  4.150 0.760 5.060 0.920 ;
        RECT  4.850 1.140 5.010 3.100 ;
        RECT  4.730 1.140 4.850 2.940 ;
        RECT  4.390 2.780 4.730 2.940 ;
        RECT  4.470 1.200 4.570 2.620 ;
        RECT  4.410 1.080 4.470 2.620 ;
        RECT  4.310 1.080 4.410 1.360 ;
        RECT  4.130 2.460 4.410 2.620 ;
        RECT  4.150 1.700 4.250 1.980 ;
        RECT  3.990 0.760 4.150 2.300 ;
        RECT  3.970 2.460 4.130 3.010 ;
        RECT  3.650 2.140 3.990 2.300 ;
        RECT  2.450 2.850 3.970 3.010 ;
        RECT  3.470 1.700 3.830 1.980 ;
        RECT  3.630 0.440 3.790 1.250 ;
        RECT  3.490 2.140 3.650 2.690 ;
        RECT  2.160 0.760 3.630 0.920 ;
        RECT  2.400 2.530 3.490 2.690 ;
        RECT  3.310 1.090 3.470 1.980 ;
        RECT  2.350 1.090 3.310 1.250 ;
        RECT  2.720 2.210 3.250 2.370 ;
        RECT  2.560 2.030 2.720 2.370 ;
        RECT  2.350 2.030 2.560 2.190 ;
        RECT  2.290 2.850 2.450 3.150 ;
        RECT  2.240 2.350 2.400 2.690 ;
        RECT  2.190 1.090 2.350 2.190 ;
        RECT  1.210 2.990 2.290 3.150 ;
        RECT  2.030 2.350 2.240 2.510 ;
        RECT  2.130 1.090 2.190 1.250 ;
        RECT  2.030 0.710 2.160 0.920 ;
        RECT  1.710 2.670 2.080 2.830 ;
        RECT  1.550 0.710 2.030 0.870 ;
        RECT  1.870 1.390 2.030 2.510 ;
        RECT  1.710 1.030 1.870 1.550 ;
        RECT  1.550 1.710 1.710 2.190 ;
        RECT  1.550 2.510 1.710 2.830 ;
        RECT  1.390 0.710 1.550 1.870 ;
        RECT  1.230 2.510 1.550 2.670 ;
        RECT  1.070 1.030 1.230 2.670 ;
        RECT  1.050 2.940 1.210 3.150 ;
        RECT  0.310 2.940 1.050 3.100 ;
        RECT  0.850 1.360 0.910 1.640 ;
        RECT  0.690 0.460 0.850 2.420 ;
        RECT  0.090 0.460 0.690 0.680 ;
        RECT  0.310 2.260 0.690 2.420 ;
        RECT  0.150 2.260 0.310 3.160 ;
    END
END CMPR32X2TR

MACRO CMPR22X4TR
    CLASS CORE ;
    FOREIGN CMPR22X4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.670 0.500 7.950 0.780 ;
        RECT  6.990 0.500 7.670 0.660 ;
        RECT  7.280 1.840 7.520 2.720 ;
        RECT  7.190 1.960 7.280 2.720 ;
        RECT  6.510 1.960 7.190 2.120 ;
        RECT  6.710 0.500 6.990 0.780 ;
        RECT  6.030 0.500 6.710 0.660 ;
        RECT  6.190 1.960 6.510 2.840 ;
        RECT  5.550 2.120 6.190 2.280 ;
        RECT  5.750 0.500 6.030 1.460 ;
        RECT  5.070 1.300 5.750 1.460 ;
        RECT  5.270 2.120 5.550 2.400 ;
        RECT  4.590 2.120 5.270 2.280 ;
        RECT  4.790 1.030 5.070 1.460 ;
        RECT  4.110 1.300 4.790 1.460 ;
        RECT  4.310 2.120 4.590 2.400 ;
        RECT  3.630 2.120 4.310 2.340 ;
        RECT  3.830 1.030 4.110 1.460 ;
        RECT  3.120 1.300 3.830 1.460 ;
        RECT  3.120 2.060 3.630 2.340 ;
        RECT  2.960 1.300 3.120 2.340 ;
        END
        ANTENNADIFFAREA 17.714 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.880 0.770 13.120 2.490 ;
        RECT  12.310 0.770 12.880 1.000 ;
        RECT  12.320 2.240 12.880 2.490 ;
        RECT  12.030 2.240 12.320 3.160 ;
        RECT  12.030 0.440 12.310 1.000 ;
        END
        ANTENNADIFFAREA 3.96 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.990 1.440 7.590 1.600 ;
        RECT  6.780 1.440 6.990 1.800 ;
        RECT  4.360 1.640 6.780 1.800 ;
        RECT  4.040 1.640 4.360 1.960 ;
        RECT  3.280 1.640 4.040 1.900 ;
        END
        ANTENNAGATEAREA 1.6608 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.760 1.480 10.590 1.760 ;
        RECT  8.480 1.240 8.760 1.760 ;
        END
        ANTENNAGATEAREA 1.632 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.790 -0.280 13.200 0.280 ;
        RECT  12.510 -0.280 12.790 0.610 ;
        RECT  11.830 -0.280 12.510 0.280 ;
        RECT  11.550 -0.280 11.830 0.680 ;
        RECT  11.010 -0.280 11.550 0.280 ;
        RECT  10.730 -0.280 11.010 1.000 ;
        RECT  10.050 -0.280 10.730 0.280 ;
        RECT  9.770 -0.280 10.050 1.000 ;
        RECT  9.090 -0.280 9.770 0.280 ;
        RECT  8.810 -0.280 9.090 1.080 ;
        RECT  2.050 -0.280 8.810 0.340 ;
        RECT  1.330 -0.280 2.050 0.280 ;
        RECT  1.050 -0.280 1.330 1.010 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.790 3.320 13.200 3.880 ;
        RECT  12.510 2.700 12.790 3.880 ;
        RECT  11.830 3.320 12.510 3.880 ;
        RECT  11.550 2.240 11.830 3.880 ;
        RECT  10.870 3.320 11.550 3.880 ;
        RECT  10.590 2.560 10.870 3.880 ;
        RECT  9.870 3.320 10.590 3.880 ;
        RECT  9.590 2.800 9.870 3.880 ;
        RECT  8.830 3.320 9.590 3.880 ;
        RECT  8.550 3.200 8.830 3.880 ;
        RECT  7.910 3.260 8.550 3.880 ;
        RECT  7.630 3.200 7.910 3.880 ;
        RECT  3.290 3.320 7.630 3.880 ;
        RECT  3.010 3.200 3.290 3.880 ;
        RECT  2.330 3.260 3.010 3.880 ;
        RECT  2.050 3.200 2.330 3.880 ;
        RECT  1.330 3.320 2.050 3.880 ;
        RECT  1.050 2.250 1.330 3.880 ;
        RECT  0.370 3.320 1.050 3.880 ;
        RECT  0.090 1.930 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.560 1.160 12.720 2.080 ;
        RECT  11.490 1.160 12.560 1.320 ;
        RECT  11.350 1.920 12.560 2.080 ;
        RECT  10.910 1.540 12.400 1.700 ;
        RECT  11.210 1.040 11.490 1.320 ;
        RECT  11.070 1.920 11.350 3.160 ;
        RECT  10.530 1.160 11.210 1.320 ;
        RECT  10.390 2.240 11.070 2.400 ;
        RECT  10.750 1.540 10.910 2.080 ;
        RECT  8.430 1.920 10.750 2.080 ;
        RECT  10.250 0.440 10.530 1.320 ;
        RECT  10.110 2.240 10.390 3.160 ;
        RECT  9.570 1.160 10.250 1.320 ;
        RECT  9.350 2.240 10.110 2.400 ;
        RECT  9.290 0.440 9.570 1.320 ;
        RECT  9.070 2.240 9.350 3.040 ;
        RECT  7.910 2.880 9.070 3.040 ;
        RECT  8.310 1.920 8.430 2.720 ;
        RECT  8.150 1.040 8.310 2.720 ;
        RECT  8.070 1.040 8.150 1.320 ;
        RECT  7.750 1.060 7.910 3.040 ;
        RECT  7.470 1.060 7.750 1.220 ;
        RECT  6.990 2.880 7.750 3.040 ;
        RECT  7.190 0.940 7.470 1.220 ;
        RECT  6.510 1.060 7.190 1.220 ;
        RECT  6.710 2.280 6.990 3.160 ;
        RECT  6.030 3.000 6.710 3.160 ;
        RECT  6.230 0.940 6.510 1.220 ;
        RECT  5.750 2.560 6.030 3.160 ;
        RECT  2.130 2.560 5.750 2.720 ;
        RECT  5.270 0.500 5.550 1.140 ;
        RECT  4.590 0.500 5.270 0.660 ;
        RECT  4.790 2.880 5.070 3.160 ;
        RECT  4.110 2.880 4.790 3.040 ;
        RECT  4.310 0.500 4.590 1.140 ;
        RECT  1.810 0.500 4.310 0.660 ;
        RECT  3.830 2.880 4.110 3.160 ;
        RECT  1.810 2.880 3.830 3.040 ;
        RECT  2.730 0.820 3.670 1.100 ;
        RECT  2.450 0.820 2.730 2.190 ;
        RECT  1.970 1.490 2.130 2.720 ;
        RECT  1.010 1.490 1.970 1.770 ;
        RECT  1.530 0.500 1.810 1.330 ;
        RECT  1.530 1.930 1.810 3.040 ;
        RECT  0.850 1.170 1.530 1.330 ;
        RECT  0.850 1.930 1.530 2.090 ;
        RECT  0.570 0.440 0.850 3.160 ;
    END
END CMPR22X4TR

MACRO CMPR22X2TR
    CLASS CORE ;
    FOREIGN CMPR22X2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 0.800 4.630 1.080 ;
        RECT  4.240 1.780 4.520 2.240 ;
        RECT  3.670 0.920 4.350 1.080 ;
        RECT  3.600 1.780 4.240 1.940 ;
        RECT  3.390 0.440 3.670 1.080 ;
        RECT  3.280 1.780 3.600 2.780 ;
        RECT  2.710 0.920 3.390 1.080 ;
        RECT  2.680 2.060 3.280 2.220 ;
        RECT  2.680 0.760 2.710 1.080 ;
        RECT  2.520 0.760 2.680 2.220 ;
        RECT  2.430 0.760 2.520 1.040 ;
        RECT  2.270 1.940 2.520 2.220 ;
        END
        ANTENNADIFFAREA 10.3795 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.280 0.440 8.320 1.560 ;
        RECT  8.000 0.440 8.280 3.160 ;
        END
        ANTENNADIFFAREA 3.52 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.240 4.970 1.620 ;
        RECT  2.840 1.240 3.120 1.890 ;
        END
        ANTENNAGATEAREA 0.8424 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.920 1.630 6.290 1.910 ;
        RECT  5.450 1.630 5.920 1.960 ;
        END
        ANTENNAGATEAREA 0.8592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.830 -0.280 8.400 0.280 ;
        RECT  7.550 -0.280 7.830 0.860 ;
        RECT  6.850 -0.280 7.550 0.280 ;
        RECT  6.570 -0.280 6.850 0.800 ;
        RECT  1.570 -0.280 6.570 0.280 ;
        RECT  1.290 -0.280 1.570 0.380 ;
        RECT  0.570 -0.280 1.290 0.280 ;
        RECT  0.290 -0.280 0.570 1.310 ;
        RECT  0.000 -0.280 0.290 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 3.320 8.400 3.880 ;
        RECT  7.520 2.400 7.800 3.880 ;
        RECT  6.780 3.320 7.520 3.880 ;
        RECT  6.500 2.880 6.780 3.880 ;
        RECT  5.780 3.320 6.500 3.880 ;
        RECT  5.500 2.880 5.780 3.880 ;
        RECT  4.860 3.260 5.500 3.880 ;
        RECT  4.580 3.200 4.860 3.880 ;
        RECT  1.570 3.260 4.580 3.880 ;
        RECT  1.290 3.200 1.570 3.880 ;
        RECT  0.570 3.320 1.290 3.880 ;
        RECT  0.290 2.930 0.570 3.880 ;
        RECT  0.000 3.320 0.290 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.680 1.120 7.840 2.040 ;
        RECT  7.370 1.120 7.680 1.280 ;
        RECT  7.260 1.880 7.680 2.040 ;
        RECT  7.240 1.440 7.520 1.720 ;
        RECT  7.090 0.440 7.370 1.280 ;
        RECT  6.980 1.880 7.260 3.160 ;
        RECT  6.720 1.560 7.240 1.720 ;
        RECT  6.330 1.120 7.090 1.280 ;
        RECT  6.300 2.560 6.980 2.720 ;
        RECT  6.530 1.560 6.720 2.400 ;
        RECT  5.290 2.120 6.530 2.400 ;
        RECT  6.050 0.440 6.330 1.280 ;
        RECT  6.020 2.560 6.300 3.060 ;
        RECT  4.150 0.440 6.050 0.600 ;
        RECT  4.840 2.560 6.020 2.720 ;
        RECT  5.130 0.920 5.290 2.400 ;
        RECT  5.090 0.920 5.130 1.080 ;
        RECT  4.810 0.800 5.090 1.080 ;
        RECT  4.680 2.560 4.840 3.040 ;
        RECT  4.040 2.880 4.680 3.040 ;
        RECT  3.870 0.440 4.150 0.720 ;
        RECT  3.760 2.100 4.040 3.100 ;
        RECT  1.890 2.940 3.760 3.100 ;
        RECT  2.910 0.440 3.190 0.720 ;
        RECT  2.750 2.380 3.030 2.660 ;
        RECT  1.890 0.440 2.910 0.600 ;
        RECT  1.570 2.380 2.750 2.540 ;
        RECT  2.090 1.260 2.360 1.540 ;
        RECT  1.810 0.860 2.090 2.210 ;
        RECT  1.730 0.440 1.890 0.700 ;
        RECT  1.730 2.700 1.890 3.100 ;
        RECT  1.570 0.540 1.730 0.700 ;
        RECT  0.890 2.700 1.730 2.860 ;
        RECT  1.410 0.540 1.570 2.540 ;
        RECT  1.050 0.540 1.410 0.700 ;
        RECT  0.770 2.040 1.410 2.320 ;
        RECT  0.610 1.600 1.250 1.880 ;
        RECT  0.770 0.440 1.050 1.310 ;
        RECT  0.730 2.480 0.890 2.860 ;
        RECT  0.610 2.480 0.730 2.640 ;
        RECT  0.450 1.600 0.610 2.640 ;
    END
END CMPR22X2TR

MACRO ACHCONX4TR
    CLASS CORE ;
    FOREIGN ACHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.520 0.950 7.760 1.310 ;
        RECT  7.460 0.950 7.520 2.040 ;
        RECT  7.280 0.950 7.460 2.500 ;
        RECT  6.800 0.950 7.280 1.200 ;
        RECT  7.180 1.800 7.280 2.500 ;
        RECT  6.600 2.340 7.180 2.500 ;
        RECT  6.520 0.440 6.800 1.200 ;
        RECT  6.440 2.340 6.600 3.160 ;
        RECT  6.220 2.880 6.440 3.160 ;
        END
        ANTENNADIFFAREA 7.35 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 1.240 8.660 1.640 ;
        END
        ANTENNAGATEAREA 0.504 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 1.570 5.320 1.960 ;
        END
        ANTENNAGATEAREA 1.056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.100 -0.280 9.200 0.280 ;
        RECT  8.820 -0.280 9.100 0.670 ;
        RECT  8.100 -0.280 8.820 0.280 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  5.520 -0.280 7.820 0.280 ;
        RECT  5.240 -0.280 5.520 0.400 ;
        RECT  0.890 -0.280 5.240 0.280 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.940 3.320 9.200 3.880 ;
        RECT  8.640 2.290 8.940 3.880 ;
        RECT  7.920 3.320 8.640 3.880 ;
        RECT  7.640 3.180 7.920 3.880 ;
        RECT  5.480 3.320 7.640 3.880 ;
        RECT  5.200 2.930 5.480 3.880 ;
        RECT  0.850 3.320 5.200 3.880 ;
        RECT  0.570 2.990 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.860 0.870 9.020 2.070 ;
        RECT  8.620 0.870 8.860 1.030 ;
        RECT  8.440 1.910 8.860 2.070 ;
        RECT  8.340 0.560 8.620 1.030 ;
        RECT  8.160 1.910 8.440 2.970 ;
        RECT  7.280 0.560 8.340 0.720 ;
        RECT  6.980 2.660 8.160 2.820 ;
        RECT  7.000 0.440 7.280 0.720 ;
        RECT  6.810 1.360 7.090 1.640 ;
        RECT  6.760 2.660 6.980 2.940 ;
        RECT  6.360 1.360 6.810 1.520 ;
        RECT  6.530 1.680 6.650 1.960 ;
        RECT  6.370 1.680 6.530 2.180 ;
        RECT  6.280 2.020 6.370 2.180 ;
        RECT  6.200 0.600 6.360 1.520 ;
        RECT  6.120 2.020 6.280 2.720 ;
        RECT  4.540 0.600 6.200 0.760 ;
        RECT  6.160 1.360 6.200 1.520 ;
        RECT  5.880 1.360 6.160 1.860 ;
        RECT  5.010 2.560 6.120 2.720 ;
        RECT  5.760 0.920 6.040 1.200 ;
        RECT  5.720 2.020 5.960 2.300 ;
        RECT  5.720 1.040 5.760 1.200 ;
        RECT  5.560 1.040 5.720 2.300 ;
        RECT  4.850 2.560 5.010 3.100 ;
        RECT  4.720 0.960 5.000 1.340 ;
        RECT  4.720 2.120 5.000 2.280 ;
        RECT  1.780 2.940 4.850 3.100 ;
        RECT  4.560 1.180 4.720 2.280 ;
        RECT  4.400 2.620 4.620 2.780 ;
        RECT  4.260 0.600 4.540 1.020 ;
        RECT  4.240 1.240 4.400 2.780 ;
        RECT  3.620 0.600 4.260 0.760 ;
        RECT  4.060 1.240 4.240 1.400 ;
        RECT  2.100 2.620 4.240 2.780 ;
        RECT  3.900 1.560 4.080 2.320 ;
        RECT  3.900 0.980 4.060 1.400 ;
        RECT  3.780 0.980 3.900 1.260 ;
        RECT  3.620 1.560 3.900 1.720 ;
        RECT  2.820 2.300 3.660 2.460 ;
        RECT  3.460 0.600 3.620 1.720 ;
        RECT  3.300 0.800 3.460 1.080 ;
        RECT  2.820 0.610 2.940 1.260 ;
        RECT  2.660 0.450 2.820 2.460 ;
        RECT  1.210 0.450 2.660 0.610 ;
        RECT  2.270 2.240 2.660 2.460 ;
        RECT  2.180 0.770 2.460 1.050 ;
        RECT  1.540 0.770 2.180 0.930 ;
        RECT  1.940 2.280 2.100 2.780 ;
        RECT  1.870 1.090 1.980 1.250 ;
        RECT  1.870 2.280 1.940 2.440 ;
        RECT  1.710 1.090 1.870 2.440 ;
        RECT  1.620 2.600 1.780 3.100 ;
        RECT  1.700 1.090 1.710 1.250 ;
        RECT  1.280 2.280 1.710 2.440 ;
        RECT  0.960 2.600 1.620 2.760 ;
        RECT  1.380 0.770 1.540 1.980 ;
        RECT  0.960 1.820 1.380 1.980 ;
        RECT  1.120 2.140 1.280 2.440 ;
        RECT  1.050 0.450 1.210 0.720 ;
        RECT  0.370 0.560 1.050 0.720 ;
        RECT  0.640 1.380 1.000 1.660 ;
        RECT  0.800 1.820 0.960 2.760 ;
        RECT  0.480 0.920 0.640 2.700 ;
        RECT  0.370 0.920 0.480 1.080 ;
        RECT  0.370 2.540 0.480 2.700 ;
        RECT  0.090 0.560 0.370 1.080 ;
        RECT  0.090 2.540 0.370 3.160 ;
    END
END ACHCONX4TR

MACRO ACHCONX2TR
    CLASS CORE ;
    FOREIGN ACHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 0.920 7.120 2.360 ;
        RECT  6.960 0.920 7.040 2.500 ;
        RECT  6.570 0.920 6.960 1.080 ;
        RECT  6.880 2.040 6.960 2.500 ;
        RECT  6.450 2.340 6.880 2.500 ;
        RECT  6.390 0.800 6.570 1.080 ;
        RECT  6.290 2.340 6.450 2.830 ;
        RECT  6.020 2.670 6.290 2.830 ;
        END
        ANTENNADIFFAREA 3.993 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.040 7.520 1.760 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.420 2.320 1.960 ;
        END
        ANTENNAGATEAREA 1.0056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.130 0.720 1.740 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.620 -0.280 8.000 0.280 ;
        RECT  7.350 -0.280 7.620 0.400 ;
        RECT  5.360 -0.280 7.350 0.280 ;
        RECT  5.070 -0.280 5.360 0.340 ;
        RECT  0.830 -0.280 5.070 0.280 ;
        RECT  0.670 -0.280 0.830 0.400 ;
        RECT  0.000 -0.280 0.670 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.370 3.320 8.000 3.880 ;
        RECT  7.070 3.130 7.370 3.880 ;
        RECT  5.360 3.320 7.070 3.880 ;
        RECT  5.040 2.930 5.360 3.880 ;
        RECT  0.800 3.320 5.040 3.880 ;
        RECT  0.640 2.490 0.800 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.680 0.600 7.840 2.820 ;
        RECT  7.050 0.600 7.680 0.760 ;
        RECT  6.770 2.660 7.680 2.820 ;
        RECT  6.870 0.480 7.050 0.760 ;
        RECT  6.620 1.240 6.780 1.640 ;
        RECT  6.610 2.660 6.770 2.940 ;
        RECT  6.230 1.240 6.620 1.400 ;
        RECT  6.210 1.570 6.370 2.180 ;
        RECT  6.070 0.500 6.230 1.400 ;
        RECT  6.130 2.020 6.210 2.180 ;
        RECT  5.970 2.020 6.130 2.510 ;
        RECT  4.260 0.500 6.070 0.660 ;
        RECT  5.970 1.240 6.070 1.400 ;
        RECT  5.810 1.240 5.970 1.860 ;
        RECT  5.230 2.350 5.970 2.510 ;
        RECT  5.650 0.910 5.890 1.070 ;
        RECT  5.650 2.020 5.810 2.180 ;
        RECT  5.490 0.910 5.650 2.180 ;
        RECT  5.070 2.350 5.230 2.770 ;
        RECT  4.800 2.610 5.070 2.770 ;
        RECT  4.640 2.610 4.800 3.110 ;
        RECT  4.570 0.930 4.730 2.380 ;
        RECT  1.120 2.950 4.640 3.110 ;
        RECT  4.210 1.250 4.570 1.560 ;
        RECT  4.210 2.630 4.430 2.790 ;
        RECT  4.100 0.500 4.260 1.000 ;
        RECT  4.050 1.800 4.210 2.790 ;
        RECT  3.420 0.500 4.100 0.660 ;
        RECT  3.890 1.390 4.050 1.960 ;
        RECT  1.790 2.630 4.050 2.790 ;
        RECT  3.780 1.390 3.890 1.550 ;
        RECT  3.730 2.190 3.890 2.470 ;
        RECT  3.620 0.820 3.780 1.550 ;
        RECT  3.570 1.710 3.730 2.470 ;
        RECT  3.420 1.710 3.570 1.870 ;
        RECT  3.240 0.500 3.420 1.870 ;
        RECT  3.250 2.170 3.410 2.460 ;
        RECT  2.820 2.300 3.250 2.460 ;
        RECT  3.080 0.760 3.240 1.170 ;
        RECT  2.660 0.450 2.820 2.460 ;
        RECT  1.150 0.450 2.660 0.610 ;
        RECT  2.220 2.300 2.660 2.460 ;
        RECT  2.180 0.770 2.340 1.050 ;
        RECT  1.470 0.770 2.180 0.930 ;
        RECT  1.790 1.090 1.920 1.250 ;
        RECT  1.630 1.090 1.790 2.790 ;
        RECT  1.280 2.500 1.630 2.790 ;
        RECT  1.310 0.770 1.470 2.190 ;
        RECT  1.120 2.030 1.310 2.190 ;
        RECT  0.990 0.450 1.150 1.660 ;
        RECT  0.960 2.030 1.120 3.110 ;
        RECT  0.250 0.620 0.990 0.780 ;
        RECT  0.250 1.900 0.320 2.990 ;
        RECT  0.090 0.620 0.250 2.990 ;
    END
END ACHCONX2TR

MACRO ACHCINX4TR
    CLASS CORE ;
    FOREIGN ACHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.520 0.950 7.760 1.310 ;
        RECT  7.460 0.950 7.520 2.040 ;
        RECT  7.280 0.950 7.460 2.500 ;
        RECT  6.800 0.950 7.280 1.200 ;
        RECT  7.180 1.800 7.280 2.500 ;
        RECT  6.600 2.340 7.180 2.500 ;
        RECT  6.520 0.440 6.800 1.200 ;
        RECT  6.440 2.340 6.600 3.160 ;
        RECT  6.220 2.880 6.440 3.160 ;
        END
        ANTENNADIFFAREA 7.35 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 1.240 8.660 1.640 ;
        END
        ANTENNAGATEAREA 0.504 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.080 1.450 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.7896 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.100 -0.280 9.200 0.280 ;
        RECT  8.820 -0.280 9.100 0.670 ;
        RECT  8.100 -0.280 8.820 0.280 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  5.520 -0.280 7.820 0.280 ;
        RECT  5.240 -0.280 5.520 0.400 ;
        RECT  0.890 -0.280 5.240 0.280 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.940 3.320 9.200 3.880 ;
        RECT  8.640 2.290 8.940 3.880 ;
        RECT  7.920 3.320 8.640 3.880 ;
        RECT  7.640 3.180 7.920 3.880 ;
        RECT  5.480 3.320 7.640 3.880 ;
        RECT  5.200 2.930 5.480 3.880 ;
        RECT  0.850 3.320 5.200 3.880 ;
        RECT  0.570 2.990 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.860 0.870 9.020 2.070 ;
        RECT  8.620 0.870 8.860 1.030 ;
        RECT  8.440 1.910 8.860 2.070 ;
        RECT  8.340 0.560 8.620 1.030 ;
        RECT  8.160 1.910 8.440 2.970 ;
        RECT  7.280 0.560 8.340 0.720 ;
        RECT  6.980 2.660 8.160 2.820 ;
        RECT  7.000 0.440 7.280 0.720 ;
        RECT  6.810 1.360 7.090 1.640 ;
        RECT  6.760 2.660 6.980 2.940 ;
        RECT  6.360 1.360 6.810 1.520 ;
        RECT  6.530 1.680 6.650 1.960 ;
        RECT  6.370 1.680 6.530 2.180 ;
        RECT  6.280 2.020 6.370 2.180 ;
        RECT  6.200 0.600 6.360 1.520 ;
        RECT  6.120 2.020 6.280 2.720 ;
        RECT  4.460 0.600 6.200 0.760 ;
        RECT  6.100 1.360 6.200 1.520 ;
        RECT  4.970 2.560 6.120 2.720 ;
        RECT  5.940 1.360 6.100 1.860 ;
        RECT  5.780 0.920 6.040 1.200 ;
        RECT  5.780 2.020 5.960 2.300 ;
        RECT  5.760 0.920 5.780 2.300 ;
        RECT  5.620 1.040 5.760 2.300 ;
        RECT  5.300 1.540 5.460 2.280 ;
        RECT  4.740 2.120 5.300 2.280 ;
        RECT  4.810 2.560 4.970 3.100 ;
        RECT  4.740 0.960 4.920 1.340 ;
        RECT  1.780 2.940 4.810 3.100 ;
        RECT  4.640 0.960 4.740 2.280 ;
        RECT  4.580 1.180 4.640 2.280 ;
        RECT  4.360 2.620 4.580 2.780 ;
        RECT  4.180 0.600 4.460 1.020 ;
        RECT  4.200 1.240 4.360 2.780 ;
        RECT  3.980 1.240 4.200 1.400 ;
        RECT  2.100 2.620 4.200 2.780 ;
        RECT  3.540 0.600 4.180 0.760 ;
        RECT  4.020 2.040 4.040 2.320 ;
        RECT  3.860 1.560 4.020 2.320 ;
        RECT  3.820 0.980 3.980 1.400 ;
        RECT  3.540 1.560 3.860 1.720 ;
        RECT  3.700 0.980 3.820 1.260 ;
        RECT  2.820 2.300 3.620 2.460 ;
        RECT  3.380 0.600 3.540 1.720 ;
        RECT  3.220 0.800 3.380 1.080 ;
        RECT  2.820 0.610 2.940 1.260 ;
        RECT  2.660 0.450 2.820 2.460 ;
        RECT  1.210 0.450 2.660 0.610 ;
        RECT  2.270 2.240 2.660 2.460 ;
        RECT  2.180 0.770 2.460 1.050 ;
        RECT  1.540 0.770 2.180 0.930 ;
        RECT  1.940 2.280 2.100 2.780 ;
        RECT  1.870 1.090 1.980 1.250 ;
        RECT  1.870 2.280 1.940 2.440 ;
        RECT  1.710 1.090 1.870 2.440 ;
        RECT  1.620 2.600 1.780 3.100 ;
        RECT  1.700 1.090 1.710 1.250 ;
        RECT  1.280 2.280 1.710 2.440 ;
        RECT  0.960 2.600 1.620 2.760 ;
        RECT  1.380 0.770 1.540 1.980 ;
        RECT  0.960 1.820 1.380 1.980 ;
        RECT  1.120 2.140 1.280 2.440 ;
        RECT  1.050 0.450 1.210 0.720 ;
        RECT  0.370 0.560 1.050 0.720 ;
        RECT  0.640 1.380 1.000 1.660 ;
        RECT  0.800 1.820 0.960 2.760 ;
        RECT  0.480 0.920 0.640 2.700 ;
        RECT  0.370 0.920 0.480 1.080 ;
        RECT  0.370 2.540 0.480 2.700 ;
        RECT  0.090 0.560 0.370 1.080 ;
        RECT  0.090 2.540 0.370 3.160 ;
    END
END ACHCINX4TR

MACRO ACHCINX2TR
    CLASS CORE ;
    FOREIGN ACHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 0.920 7.120 2.360 ;
        RECT  6.960 0.920 7.040 2.500 ;
        RECT  6.550 0.920 6.960 1.080 ;
        RECT  6.880 2.040 6.960 2.500 ;
        RECT  6.450 2.340 6.880 2.500 ;
        RECT  6.390 0.800 6.550 1.080 ;
        RECT  6.290 2.340 6.450 2.830 ;
        RECT  6.020 2.670 6.290 2.830 ;
        END
        ANTENNADIFFAREA 3.993 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.280 1.040 7.520 1.760 ;
        END
        ANTENNAGATEAREA 0.2568 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.420 2.320 1.960 ;
        END
        ANTENNAGATEAREA 0.7392 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.130 0.720 1.740 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.550 -0.280 8.000 0.280 ;
        RECT  7.390 -0.280 7.550 0.400 ;
        RECT  5.360 -0.280 7.390 0.280 ;
        RECT  5.070 -0.280 5.360 0.340 ;
        RECT  0.830 -0.280 5.070 0.280 ;
        RECT  0.670 -0.280 0.830 0.400 ;
        RECT  0.000 -0.280 0.670 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.290 3.320 8.000 3.880 ;
        RECT  7.130 3.180 7.290 3.880 ;
        RECT  5.270 3.320 7.130 3.880 ;
        RECT  5.110 2.930 5.270 3.880 ;
        RECT  0.800 3.320 5.110 3.880 ;
        RECT  0.640 2.490 0.800 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.680 0.600 7.840 2.820 ;
        RECT  7.030 0.600 7.680 0.760 ;
        RECT  6.770 2.660 7.680 2.820 ;
        RECT  6.870 0.480 7.030 0.760 ;
        RECT  6.620 1.240 6.780 1.640 ;
        RECT  6.610 2.660 6.770 2.940 ;
        RECT  6.230 1.240 6.620 1.400 ;
        RECT  6.210 1.570 6.370 2.180 ;
        RECT  6.070 0.500 6.230 1.400 ;
        RECT  6.130 2.020 6.210 2.180 ;
        RECT  5.970 2.020 6.130 2.510 ;
        RECT  4.260 0.500 6.070 0.660 ;
        RECT  5.970 1.240 6.070 1.400 ;
        RECT  5.810 1.240 5.970 1.860 ;
        RECT  5.230 2.350 5.970 2.510 ;
        RECT  5.650 0.910 5.890 1.070 ;
        RECT  5.650 2.020 5.810 2.180 ;
        RECT  5.490 0.910 5.650 2.180 ;
        RECT  5.170 0.820 5.330 1.650 ;
        RECT  5.070 2.350 5.230 2.770 ;
        RECT  4.730 0.820 5.170 0.980 ;
        RECT  4.950 2.610 5.070 2.770 ;
        RECT  4.790 2.610 4.950 3.110 ;
        RECT  1.120 2.950 4.790 3.110 ;
        RECT  4.570 0.820 4.730 2.380 ;
        RECT  4.210 1.360 4.570 1.640 ;
        RECT  4.210 2.630 4.430 2.790 ;
        RECT  4.100 0.500 4.260 1.180 ;
        RECT  4.050 1.800 4.210 2.790 ;
        RECT  3.420 0.500 4.100 0.660 ;
        RECT  3.890 1.390 4.050 1.960 ;
        RECT  1.790 2.630 4.050 2.790 ;
        RECT  3.780 1.390 3.890 1.550 ;
        RECT  3.730 2.190 3.890 2.470 ;
        RECT  3.620 0.960 3.780 1.550 ;
        RECT  3.570 1.710 3.730 2.470 ;
        RECT  3.420 1.710 3.570 1.870 ;
        RECT  3.240 0.500 3.420 1.870 ;
        RECT  3.250 2.170 3.410 2.460 ;
        RECT  2.820 2.300 3.250 2.460 ;
        RECT  3.080 1.010 3.240 1.170 ;
        RECT  2.660 0.450 2.820 2.460 ;
        RECT  1.150 0.450 2.660 0.610 ;
        RECT  2.220 2.300 2.660 2.460 ;
        RECT  2.180 0.770 2.340 1.050 ;
        RECT  1.470 0.770 2.180 0.930 ;
        RECT  1.790 1.090 1.920 1.250 ;
        RECT  1.630 1.090 1.790 2.790 ;
        RECT  1.280 2.500 1.630 2.790 ;
        RECT  1.310 0.770 1.470 2.190 ;
        RECT  1.120 2.030 1.310 2.190 ;
        RECT  0.990 0.450 1.150 1.660 ;
        RECT  0.960 2.030 1.120 3.110 ;
        RECT  0.250 0.620 0.990 0.780 ;
        RECT  0.250 1.900 0.320 2.990 ;
        RECT  0.090 0.620 0.250 2.990 ;
    END
END ACHCINX2TR

MACRO ACCSIHCONX4TR
    CLASS CORE ;
    FOREIGN ACCSIHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.920 4.320 2.280 ;
        RECT  3.680 0.920 4.000 1.080 ;
        RECT  3.200 2.120 4.000 2.280 ;
        RECT  3.400 0.800 3.680 1.080 ;
        RECT  2.640 0.920 3.400 1.080 ;
        RECT  2.880 2.120 3.200 3.160 ;
        RECT  2.360 0.800 2.640 1.080 ;
        END
        ANTENNADIFFAREA 5.236 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 2.120 1.920 2.960 ;
        RECT  0.880 2.120 1.560 2.280 ;
        RECT  0.920 0.440 1.200 1.080 ;
        RECT  0.320 0.920 0.920 1.080 ;
        RECT  0.600 2.120 0.880 2.950 ;
        RECT  0.320 2.120 0.600 2.280 ;
        RECT  0.080 0.920 0.320 2.280 ;
        END
        ANTENNADIFFAREA 5.004 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.240 3.840 1.640 ;
        RECT  2.520 1.240 3.560 1.400 ;
        RECT  2.240 1.240 2.520 1.640 ;
        RECT  1.520 1.240 2.240 1.400 ;
        RECT  0.880 1.240 1.520 1.640 ;
        END
        ANTENNAGATEAREA 0.912 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.580 3.400 1.860 ;
        RECT  2.680 1.580 2.840 1.960 ;
        RECT  2.040 1.800 2.680 1.960 ;
        RECT  1.760 1.560 2.040 1.960 ;
        RECT  0.720 1.800 1.760 1.960 ;
        RECT  0.480 1.240 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.912 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.200 -0.280 4.400 0.280 ;
        RECT  3.920 -0.280 4.200 0.400 ;
        RECT  3.160 -0.280 3.920 0.340 ;
        RECT  2.880 -0.280 3.160 0.400 ;
        RECT  2.000 -0.280 2.880 0.340 ;
        RECT  1.720 -0.280 2.000 1.080 ;
        RECT  0.400 -0.280 1.720 0.280 ;
        RECT  0.120 -0.280 0.400 0.760 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.000 3.320 4.400 3.880 ;
        RECT  3.720 2.440 4.000 3.880 ;
        RECT  2.320 3.320 3.720 3.880 ;
        RECT  2.100 2.120 2.320 3.880 ;
        RECT  1.360 3.320 2.100 3.880 ;
        RECT  1.080 2.670 1.360 3.880 ;
        RECT  0.400 3.320 1.080 3.880 ;
        RECT  0.120 2.670 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END ACCSIHCONX4TR

MACRO ACCSIHCONX2TR
    CLASS CORE ;
    FOREIGN ACCSIHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 2.040 2.320 3.160 ;
        RECT  2.080 1.190 2.240 3.160 ;
        RECT  1.770 1.190 2.080 1.360 ;
        RECT  1.890 2.190 2.080 3.160 ;
        RECT  1.610 0.760 1.770 1.360 ;
        RECT  1.480 0.760 1.610 1.040 ;
        END
        ANTENNADIFFAREA 3.376 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 2.180 0.850 2.870 ;
        RECT  0.480 1.850 0.640 2.870 ;
        RECT  0.260 1.850 0.480 2.010 ;
        RECT  0.260 0.440 0.440 1.070 ;
        RECT  0.100 0.440 0.260 2.010 ;
        END
        ANTENNADIFFAREA 3.2 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.240 1.440 1.640 ;
        RECT  1.120 1.240 1.280 1.400 ;
        RECT  0.880 0.840 1.120 1.400 ;
        RECT  0.580 1.240 0.880 1.400 ;
        RECT  0.420 1.240 0.580 1.690 ;
        END
        ANTENNAGATEAREA 0.468 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.520 1.920 2.020 ;
        RECT  1.040 1.860 1.680 2.020 ;
        RECT  0.880 1.580 1.040 2.020 ;
        END
        ANTENNAGATEAREA 0.468 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 -0.280 2.400 0.280 ;
        RECT  1.960 -0.280 2.240 0.990 ;
        RECT  1.240 -0.280 1.960 0.280 ;
        RECT  0.960 -0.280 1.240 0.680 ;
        RECT  0.000 -0.280 0.960 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 3.320 2.400 3.880 ;
        RECT  1.090 2.450 1.370 3.880 ;
        RECT  0.310 3.260 1.090 3.880 ;
        RECT  0.090 2.170 0.310 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END ACCSIHCONX2TR

MACRO ACCSHCONX4TR
    CLASS CORE ;
    FOREIGN ACCSHCONX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.400 0.900 8.440 1.060 ;
        RECT  8.280 0.900 8.400 2.190 ;
        RECT  8.120 0.760 8.280 2.190 ;
        RECT  7.520 0.760 8.120 0.920 ;
        RECT  7.380 0.760 7.520 1.760 ;
        RECT  7.260 0.760 7.380 2.190 ;
        RECT  7.220 0.760 7.260 2.500 ;
        RECT  7.100 2.030 7.220 2.500 ;
        RECT  6.400 2.340 7.100 2.500 ;
        RECT  6.400 0.440 6.470 1.870 ;
        RECT  6.310 0.440 6.400 2.500 ;
        RECT  6.300 0.440 6.310 1.130 ;
        RECT  6.240 1.720 6.310 2.500 ;
        RECT  6.080 2.020 6.240 2.180 ;
        END
        ANTENNADIFFAREA 8.568 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.920 0.950 11.080 1.110 ;
        RECT  10.760 0.760 10.920 1.110 ;
        RECT  10.060 0.760 10.760 0.920 ;
        RECT  10.560 2.480 10.720 3.160 ;
        RECT  9.920 3.000 10.560 3.160 ;
        RECT  9.920 0.760 10.060 1.750 ;
        RECT  9.900 0.760 9.920 3.160 ;
        RECT  9.100 0.760 9.900 0.920 ;
        RECT  9.760 1.580 9.900 3.160 ;
        RECT  9.580 2.240 9.760 3.160 ;
        RECT  8.860 3.000 9.580 3.160 ;
        RECT  8.940 0.760 9.100 1.150 ;
        RECT  8.580 2.670 8.860 3.160 ;
        END
        ANTENNADIFFAREA 8.138 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.720 1.260 12.880 1.640 ;
        RECT  12.480 0.840 12.720 1.420 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.080 1.470 12.320 1.960 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.840 4.720 1.160 ;
        RECT  4.480 0.840 4.640 1.840 ;
        END
        ANTENNAGATEAREA 0.7824 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.240 0.560 2.360 ;
        END
        ANTENNAGATEAREA 0.5256 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.720 -0.280 14.000 0.280 ;
        RECT  13.560 -0.280 13.720 1.310 ;
        RECT  12.740 -0.280 13.560 0.280 ;
        RECT  12.460 -0.280 12.740 0.340 ;
        RECT  11.700 -0.280 12.460 0.280 ;
        RECT  11.420 -0.280 11.700 0.340 ;
        RECT  5.960 -0.280 11.420 0.280 ;
        RECT  5.680 -0.280 5.960 0.590 ;
        RECT  4.560 -0.280 5.680 0.280 ;
        RECT  4.400 -0.280 4.560 0.670 ;
        RECT  1.840 -0.280 4.400 0.280 ;
        RECT  1.560 -0.280 1.840 0.340 ;
        RECT  0.460 -0.280 1.560 0.280 ;
        RECT  0.180 -0.280 0.460 1.070 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.720 3.320 14.000 3.880 ;
        RECT  13.560 2.120 13.720 3.880 ;
        RECT  12.680 3.320 13.560 3.880 ;
        RECT  12.520 2.340 12.680 3.880 ;
        RECT  11.640 3.320 12.520 3.880 ;
        RECT  11.480 2.520 11.640 3.880 ;
        RECT  5.420 3.320 11.480 3.880 ;
        RECT  5.140 2.990 5.420 3.880 ;
        RECT  4.600 3.320 5.140 3.880 ;
        RECT  4.320 2.990 4.600 3.880 ;
        RECT  1.740 3.320 4.320 3.880 ;
        RECT  1.580 2.930 1.740 3.880 ;
        RECT  0.460 3.320 1.580 3.880 ;
        RECT  0.180 2.530 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.040 0.440 13.200 3.160 ;
        RECT  11.240 0.500 13.040 0.660 ;
        RECT  12.000 1.030 12.160 1.310 ;
        RECT  12.000 2.120 12.160 3.160 ;
        RECT  11.920 1.150 12.000 1.310 ;
        RECT  11.920 2.120 12.000 2.280 ;
        RECT  11.760 1.150 11.920 2.280 ;
        RECT  10.480 2.120 11.760 2.280 ;
        RECT  11.080 0.440 11.240 0.660 ;
        RECT  6.940 0.440 11.080 0.600 ;
        RECT  10.480 1.080 10.600 1.240 ;
        RECT  10.320 1.080 10.480 2.280 ;
        RECT  10.240 2.120 10.320 2.280 ;
        RECT  10.080 2.120 10.240 2.840 ;
        RECT  9.520 1.090 9.640 1.250 ;
        RECT  9.360 1.090 9.520 1.800 ;
        RECT  9.280 1.610 9.360 1.800 ;
        RECT  9.120 1.610 9.280 2.560 ;
        RECT  8.160 2.350 9.120 2.510 ;
        RECT  8.000 2.350 8.160 3.140 ;
        RECT  5.740 2.980 8.000 3.140 ;
        RECT  7.840 1.080 7.960 1.240 ;
        RECT  7.680 1.080 7.840 2.820 ;
        RECT  6.060 2.660 7.680 2.820 ;
        RECT  6.780 0.440 6.940 2.180 ;
        RECT  6.560 2.020 6.780 2.180 ;
        RECT  5.920 1.290 6.150 1.570 ;
        RECT  5.900 2.350 6.060 2.820 ;
        RECT  5.760 0.750 5.920 2.190 ;
        RECT  5.280 2.350 5.900 2.510 ;
        RECT  5.440 0.750 5.760 0.910 ;
        RECT  5.620 2.030 5.760 2.190 ;
        RECT  5.580 2.670 5.740 3.140 ;
        RECT  5.440 1.070 5.600 1.870 ;
        RECT  3.980 2.670 5.580 2.830 ;
        RECT  5.280 0.450 5.440 0.910 ;
        RECT  5.040 1.070 5.440 1.230 ;
        RECT  5.280 1.710 5.440 1.870 ;
        RECT  5.160 0.450 5.280 0.610 ;
        RECT  4.960 1.390 5.280 1.550 ;
        RECT  5.120 1.710 5.280 2.510 ;
        RECT  4.800 2.320 5.120 2.510 ;
        RECT  4.880 0.950 5.040 1.230 ;
        RECT  4.800 1.390 4.960 2.160 ;
        RECT  4.440 2.000 4.800 2.160 ;
        RECT  4.280 2.000 4.440 2.450 ;
        RECT  3.660 2.290 4.280 2.450 ;
        RECT  3.960 0.440 4.120 2.130 ;
        RECT  3.820 2.670 3.980 3.160 ;
        RECT  3.920 0.440 3.960 0.720 ;
        RECT  3.840 1.970 3.960 2.130 ;
        RECT  3.480 0.560 3.920 0.720 ;
        RECT  2.060 3.000 3.820 3.160 ;
        RECT  3.660 1.030 3.800 1.190 ;
        RECT  3.500 1.030 3.660 2.840 ;
        RECT  2.720 2.680 3.500 2.840 ;
        RECT  3.320 0.440 3.480 0.720 ;
        RECT  3.160 0.880 3.320 1.040 ;
        RECT  3.160 2.230 3.180 2.510 ;
        RECT  3.000 0.650 3.160 2.510 ;
        RECT  1.320 0.650 3.000 0.810 ;
        RECT  2.720 1.030 2.840 1.190 ;
        RECT  2.560 1.030 2.720 2.840 ;
        RECT  2.540 2.560 2.560 2.840 ;
        RECT  2.140 0.970 2.300 2.190 ;
        RECT  2.060 1.910 2.140 2.190 ;
        RECT  1.900 2.610 2.060 3.160 ;
        RECT  1.320 1.380 1.980 1.540 ;
        RECT  0.880 2.610 1.900 2.770 ;
        RECT  1.160 0.650 1.320 2.130 ;
        RECT  1.100 0.970 1.160 1.250 ;
        RECT  1.040 1.970 1.160 2.130 ;
        RECT  0.720 0.440 0.880 3.160 ;
    END
END ACCSHCONX4TR

MACRO ACCSHCONX2TR
    CLASS CORE ;
    FOREIGN ACCSHCONX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.960 0.840 8.120 1.120 ;
        RECT  7.800 0.760 7.960 2.460 ;
        RECT  7.160 0.760 7.800 0.920 ;
        RECT  7.680 2.300 7.800 2.460 ;
        RECT  7.000 0.760 7.160 1.760 ;
        RECT  6.840 0.840 7.000 2.190 ;
        RECT  6.720 1.970 6.840 2.190 ;
        END
        ANTENNADIFFAREA 4.83 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.440 0.870 9.560 3.100 ;
        RECT  9.280 0.770 9.440 3.100 ;
        RECT  8.600 0.770 9.280 0.930 ;
        RECT  9.240 2.230 9.280 3.100 ;
        RECT  8.240 2.940 9.240 3.100 ;
        RECT  8.440 0.770 8.600 1.250 ;
        RECT  8.320 0.870 8.440 1.250 ;
        END
        ANTENNADIFFAREA 5.208 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.480 1.240 10.720 1.960 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.040 1.240 10.320 1.680 ;
        END
        ANTENNAGATEAREA 0.2592 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 0.840 4.760 1.160 ;
        RECT  4.440 0.840 4.680 1.750 ;
        RECT  4.400 1.470 4.440 1.750 ;
        END
        ANTENNAGATEAREA 0.7824 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.640 1.640 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.5256 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.580 -0.280 11.200 0.280 ;
        RECT  10.300 -0.280 10.580 0.340 ;
        RECT  6.120 -0.280 10.300 0.280 ;
        RECT  5.840 -0.280 6.120 0.590 ;
        RECT  4.720 -0.280 5.840 0.280 ;
        RECT  4.440 -0.280 4.720 0.670 ;
        RECT  1.940 -0.280 4.440 0.280 ;
        RECT  1.660 -0.280 1.940 0.400 ;
        RECT  0.600 -0.280 1.660 0.280 ;
        RECT  0.320 -0.280 0.600 1.080 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.520 3.320 11.200 3.880 ;
        RECT  10.240 2.380 10.520 3.880 ;
        RECT  5.580 3.260 10.240 3.880 ;
        RECT  5.300 2.990 5.580 3.880 ;
        RECT  4.720 3.320 5.300 3.880 ;
        RECT  4.440 2.990 4.720 3.880 ;
        RECT  1.900 3.320 4.440 3.880 ;
        RECT  1.620 2.930 1.900 3.880 ;
        RECT  0.600 3.320 1.620 3.880 ;
        RECT  0.320 2.520 0.600 3.880 ;
        RECT  0.000 3.320 0.320 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.040 0.500 11.100 1.250 ;
        RECT  10.880 0.500 11.040 3.160 ;
        RECT  9.760 0.500 10.880 0.660 ;
        RECT  10.760 2.230 10.880 3.160 ;
        RECT  9.880 0.860 10.060 1.080 ;
        RECT  9.880 2.240 10.000 3.100 ;
        RECT  9.720 0.860 9.880 3.100 ;
        RECT  9.600 0.440 9.760 0.660 ;
        RECT  6.680 0.440 9.600 0.600 ;
        RECT  8.960 1.090 9.080 1.310 ;
        RECT  8.960 2.620 9.040 2.780 ;
        RECT  8.800 1.090 8.960 2.780 ;
        RECT  7.950 2.620 8.800 2.780 ;
        RECT  7.790 2.620 7.950 2.830 ;
        RECT  4.180 2.670 7.790 2.830 ;
        RECT  7.480 1.080 7.640 1.300 ;
        RECT  7.320 1.080 7.480 2.510 ;
        RECT  5.320 2.350 7.320 2.510 ;
        RECT  6.520 0.440 6.680 1.810 ;
        RECT  6.400 0.440 6.520 1.050 ;
        RECT  6.360 1.650 6.520 2.150 ;
        RECT  6.080 1.270 6.360 1.490 ;
        RECT  6.240 1.930 6.360 2.150 ;
        RECT  5.920 0.750 6.080 2.190 ;
        RECT  5.600 0.750 5.920 0.910 ;
        RECT  5.780 2.030 5.920 2.190 ;
        RECT  5.600 1.070 5.760 1.870 ;
        RECT  5.440 0.440 5.600 0.910 ;
        RECT  5.200 1.070 5.600 1.230 ;
        RECT  5.320 1.710 5.600 1.870 ;
        RECT  5.320 0.440 5.440 0.720 ;
        RECT  5.000 1.390 5.440 1.550 ;
        RECT  5.160 1.710 5.320 2.510 ;
        RECT  4.920 0.950 5.200 1.230 ;
        RECT  4.920 2.230 5.160 2.510 ;
        RECT  4.840 1.390 5.000 2.070 ;
        RECT  4.560 1.910 4.840 2.070 ;
        RECT  4.400 1.910 4.560 2.510 ;
        RECT  3.860 2.350 4.400 2.510 ;
        RECT  4.080 0.440 4.240 2.190 ;
        RECT  4.020 2.670 4.180 3.160 ;
        RECT  3.960 0.440 4.080 0.720 ;
        RECT  3.960 1.910 4.080 2.190 ;
        RECT  2.220 3.000 4.020 3.160 ;
        RECT  3.700 0.560 3.960 0.720 ;
        RECT  3.740 0.970 3.900 1.250 ;
        RECT  3.740 2.350 3.860 2.840 ;
        RECT  3.580 0.970 3.740 2.840 ;
        RECT  3.420 0.440 3.700 0.720 ;
        RECT  2.900 2.680 3.580 2.840 ;
        RECT  3.260 0.880 3.420 1.160 ;
        RECT  3.260 2.230 3.380 2.510 ;
        RECT  3.100 0.650 3.260 2.510 ;
        RECT  1.420 0.650 3.100 0.810 ;
        RECT  2.820 0.970 2.940 1.250 ;
        RECT  2.820 2.560 2.900 2.840 ;
        RECT  2.660 0.970 2.820 2.840 ;
        RECT  2.620 2.560 2.660 2.840 ;
        RECT  2.380 0.970 2.460 1.250 ;
        RECT  2.180 0.970 2.380 2.190 ;
        RECT  2.060 2.610 2.220 3.160 ;
        RECT  2.100 1.910 2.180 2.190 ;
        RECT  1.080 2.610 2.060 2.770 ;
        RECT  1.420 1.320 2.020 1.600 ;
        RECT  1.260 0.650 1.420 2.190 ;
        RECT  1.140 0.970 1.260 1.250 ;
        RECT  1.140 1.910 1.260 2.190 ;
        RECT  0.960 0.440 1.080 0.720 ;
        RECT  0.960 2.610 1.080 3.160 ;
        RECT  0.800 0.440 0.960 3.160 ;
    END
END ACCSHCONX2TR

MACRO ACCSHCINX4TR
    CLASS CORE ;
    FOREIGN ACCSHCINX4TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.250 0.970 10.450 1.250 ;
        RECT  10.170 0.970 10.250 2.510 ;
        RECT  10.090 1.090 10.170 2.510 ;
        RECT  9.970 2.270 10.090 2.510 ;
        RECT  8.530 2.350 9.970 2.510 ;
        RECT  9.490 0.640 9.520 1.360 ;
        RECT  9.270 0.440 9.490 1.750 ;
        RECT  8.530 1.590 9.270 1.750 ;
        RECT  8.370 1.590 8.530 2.510 ;
        RECT  8.080 1.590 8.370 2.080 ;
        END
        ANTENNADIFFAREA 9.786 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.050 2.290 13.330 3.160 ;
        RECT  12.730 1.090 13.050 1.360 ;
        RECT  12.370 3.000 13.050 3.160 ;
        RECT  12.370 1.200 12.730 1.360 ;
        RECT  12.090 1.200 12.370 3.160 ;
        RECT  12.050 1.030 12.090 3.160 ;
        RECT  11.810 1.030 12.050 1.360 ;
        RECT  11.410 3.000 12.050 3.160 ;
        RECT  11.250 2.290 11.410 3.160 ;
        RECT  11.130 2.290 11.250 2.890 ;
        END
        ANTENNADIFFAREA 7.056 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  16.080 1.240 16.320 2.360 ;
        RECT  15.830 1.240 16.080 1.750 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.440 1.240 14.760 1.660 ;
        END
        ANTENNAGATEAREA 0.5328 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.560 1.100 6.720 1.380 ;
        RECT  6.360 1.220 6.560 1.380 ;
        RECT  6.060 1.220 6.360 1.560 ;
        RECT  6.000 0.850 6.060 1.560 ;
        RECT  5.780 0.850 6.000 1.850 ;
        RECT  5.720 1.570 5.780 1.850 ;
        END
        ANTENNAGATEAREA 0.7824 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.240 0.490 1.630 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.310 -0.280 16.400 0.280 ;
        RECT  16.030 -0.280 16.310 1.080 ;
        RECT  15.350 -0.280 16.030 0.280 ;
        RECT  15.130 -0.280 15.350 0.760 ;
        RECT  14.130 -0.280 15.130 0.280 ;
        RECT  13.850 -0.280 14.130 0.320 ;
        RECT  8.780 -0.280 13.850 0.280 ;
        RECT  8.500 -0.280 8.780 0.400 ;
        RECT  7.860 -0.280 8.500 0.340 ;
        RECT  7.580 -0.280 7.860 0.390 ;
        RECT  6.340 -0.280 7.580 0.280 ;
        RECT  6.060 -0.280 6.340 0.370 ;
        RECT  0.890 -0.280 6.060 0.280 ;
        RECT  0.610 -0.280 0.890 0.400 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.310 3.320 16.400 3.880 ;
        RECT  16.030 2.530 16.310 3.880 ;
        RECT  15.350 3.320 16.030 3.880 ;
        RECT  15.070 1.910 15.350 3.880 ;
        RECT  14.390 3.320 15.070 3.880 ;
        RECT  14.110 2.290 14.390 3.880 ;
        RECT  7.530 3.320 14.110 3.880 ;
        RECT  6.600 3.260 7.530 3.880 ;
        RECT  1.710 3.320 6.600 3.880 ;
        RECT  1.430 3.180 1.710 3.880 ;
        RECT  0.370 3.320 1.430 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.670 0.440 15.830 1.080 ;
        RECT  15.670 1.910 15.830 3.160 ;
        RECT  15.510 0.440 15.670 3.160 ;
        RECT  14.970 0.920 15.510 1.080 ;
        RECT  14.810 0.480 14.970 1.080 ;
        RECT  14.590 1.910 14.870 3.160 ;
        RECT  13.690 0.480 14.810 0.640 ;
        RECT  14.280 0.800 14.650 1.080 ;
        RECT  14.280 1.910 14.590 2.130 ;
        RECT  14.120 0.800 14.280 2.130 ;
        RECT  13.370 0.800 14.120 0.960 ;
        RECT  13.810 1.970 14.120 2.130 ;
        RECT  13.530 1.970 13.810 2.920 ;
        RECT  13.530 0.440 13.690 0.640 ;
        RECT  9.970 0.440 13.530 0.600 ;
        RECT  12.850 1.970 13.530 2.130 ;
        RECT  13.210 0.760 13.370 0.960 ;
        RECT  12.570 0.760 13.210 0.920 ;
        RECT  12.690 1.970 12.850 2.840 ;
        RECT  12.570 2.290 12.690 2.840 ;
        RECT  12.290 0.760 12.570 1.040 ;
        RECT  11.770 2.290 11.890 2.840 ;
        RECT  11.610 1.520 11.770 2.840 ;
        RECT  11.330 0.760 11.610 1.680 ;
        RECT  10.770 0.760 11.330 0.920 ;
        RECT  10.950 1.350 11.150 1.890 ;
        RECT  10.930 1.350 10.950 3.150 ;
        RECT  10.730 1.730 10.930 3.150 ;
        RECT  10.610 0.760 10.770 1.570 ;
        RECT  7.850 2.990 10.730 3.150 ;
        RECT  10.570 1.410 10.610 1.570 ;
        RECT  10.410 1.410 10.570 2.830 ;
        RECT  8.210 2.670 10.410 2.830 ;
        RECT  9.840 0.440 9.970 0.720 ;
        RECT  9.680 0.440 9.840 2.070 ;
        RECT  8.910 1.910 9.680 2.070 ;
        RECT  8.890 0.560 9.110 1.430 ;
        RECT  8.690 1.910 8.910 2.190 ;
        RECT  7.420 0.560 8.890 0.720 ;
        RECT  7.540 0.880 8.260 1.040 ;
        RECT  8.050 2.240 8.210 2.830 ;
        RECT  6.690 2.240 8.050 2.400 ;
        RECT  5.560 2.560 7.890 2.780 ;
        RECT  7.690 2.940 7.850 3.150 ;
        RECT  5.880 2.940 7.690 3.100 ;
        RECT  7.260 0.880 7.540 2.080 ;
        RECT  7.260 0.450 7.420 0.720 ;
        RECT  6.660 0.450 7.260 0.610 ;
        RECT  6.850 1.860 7.260 2.080 ;
        RECT  6.940 0.770 7.100 1.700 ;
        RECT  6.820 0.770 6.940 0.930 ;
        RECT  6.690 1.540 6.940 1.700 ;
        RECT  6.530 1.540 6.690 2.400 ;
        RECT  6.500 0.450 6.660 0.690 ;
        RECT  5.970 2.120 6.530 2.400 ;
        RECT  5.620 0.530 6.500 0.690 ;
        RECT  5.720 2.940 5.880 3.160 ;
        RECT  5.560 2.010 5.720 2.290 ;
        RECT  2.030 3.000 5.720 3.160 ;
        RECT  5.560 0.530 5.620 1.040 ;
        RECT  5.440 0.530 5.560 2.290 ;
        RECT  5.400 2.560 5.560 2.840 ;
        RECT  5.400 0.530 5.440 2.170 ;
        RECT  4.600 0.530 5.400 0.690 ;
        RECT  2.350 2.620 5.400 2.840 ;
        RECT  5.140 1.920 5.240 2.200 ;
        RECT  5.020 0.900 5.140 2.200 ;
        RECT  4.860 0.900 5.020 2.460 ;
        RECT  2.670 2.300 4.860 2.460 ;
        RECT  4.600 1.980 4.700 2.140 ;
        RECT  4.440 0.530 4.600 2.140 ;
        RECT  4.320 0.760 4.440 1.040 ;
        RECT  4.420 1.980 4.440 2.140 ;
        RECT  4.120 1.920 4.220 2.140 ;
        RECT  3.940 0.440 4.120 2.140 ;
        RECT  2.800 0.440 3.940 0.720 ;
        RECT  2.950 1.920 3.940 2.140 ;
        RECT  2.490 1.020 3.650 1.300 ;
        RECT  1.210 0.440 2.800 0.600 ;
        RECT  2.510 2.080 2.670 2.460 ;
        RECT  2.230 2.080 2.510 2.240 ;
        RECT  2.330 0.760 2.490 1.300 ;
        RECT  2.190 2.400 2.350 2.840 ;
        RECT  1.690 0.760 2.330 0.920 ;
        RECT  2.130 1.960 2.230 2.240 ;
        RECT  1.690 2.400 2.190 2.560 ;
        RECT  1.970 1.080 2.130 2.240 ;
        RECT  1.870 2.860 2.030 3.160 ;
        RECT  1.850 1.080 1.970 1.300 ;
        RECT  1.950 1.960 1.970 2.240 ;
        RECT  1.370 2.860 1.870 3.020 ;
        RECT  1.530 0.760 1.690 2.560 ;
        RECT  1.250 1.030 1.370 3.020 ;
        RECT  1.210 0.910 1.250 3.020 ;
        RECT  1.050 0.440 1.210 0.720 ;
        RECT  0.970 0.910 1.210 1.190 ;
        RECT  1.190 2.860 1.210 3.020 ;
        RECT  0.910 2.860 1.190 3.160 ;
        RECT  0.370 0.560 1.050 0.720 ;
        RECT  0.850 1.350 1.050 1.630 ;
        RECT  0.810 1.350 0.850 2.700 ;
        RECT  0.650 0.920 0.810 2.700 ;
        RECT  0.370 0.920 0.650 1.080 ;
        RECT  0.570 1.910 0.650 2.700 ;
        RECT  0.090 0.560 0.370 1.080 ;
    END
END ACCSHCINX4TR

MACRO ACCSHCINX2TR
    CLASS CORE ;
    FOREIGN ACCSHCINX2TR 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.600 ;
    SYMMETRY X Y ;
    SITE IBM13SITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.710 0.980 9.930 2.520 ;
        RECT  9.680 2.040 9.710 2.520 ;
        RECT  8.730 2.360 9.680 2.520 ;
        RECT  8.570 1.860 8.730 2.520 ;
        RECT  8.310 1.860 8.570 2.140 ;
        END
        ANTENNADIFFAREA 5.5535 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.190 1.030 12.350 1.310 ;
        RECT  12.030 1.030 12.190 2.890 ;
        RECT  11.680 1.290 12.030 2.890 ;
        RECT  11.390 1.290 11.680 1.450 ;
        RECT  11.100 2.730 11.680 2.890 ;
        RECT  11.230 1.090 11.390 1.450 ;
        RECT  11.110 1.090 11.230 1.310 ;
        RECT  10.820 2.610 11.100 2.890 ;
        END
        ANTENNADIFFAREA 5.0275 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.680 1.240 13.920 2.360 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.830 1.240 13.160 1.640 ;
        END
        ANTENNAGATEAREA 0.2664 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.360 1.340 7.080 1.500 ;
        RECT  6.080 0.850 6.360 1.850 ;
        RECT  5.960 1.570 6.080 1.850 ;
        END
        ANTENNAGATEAREA 0.7824 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.530 0.740 1.810 ;
        RECT  0.440 1.530 0.720 1.960 ;
        END
        ANTENNAGATEAREA 0.264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.370 -0.280 14.000 0.280 ;
        RECT  13.090 -0.280 13.370 0.380 ;
        RECT  8.760 -0.280 13.090 0.280 ;
        RECT  8.480 -0.280 8.760 0.400 ;
        RECT  8.160 -0.280 8.480 0.280 ;
        RECT  7.880 -0.280 8.160 0.400 ;
        RECT  6.640 -0.280 7.880 0.280 ;
        RECT  6.360 -0.280 6.640 0.370 ;
        RECT  1.140 -0.280 6.360 0.280 ;
        RECT  0.860 -0.280 1.140 0.400 ;
        RECT  0.000 -0.280 0.860 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.170 3.320 14.000 3.880 ;
        RECT  12.890 2.120 13.170 3.880 ;
        RECT  7.760 3.320 12.890 3.880 ;
        RECT  7.480 3.260 7.760 3.880 ;
        RECT  2.020 3.320 7.480 3.880 ;
        RECT  1.740 3.200 2.020 3.880 ;
        RECT  0.620 3.320 1.740 3.880 ;
        RECT  0.340 2.120 0.620 3.880 ;
        RECT  0.000 3.320 0.340 3.880 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  13.480 0.540 13.890 0.820 ;
        RECT  13.520 2.540 13.650 3.160 ;
        RECT  13.480 1.800 13.520 3.160 ;
        RECT  13.360 0.540 13.480 3.160 ;
        RECT  13.320 0.540 13.360 1.960 ;
        RECT  12.190 0.540 13.320 0.700 ;
        RECT  12.670 0.860 12.850 1.080 ;
        RECT  12.510 0.860 12.670 3.160 ;
        RECT  12.390 1.910 12.510 3.160 ;
        RECT  12.030 0.450 12.190 0.700 ;
        RECT  9.520 0.450 12.030 0.610 ;
        RECT  11.590 0.770 11.870 1.130 ;
        RECT  10.950 0.770 11.590 0.930 ;
        RECT  11.300 2.240 11.520 2.520 ;
        RECT  10.950 2.240 11.300 2.400 ;
        RECT  10.790 0.770 10.950 2.400 ;
        RECT  10.250 0.770 10.790 0.930 ;
        RECT  10.410 1.300 10.630 3.160 ;
        RECT  8.040 3.000 10.410 3.160 ;
        RECT  10.090 0.770 10.250 2.840 ;
        RECT  8.410 2.680 10.090 2.840 ;
        RECT  9.360 0.450 9.520 1.260 ;
        RECT  9.170 0.980 9.360 1.260 ;
        RECT  8.920 0.440 9.200 0.720 ;
        RECT  9.110 1.100 9.170 1.260 ;
        RECT  8.890 1.100 9.110 2.140 ;
        RECT  7.720 0.560 8.920 0.720 ;
        RECT  7.780 0.890 8.470 1.170 ;
        RECT  8.250 2.300 8.410 2.840 ;
        RECT  6.920 2.300 8.250 2.460 ;
        RECT  6.280 2.620 8.090 2.780 ;
        RECT  7.900 2.940 8.040 3.160 ;
        RECT  6.600 2.940 7.900 3.100 ;
        RECT  7.560 0.890 7.780 2.140 ;
        RECT  7.560 0.440 7.720 0.720 ;
        RECT  6.960 0.440 7.560 0.600 ;
        RECT  7.080 1.980 7.560 2.140 ;
        RECT  7.240 0.760 7.400 1.820 ;
        RECT  7.120 0.760 7.240 1.040 ;
        RECT  6.920 1.660 7.240 1.820 ;
        RECT  6.800 0.440 6.960 0.690 ;
        RECT  6.760 1.660 6.920 2.460 ;
        RECT  5.920 0.530 6.800 0.690 ;
        RECT  6.200 2.180 6.760 2.460 ;
        RECT  6.440 2.940 6.600 3.160 ;
        RECT  2.340 3.000 6.440 3.160 ;
        RECT  2.660 2.620 6.280 2.840 ;
        RECT  5.800 2.010 5.960 2.290 ;
        RECT  5.800 0.530 5.920 1.040 ;
        RECT  5.640 0.530 5.800 2.290 ;
        RECT  4.880 0.530 5.640 0.690 ;
        RECT  5.440 1.920 5.480 2.200 ;
        RECT  5.320 0.900 5.440 2.200 ;
        RECT  5.160 0.900 5.320 2.460 ;
        RECT  2.980 2.300 5.160 2.460 ;
        RECT  4.880 1.980 5.000 2.140 ;
        RECT  4.720 0.530 4.880 2.140 ;
        RECT  4.560 0.760 4.720 1.040 ;
        RECT  4.360 1.920 4.520 2.140 ;
        RECT  4.200 0.440 4.360 2.140 ;
        RECT  3.050 0.440 4.200 0.720 ;
        RECT  3.260 1.920 4.200 2.140 ;
        RECT  2.740 1.020 3.890 1.300 ;
        RECT  1.460 0.440 3.050 0.600 ;
        RECT  2.820 2.080 2.980 2.460 ;
        RECT  2.540 2.080 2.820 2.240 ;
        RECT  2.580 0.760 2.740 1.300 ;
        RECT  2.500 2.400 2.660 2.840 ;
        RECT  1.940 0.760 2.580 0.920 ;
        RECT  2.420 1.960 2.540 2.240 ;
        RECT  1.940 2.400 2.500 2.560 ;
        RECT  2.260 1.080 2.420 2.240 ;
        RECT  2.180 2.880 2.340 3.160 ;
        RECT  2.100 1.080 2.260 1.300 ;
        RECT  1.620 2.880 2.180 3.040 ;
        RECT  1.780 0.760 1.940 2.560 ;
        RECT  1.500 1.030 1.620 3.040 ;
        RECT  1.460 0.910 1.500 3.040 ;
        RECT  1.300 0.440 1.460 0.720 ;
        RECT  1.220 0.910 1.460 1.190 ;
        RECT  1.220 2.760 1.460 3.040 ;
        RECT  0.620 0.560 1.300 0.720 ;
        RECT  1.160 1.350 1.300 1.630 ;
        RECT  1.060 1.350 1.160 2.580 ;
        RECT  0.900 1.140 1.060 2.580 ;
        RECT  0.620 1.140 0.900 1.300 ;
        RECT  0.880 1.910 0.900 2.580 ;
        RECT  0.340 0.560 0.620 1.300 ;
    END
END ACCSHCINX2TR

END LIBRARY
